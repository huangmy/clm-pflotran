netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "timestep fractional area burned for crop" ;
		BAF_CROP:units = "proportion" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "timestep fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned in this timestep" ;
		LFC2:units = "per timestep" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "timestep fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/timestep" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/14/14 18:41:51" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "bandre" ;
		:version = "clm4_5_67" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c130821.nc" ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/14/14" ;

 time_written =
  "18:41:51" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.484872e-14, 4.497019e-14, 4.49466e-14, 4.504447e-14, 4.49902e-14, 
    4.505427e-14, 4.487338e-14, 4.497499e-14, 4.491014e-14, 4.485969e-14, 
    4.523413e-14, 4.504884e-14, 4.542646e-14, 4.530849e-14, 4.560464e-14, 
    4.540809e-14, 4.564424e-14, 4.559901e-14, 4.573518e-14, 4.569619e-14, 
    4.587009e-14, 4.575318e-14, 4.59602e-14, 4.584221e-14, 4.586065e-14, 
    4.574931e-14, 4.508619e-14, 4.521107e-14, 4.507878e-14, 4.50966e-14, 
    4.508862e-14, 4.499131e-14, 4.494222e-14, 4.483946e-14, 4.485813e-14, 
    4.493362e-14, 4.510461e-14, 4.504662e-14, 4.51928e-14, 4.51895e-14, 
    4.5352e-14, 4.527876e-14, 4.555155e-14, 4.547411e-14, 4.569782e-14, 
    4.564159e-14, 4.569517e-14, 4.567893e-14, 4.569538e-14, 4.56129e-14, 
    4.564825e-14, 4.557566e-14, 4.529247e-14, 4.537577e-14, 4.512715e-14, 
    4.497733e-14, 4.487783e-14, 4.480714e-14, 4.481714e-14, 4.483618e-14, 
    4.493406e-14, 4.502604e-14, 4.509608e-14, 4.514291e-14, 4.518903e-14, 
    4.532841e-14, 4.540221e-14, 4.556718e-14, 4.553746e-14, 4.558784e-14, 
    4.563599e-14, 4.571675e-14, 4.570347e-14, 4.573903e-14, 4.558653e-14, 
    4.568789e-14, 4.552054e-14, 4.556632e-14, 4.520142e-14, 4.506227e-14, 
    4.500296e-14, 4.495113e-14, 4.482482e-14, 4.491205e-14, 4.487767e-14, 
    4.495948e-14, 4.501142e-14, 4.498574e-14, 4.514419e-14, 4.508261e-14, 
    4.540658e-14, 4.526715e-14, 4.563038e-14, 4.554357e-14, 4.565118e-14, 
    4.559629e-14, 4.569032e-14, 4.560569e-14, 4.575227e-14, 4.578414e-14, 
    4.576236e-14, 4.584606e-14, 4.5601e-14, 4.569516e-14, 4.498502e-14, 
    4.49892e-14, 4.500873e-14, 4.492288e-14, 4.491763e-14, 4.483895e-14, 
    4.490898e-14, 4.493877e-14, 4.501444e-14, 4.505915e-14, 4.510164e-14, 
    4.519502e-14, 4.529919e-14, 4.544474e-14, 4.554919e-14, 4.561917e-14, 
    4.557627e-14, 4.561414e-14, 4.55718e-14, 4.555196e-14, 4.577219e-14, 
    4.564857e-14, 4.583403e-14, 4.582378e-14, 4.573986e-14, 4.582493e-14, 
    4.499214e-14, 4.496804e-14, 4.488427e-14, 4.494983e-14, 4.483037e-14, 
    4.489724e-14, 4.493566e-14, 4.508386e-14, 4.511643e-14, 4.514659e-14, 
    4.520614e-14, 4.528251e-14, 4.541635e-14, 4.553267e-14, 4.56388e-14, 
    4.563103e-14, 4.563376e-14, 4.565745e-14, 4.559876e-14, 4.566708e-14, 
    4.567853e-14, 4.564857e-14, 4.582241e-14, 4.577277e-14, 4.582356e-14, 
    4.579125e-14, 4.497588e-14, 4.501644e-14, 4.499452e-14, 4.503573e-14, 
    4.500669e-14, 4.513571e-14, 4.517436e-14, 4.535511e-14, 4.5281e-14, 
    4.539896e-14, 4.5293e-14, 4.531177e-14, 4.540274e-14, 4.529874e-14, 
    4.552626e-14, 4.5372e-14, 4.565837e-14, 4.550447e-14, 4.5668e-14, 
    4.563834e-14, 4.568746e-14, 4.573142e-14, 4.578672e-14, 4.588865e-14, 
    4.586506e-14, 4.595027e-14, 4.507689e-14, 4.512944e-14, 4.512484e-14, 
    4.517983e-14, 4.522047e-14, 4.530854e-14, 4.544963e-14, 4.53966e-14, 
    4.549396e-14, 4.551349e-14, 4.536558e-14, 4.545639e-14, 4.516461e-14, 
    4.521178e-14, 4.518372e-14, 4.508102e-14, 4.540879e-14, 4.524068e-14, 
    4.555091e-14, 4.546002e-14, 4.572515e-14, 4.559333e-14, 4.585207e-14, 
    4.596242e-14, 4.60663e-14, 4.618743e-14, 4.515814e-14, 4.512244e-14, 
    4.518637e-14, 4.527471e-14, 4.53567e-14, 4.546556e-14, 4.547671e-14, 
    4.549708e-14, 4.554984e-14, 4.559419e-14, 4.550349e-14, 4.560531e-14, 
    4.522266e-14, 4.542338e-14, 4.510892e-14, 4.520366e-14, 4.526952e-14, 
    4.524066e-14, 4.539055e-14, 4.542584e-14, 4.556909e-14, 4.549509e-14, 
    4.593517e-14, 4.574066e-14, 4.627966e-14, 4.612929e-14, 4.510996e-14, 
    4.515802e-14, 4.532512e-14, 4.524565e-14, 4.547284e-14, 4.552868e-14, 
    4.557405e-14, 4.563201e-14, 4.563829e-14, 4.567262e-14, 4.561636e-14, 
    4.567041e-14, 4.546579e-14, 4.555727e-14, 4.530606e-14, 4.536724e-14, 
    4.533911e-14, 4.530823e-14, 4.540352e-14, 4.550492e-14, 4.550713e-14, 
    4.553958e-14, 4.5631e-14, 4.547376e-14, 4.596017e-14, 4.565993e-14, 
    4.521041e-14, 4.530284e-14, 4.531609e-14, 4.528029e-14, 4.552308e-14, 
    4.543516e-14, 4.567179e-14, 4.560789e-14, 4.571258e-14, 4.566056e-14, 
    4.565291e-14, 4.558607e-14, 4.554443e-14, 4.543919e-14, 4.535347e-14, 
    4.528549e-14, 4.53013e-14, 4.537598e-14, 4.551112e-14, 4.563884e-14, 
    4.561086e-14, 4.570463e-14, 4.545638e-14, 4.55605e-14, 4.552027e-14, 
    4.562519e-14, 4.539518e-14, 4.559095e-14, 4.534507e-14, 4.536666e-14, 
    4.543342e-14, 4.556753e-14, 4.559726e-14, 4.56289e-14, 4.560939e-14, 
    4.551456e-14, 4.549904e-14, 4.54318e-14, 4.541321e-14, 4.536197e-14, 
    4.53195e-14, 4.535829e-14, 4.5399e-14, 4.551462e-14, 4.561866e-14, 
    4.573204e-14, 4.575978e-14, 4.589195e-14, 4.578431e-14, 4.596183e-14, 
    4.581083e-14, 4.607213e-14, 4.560234e-14, 4.580648e-14, 4.543647e-14, 
    4.54764e-14, 4.554852e-14, 4.571391e-14, 4.56247e-14, 4.572905e-14, 
    4.549843e-14, 4.537853e-14, 4.534754e-14, 4.528962e-14, 4.534887e-14, 
    4.534405e-14, 4.540072e-14, 4.538251e-14, 4.551846e-14, 4.544546e-14, 
    4.56527e-14, 4.572824e-14, 4.594133e-14, 4.607172e-14, 4.620437e-14, 
    4.626286e-14, 4.628066e-14, 4.628809e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.895644e-14, -1.897863e-14, -1.89743e-14, -1.89922e-14, -1.898225e-14, 
    -1.899399e-14, -1.896091e-14, -1.897953e-14, -1.896763e-14, -1.89584e-14, 
    -1.902693e-14, -1.8993e-14, -1.906175e-14, -1.904026e-14, -1.909404e-14, 
    -1.905844e-14, -1.910119e-14, -1.909295e-14, -1.911756e-14, 
    -1.911051e-14, -1.914205e-14, -1.912081e-14, -1.915824e-14, 
    -1.913695e-14, -1.914031e-14, -1.912012e-14, -1.899977e-14, 
    -1.902273e-14, -1.899842e-14, -1.90017e-14, -1.900021e-14, -1.898248e-14, 
    -1.897358e-14, -1.895469e-14, -1.895811e-14, -1.897195e-14, 
    -1.900317e-14, -1.899254e-14, -1.901917e-14, -1.901857e-14, 
    -1.904816e-14, -1.903483e-14, -1.908436e-14, -1.907029e-14, -1.91108e-14, 
    -1.910065e-14, -1.911034e-14, -1.910739e-14, -1.911038e-14, 
    -1.909547e-14, -1.910187e-14, -1.908871e-14, -1.903734e-14, 
    -1.905249e-14, -1.900726e-14, -1.898003e-14, -1.896174e-14, 
    -1.894879e-14, -1.895062e-14, -1.895413e-14, -1.897204e-14, 
    -1.898879e-14, -1.900155e-14, -1.901009e-14, -1.901848e-14, 
    -1.904401e-14, -1.905734e-14, -1.908723e-14, -1.908179e-14, 
    -1.909096e-14, -1.909963e-14, -1.911425e-14, -1.911184e-14, 
    -1.911828e-14, -1.909068e-14, -1.910905e-14, -1.90787e-14, -1.908702e-14, 
    -1.902099e-14, -1.89954e-14, -1.89847e-14, -1.897514e-14, -1.895203e-14, 
    -1.896801e-14, -1.896172e-14, -1.897663e-14, -1.898612e-14, 
    -1.898142e-14, -1.901032e-14, -1.89991e-14, -1.905813e-14, -1.903276e-14, 
    -1.909862e-14, -1.90829e-14, -1.910238e-14, -1.909243e-14, -1.910948e-14, 
    -1.909414e-14, -1.912066e-14, -1.912645e-14, -1.91225e-14, -1.913759e-14, 
    -1.909329e-14, -1.911036e-14, -1.89813e-14, -1.898207e-14, -1.898562e-14, 
    -1.896999e-14, -1.896902e-14, -1.895461e-14, -1.896742e-14, 
    -1.897288e-14, -1.898665e-14, -1.899483e-14, -1.900258e-14, -1.90196e-14, 
    -1.90386e-14, -1.906502e-14, -1.908392e-14, -1.909657e-14, -1.90888e-14, 
    -1.909567e-14, -1.9088e-14, -1.90844e-14, -1.91243e-14, -1.910194e-14, 
    -1.913543e-14, -1.913357e-14, -1.911845e-14, -1.913378e-14, -1.89826e-14, 
    -1.897818e-14, -1.896291e-14, -1.897487e-14, -1.895304e-14, 
    -1.896529e-14, -1.897235e-14, -1.899939e-14, -1.900526e-14, 
    -1.901078e-14, -1.902161e-14, -1.903552e-14, -1.905986e-14, 
    -1.908096e-14, -1.910013e-14, -1.909872e-14, -1.909922e-14, 
    -1.910352e-14, -1.909289e-14, -1.910526e-14, -1.910735e-14, 
    -1.910191e-14, -1.913332e-14, -1.912436e-14, -1.913353e-14, 
    -1.912769e-14, -1.897961e-14, -1.898703e-14, -1.898303e-14, 
    -1.899057e-14, -1.898528e-14, -1.900886e-14, -1.901591e-14, 
    -1.904879e-14, -1.903526e-14, -1.905672e-14, -1.903742e-14, 
    -1.904086e-14, -1.905751e-14, -1.903845e-14, -1.907983e-14, 
    -1.905189e-14, -1.910368e-14, -1.907594e-14, -1.910542e-14, 
    -1.910004e-14, -1.910893e-14, -1.91169e-14, -1.912688e-14, -1.914532e-14, 
    -1.914105e-14, -1.915641e-14, -1.899806e-14, -1.900768e-14, 
    -1.900679e-14, -1.901682e-14, -1.902424e-14, -1.904024e-14, 
    -1.906588e-14, -1.905623e-14, -1.907389e-14, -1.907744e-14, 
    -1.905059e-14, -1.906713e-14, -1.901408e-14, -1.902272e-14, 
    -1.901755e-14, -1.899884e-14, -1.905852e-14, -1.902798e-14, 
    -1.908424e-14, -1.906775e-14, -1.911577e-14, -1.909197e-14, -1.91387e-14, 
    -1.915871e-14, -1.917729e-14, -1.919919e-14, -1.901288e-14, 
    -1.900635e-14, -1.9018e-14, -1.903416e-14, -1.904901e-14, -1.906877e-14, 
    -1.907076e-14, -1.907447e-14, -1.908402e-14, -1.909206e-14, 
    -1.907568e-14, -1.909407e-14, -1.902481e-14, -1.906114e-14, 
    -1.900392e-14, -1.902125e-14, -1.903319e-14, -1.902791e-14, 
    -1.905512e-14, -1.906153e-14, -1.908756e-14, -1.907409e-14, 
    -1.915381e-14, -1.911864e-14, -1.921567e-14, -1.918871e-14, 
    -1.900408e-14, -1.901284e-14, -1.90433e-14, -1.902882e-14, -1.907006e-14, 
    -1.90802e-14, -1.90884e-14, -1.909894e-14, -1.910004e-14, -1.910627e-14, 
    -1.909607e-14, -1.910585e-14, -1.906881e-14, -1.908538e-14, 
    -1.903977e-14, -1.905092e-14, -1.904578e-14, -1.904017e-14, 
    -1.905748e-14, -1.907595e-14, -1.907628e-14, -1.908221e-14, 
    -1.909901e-14, -1.907023e-14, -1.915847e-14, -1.910421e-14, 
    -1.902238e-14, -1.903929e-14, -1.904162e-14, -1.903509e-14, 
    -1.907919e-14, -1.906325e-14, -1.910611e-14, -1.909453e-14, 
    -1.911348e-14, -1.910408e-14, -1.91027e-14, -1.909059e-14, -1.908306e-14, 
    -1.906399e-14, -1.904843e-14, -1.903603e-14, -1.903891e-14, 
    -1.905252e-14, -1.907707e-14, -1.910017e-14, -1.909513e-14, 
    -1.911204e-14, -1.906708e-14, -1.9086e-14, -1.907871e-14, -1.909768e-14, 
    -1.905599e-14, -1.909171e-14, -1.904686e-14, -1.905079e-14, 
    -1.906293e-14, -1.908733e-14, -1.909261e-14, -1.909838e-14, -1.90948e-14, 
    -1.907768e-14, -1.907483e-14, -1.906262e-14, -1.905927e-14, 
    -1.904993e-14, -1.904221e-14, -1.904928e-14, -1.905671e-14, 
    -1.907765e-14, -1.909653e-14, -1.911703e-14, -1.912201e-14, 
    -1.914605e-14, -1.912658e-14, -1.915878e-14, -1.913155e-14, 
    -1.917856e-14, -1.909368e-14, -1.913061e-14, -1.906346e-14, -1.90707e-14, 
    -1.908386e-14, -1.911382e-14, -1.909759e-14, -1.911654e-14, 
    -1.907472e-14, -1.905302e-14, -1.904731e-14, -1.90368e-14, -1.904756e-14, 
    -1.904668e-14, -1.905697e-14, -1.905366e-14, -1.907835e-14, 
    -1.906509e-14, -1.910268e-14, -1.911637e-14, -1.915483e-14, 
    -1.917835e-14, -1.920212e-14, -1.921263e-14, -1.921581e-14, -1.921715e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.516502e-11, 1.515783e-11, 1.515932e-11, 1.515286e-11, 1.515655e-11, 
    1.515217e-11, 1.516366e-11, 1.515751e-11, 1.516153e-11, 1.516443e-11, 
    1.513794e-11, 1.515256e-11, 1.503708e-11, 1.503615e-11, 1.503342e-11, 
    1.503709e-11, 1.503173e-11, 1.503366e-11, 1.502656e-11, 1.502901e-11, 
    1.501535e-11, 1.502531e-11, 1.500548e-11, 1.501803e-11, 1.501629e-11, 
    1.502558e-11, 1.514989e-11, 1.513993e-11, 1.515043e-11, 1.514911e-11, 
    1.514971e-11, 1.515646e-11, 1.515957e-11, 1.516554e-11, 1.516452e-11, 
    1.516011e-11, 1.514851e-11, 1.515273e-11, 1.514155e-11, 1.514182e-11, 
    1.50368e-11, 1.503552e-11, 1.50352e-11, 1.503675e-11, 1.502891e-11, 
    1.503187e-11, 1.502906e-11, 1.502998e-11, 1.502905e-11, 1.503311e-11, 
    1.503155e-11, 1.503448e-11, 1.503583e-11, 1.5037e-11, 1.51468e-11, 
    1.515734e-11, 1.51634e-11, 1.516726e-11, 1.516673e-11, 1.516571e-11, 
    1.516008e-11, 1.515415e-11, 1.514916e-11, 1.514558e-11, 1.514186e-11, 
    1.503645e-11, 1.503709e-11, 1.503473e-11, 1.503558e-11, 1.503405e-11, 
    1.503213e-11, 1.502775e-11, 1.502857e-11, 1.502629e-11, 1.503411e-11, 
    1.502947e-11, 1.503597e-11, 1.503478e-11, 1.514074e-11, 1.515162e-11, 
    1.515567e-11, 1.515903e-11, 1.516632e-11, 1.516141e-11, 1.516341e-11, 
    1.515852e-11, 1.515514e-11, 1.515684e-11, 1.514548e-11, 1.515015e-11, 
    1.50371e-11, 1.503522e-11, 1.503238e-11, 1.503542e-11, 1.503142e-11, 
    1.503377e-11, 1.502934e-11, 1.503341e-11, 1.502537e-11, 1.502298e-11, 
    1.502464e-11, 1.501769e-11, 1.503359e-11, 1.502906e-11, 1.515689e-11, 
    1.515661e-11, 1.515532e-11, 1.516076e-11, 1.516108e-11, 1.516557e-11, 
    1.51616e-11, 1.51598e-11, 1.515495e-11, 1.515184e-11, 1.514874e-11, 
    1.514135e-11, 1.503596e-11, 1.5037e-11, 1.503527e-11, 1.503287e-11, 
    1.503446e-11, 1.503307e-11, 1.503461e-11, 1.50352e-11, 1.50239e-11, 
    1.503153e-11, 1.501879e-11, 1.50197e-11, 1.502623e-11, 1.50196e-11, 
    1.515642e-11, 1.515798e-11, 1.516304e-11, 1.515913e-11, 1.516603e-11, 
    1.516228e-11, 1.515998e-11, 1.515004e-11, 1.514763e-11, 1.514529e-11, 
    1.514042e-11, 1.50356e-11, 1.503711e-11, 1.503568e-11, 1.5032e-11, 
    1.503236e-11, 1.503223e-11, 1.50311e-11, 1.503367e-11, 1.503061e-11, 
    1.503e-11, 1.503154e-11, 1.501982e-11, 1.502387e-11, 1.501972e-11, 
    1.502243e-11, 1.515748e-11, 1.51548e-11, 1.515627e-11, 1.515348e-11, 
    1.515545e-11, 1.514612e-11, 1.514303e-11, 1.503681e-11, 1.503556e-11, 
    1.50371e-11, 1.503584e-11, 1.503621e-11, 1.503708e-11, 1.503597e-11, 
    1.503582e-11, 1.503695e-11, 1.503106e-11, 1.503625e-11, 1.503057e-11, 
    1.503202e-11, 1.502951e-11, 1.50268e-11, 1.502279e-11, 1.50135e-11, 
    1.501587e-11, 1.500668e-11, 1.515057e-11, 1.514662e-11, 1.514699e-11, 
    1.514262e-11, 1.51392e-11, 1.503616e-11, 1.503698e-11, 1.503711e-11, 
    1.503647e-11, 1.503611e-11, 1.503694e-11, 1.503692e-11, 1.514384e-11, 
    1.513992e-11, 1.514229e-11, 1.515026e-11, 1.503711e-11, 1.513742e-11, 
    1.503522e-11, 1.503689e-11, 1.502721e-11, 1.503385e-11, 1.501712e-11, 
    1.500519e-11, 1.499124e-11, 1.497129e-11, 1.514437e-11, 1.514717e-11, 
    1.514208e-11, 1.50354e-11, 1.503685e-11, 1.503684e-11, 1.503671e-11, 
    1.503641e-11, 1.503526e-11, 1.503384e-11, 1.503629e-11, 1.503342e-11, 
    1.513895e-11, 1.50371e-11, 1.514819e-11, 1.51406e-11, 1.503528e-11, 
    1.513744e-11, 1.503709e-11, 1.503711e-11, 1.503468e-11, 1.503645e-11, 
    1.50084e-11, 1.502616e-11, 1.495345e-11, 1.498135e-11, 1.514812e-11, 
    1.514439e-11, 1.503643e-11, 1.5137e-11, 1.503676e-11, 1.503578e-11, 
    1.503454e-11, 1.50323e-11, 1.503202e-11, 1.503032e-11, 1.503298e-11, 
    1.503044e-11, 1.503683e-11, 1.503504e-11, 1.503611e-11, 1.503694e-11, 
    1.503665e-11, 1.503615e-11, 1.503712e-11, 1.503626e-11, 1.503624e-11, 
    1.503551e-11, 1.503227e-11, 1.503675e-11, 1.500542e-11, 1.503091e-11, 
    1.514006e-11, 1.503602e-11, 1.503629e-11, 1.503556e-11, 1.503591e-11, 
    1.503707e-11, 1.503037e-11, 1.503332e-11, 1.502802e-11, 1.503095e-11, 
    1.503133e-11, 1.503413e-11, 1.50354e-11, 1.503704e-11, 1.503681e-11, 
    1.503568e-11, 1.503602e-11, 1.5037e-11, 1.503614e-11, 1.503199e-11, 
    1.503319e-11, 1.502851e-11, 1.503693e-11, 1.503494e-11, 1.503596e-11, 
    1.503261e-11, 1.50371e-11, 1.503389e-11, 1.503673e-11, 1.503695e-11, 
    1.503708e-11, 1.503471e-11, 1.503373e-11, 1.503244e-11, 1.503326e-11, 
    1.503608e-11, 1.503638e-11, 1.503709e-11, 1.503712e-11, 1.503691e-11, 
    1.503635e-11, 1.503687e-11, 1.50371e-11, 1.503609e-11, 1.503287e-11, 
    1.502676e-11, 1.502484e-11, 1.501312e-11, 1.502294e-11, 1.500521e-11, 
    1.502072e-11, 1.49903e-11, 1.50335e-11, 1.502114e-11, 1.503707e-11, 
    1.503672e-11, 1.503527e-11, 1.502791e-11, 1.503263e-11, 1.502694e-11, 
    1.503639e-11, 1.503701e-11, 1.503675e-11, 1.503577e-11, 1.503677e-11, 
    1.503671e-11, 1.503712e-11, 1.503705e-11, 1.503601e-11, 1.503702e-11, 
    1.503133e-11, 1.5027e-11, 1.500772e-11, 1.49904e-11, 1.496822e-11, 
    1.495689e-11, 1.495326e-11, 1.495171e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931945e-23, 1.931947e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.93194e-23, 1.931941e-23, 1.931939e-23, 1.93194e-23, 1.93194e-23, 
    1.931941e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931945e-23, 1.931944e-23, 1.931946e-23, 
    1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931945e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.931941e-23, 1.93194e-23, 1.931942e-23, 1.931941e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.93194e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931941e-23, 1.931942e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931941e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931944e-23, 1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.93194e-23, 
    1.93194e-23, 1.931939e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931943e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.93194e-23, 
    1.931939e-23, 1.931938e-23, 1.931937e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931945e-23, 1.931944e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 
    1.931939e-23, 1.931941e-23, 1.931936e-23, 1.931938e-23, 1.931946e-23, 
    1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931939e-23, 1.931942e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 
    1.931944e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 
    1.931942e-23, 1.931944e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931941e-23, 1.931941e-23, 1.93194e-23, 1.931941e-23, 1.931939e-23, 
    1.93194e-23, 1.931938e-23, 1.931942e-23, 1.93194e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 
    1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931941e-23, 1.931939e-23, 1.931938e-23, 1.931937e-23, 
    1.931937e-23, 1.931936e-23, 1.931936e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.975377e-24, 1.975379e-24, 1.975374e-24, 1.975376e-24, 1.975372e-24, 
    1.975375e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975371e-24, 
    1.975369e-24, 1.975371e-24, 1.975368e-24, 1.97537e-24, 1.975369e-24, 
    1.975371e-24, 1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975378e-24, 
    1.975378e-24, 1.975379e-24, 1.97538e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 
    1.975375e-24, 1.975376e-24, 1.975373e-24, 1.975374e-24, 1.975371e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 1.975378e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975377e-24, 
    1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975373e-24, 
    1.975371e-24, 1.975373e-24, 1.975373e-24, 1.975377e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975375e-24, 1.975376e-24, 1.975372e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 1.97537e-24, 
    1.975371e-24, 1.97537e-24, 1.975372e-24, 1.975371e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 1.975372e-24, 
    1.975373e-24, 1.975372e-24, 1.975373e-24, 1.975373e-24, 1.97537e-24, 
    1.975372e-24, 1.97537e-24, 1.97537e-24, 1.975371e-24, 1.97537e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975371e-24, 1.975372e-24, 1.97537e-24, 1.97537e-24, 1.97537e-24, 
    1.97537e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975375e-24, 1.975376e-24, 
    1.975375e-24, 1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975376e-24, 
    1.975373e-24, 1.975375e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.97537e-24, 1.975369e-24, 
    1.975369e-24, 1.975368e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975375e-24, 1.975374e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 
    1.975373e-24, 1.975374e-24, 1.975371e-24, 1.975372e-24, 1.975369e-24, 
    1.975368e-24, 1.975367e-24, 1.975365e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975377e-24, 1.975374e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975374e-24, 
    1.975368e-24, 1.975371e-24, 1.975365e-24, 1.975366e-24, 1.975378e-24, 
    1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975374e-24, 1.975373e-24, 
    1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975372e-24, 1.975374e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975368e-24, 1.975372e-24, 
    1.975377e-24, 1.975376e-24, 1.975376e-24, 1.975376e-24, 1.975373e-24, 
    1.975374e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975373e-24, 1.975374e-24, 1.975375e-24, 
    1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975374e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975375e-24, 1.975373e-24, 1.975375e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975373e-24, 1.975374e-24, 1.975374e-24, 1.975375e-24, 1.975375e-24, 
    1.975376e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975371e-24, 1.975371e-24, 1.975369e-24, 1.97537e-24, 1.975368e-24, 
    1.97537e-24, 1.975367e-24, 1.975372e-24, 1.97537e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 
    1.975374e-24, 1.975375e-24, 1.975375e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975374e-24, 
    1.975372e-24, 1.975371e-24, 1.975368e-24, 1.975367e-24, 1.975365e-24, 
    1.975365e-24, 1.975365e-24, 1.975364e-24 ;

 CONC_CH4_SAT =
  8.459784e-08, 8.470361e-08, 8.468301e-08, 8.47683e-08, 8.472092e-08, 
    8.477681e-08, 8.461919e-08, 8.47079e-08, 8.465123e-08, 8.460722e-08, 
    8.493365e-08, 8.477208e-08, 8.509976e-08, 8.499739e-08, 8.525374e-08, 
    8.508398e-08, 8.528783e-08, 8.52486e-08, 8.536595e-08, 8.533235e-08, 
    8.54826e-08, 8.538145e-08, 8.555985e-08, 8.545833e-08, 8.547433e-08, 
    8.537815e-08, 8.480441e-08, 8.491364e-08, 8.479798e-08, 8.481356e-08, 
    8.480652e-08, 8.472198e-08, 8.467948e-08, 8.458957e-08, 8.460587e-08, 
    8.46718e-08, 8.482056e-08, 8.476997e-08, 8.48969e-08, 8.489403e-08, 
    8.503504e-08, 8.497153e-08, 8.520762e-08, 8.514061e-08, 8.533375e-08, 
    8.528531e-08, 8.533152e-08, 8.531748e-08, 8.533171e-08, 8.526061e-08, 
    8.52911e-08, 8.52284e-08, 8.498348e-08, 8.50557e-08, 8.484006e-08, 
    8.471021e-08, 8.462313e-08, 8.456142e-08, 8.457015e-08, 8.458684e-08, 
    8.467219e-08, 8.475207e-08, 8.481292e-08, 8.48536e-08, 8.489362e-08, 
    8.501514e-08, 8.507877e-08, 8.522128e-08, 8.519539e-08, 8.523908e-08, 
    8.528047e-08, 8.535015e-08, 8.533866e-08, 8.536938e-08, 8.523777e-08, 
    8.532536e-08, 8.518069e-08, 8.522034e-08, 8.490532e-08, 8.478358e-08, 
    8.473244e-08, 8.4687e-08, 8.457688e-08, 8.4653e-08, 8.462303e-08, 
    8.469412e-08, 8.473936e-08, 8.471696e-08, 8.485471e-08, 8.480124e-08, 
    8.508254e-08, 8.496161e-08, 8.527564e-08, 8.520069e-08, 8.529356e-08, 
    8.524616e-08, 8.532741e-08, 8.525429e-08, 8.538074e-08, 8.540832e-08, 
    8.538949e-08, 8.546148e-08, 8.525025e-08, 8.53316e-08, 8.471637e-08, 
    8.472003e-08, 8.473697e-08, 8.466245e-08, 8.465783e-08, 8.458917e-08, 
    8.46502e-08, 8.467623e-08, 8.474191e-08, 8.478087e-08, 8.481782e-08, 
    8.489891e-08, 8.498944e-08, 8.511542e-08, 8.520556e-08, 8.526591e-08, 
    8.522886e-08, 8.526158e-08, 8.522503e-08, 8.520786e-08, 8.539804e-08, 
    8.529143e-08, 8.545113e-08, 8.544228e-08, 8.537014e-08, 8.544328e-08, 
    8.472259e-08, 8.470155e-08, 8.462871e-08, 8.468572e-08, 8.458167e-08, 
    8.464005e-08, 8.467364e-08, 8.480254e-08, 8.483061e-08, 8.485688e-08, 
    8.490852e-08, 8.497479e-08, 8.509083e-08, 8.519139e-08, 8.528284e-08, 
    8.527613e-08, 8.52785e-08, 8.529899e-08, 8.524833e-08, 8.53073e-08, 
    8.531726e-08, 8.529132e-08, 8.54411e-08, 8.539836e-08, 8.54421e-08, 
    8.541425e-08, 8.470837e-08, 8.474371e-08, 8.472463e-08, 8.476055e-08, 
    8.473531e-08, 8.484765e-08, 8.488127e-08, 8.503797e-08, 8.497354e-08, 
    8.507582e-08, 8.498387e-08, 8.500022e-08, 8.507951e-08, 8.498879e-08, 
    8.518601e-08, 8.505272e-08, 8.529979e-08, 8.51674e-08, 8.530809e-08, 
    8.528245e-08, 8.532481e-08, 8.53628e-08, 8.541039e-08, 8.549829e-08, 
    8.547791e-08, 8.555118e-08, 8.479627e-08, 8.484209e-08, 8.483789e-08, 
    8.488568e-08, 8.492102e-08, 8.49973e-08, 8.511954e-08, 8.507357e-08, 
    8.515774e-08, 8.517468e-08, 8.504668e-08, 8.512546e-08, 8.48726e-08, 
    8.491372e-08, 8.488912e-08, 8.479997e-08, 8.508438e-08, 8.493878e-08, 
    8.520708e-08, 8.512848e-08, 8.535741e-08, 8.524388e-08, 8.546674e-08, 
    8.556202e-08, 8.565076e-08, 8.575505e-08, 8.486689e-08, 8.48358e-08, 
    8.489131e-08, 8.496827e-08, 8.503909e-08, 8.51333e-08, 8.514284e-08, 
    8.516051e-08, 8.520604e-08, 8.524436e-08, 8.516624e-08, 8.525394e-08, 
    8.492357e-08, 8.509692e-08, 8.482419e-08, 8.490672e-08, 8.496367e-08, 
    8.493854e-08, 8.506827e-08, 8.509883e-08, 8.522287e-08, 8.515871e-08, 
    8.553867e-08, 8.537104e-08, 8.583374e-08, 8.57051e-08, 8.482498e-08, 
    8.486671e-08, 8.501186e-08, 8.494284e-08, 8.51395e-08, 8.518783e-08, 
    8.522694e-08, 8.527714e-08, 8.528243e-08, 8.531212e-08, 8.526348e-08, 
    8.531014e-08, 8.51335e-08, 8.521251e-08, 8.499511e-08, 8.504822e-08, 
    8.502374e-08, 8.499699e-08, 8.507952e-08, 8.516751e-08, 8.516914e-08, 
    8.519736e-08, 8.527721e-08, 8.514029e-08, 8.556071e-08, 8.530203e-08, 
    8.491219e-08, 8.499271e-08, 8.500389e-08, 8.497278e-08, 8.5183e-08, 
    8.510699e-08, 8.531136e-08, 8.525618e-08, 8.534649e-08, 8.530166e-08, 
    8.529507e-08, 8.523735e-08, 8.520144e-08, 8.511052e-08, 8.503633e-08, 
    8.497727e-08, 8.499099e-08, 8.505583e-08, 8.517284e-08, 8.528303e-08, 
    8.525895e-08, 8.533963e-08, 8.512528e-08, 8.521543e-08, 8.518069e-08, 
    8.527116e-08, 8.507239e-08, 8.524248e-08, 8.502889e-08, 8.504762e-08, 
    8.510548e-08, 8.522171e-08, 8.5247e-08, 8.527445e-08, 8.525746e-08, 
    8.517575e-08, 8.516223e-08, 8.510401e-08, 8.508804e-08, 8.504352e-08, 
    8.500675e-08, 8.504041e-08, 8.507579e-08, 8.517569e-08, 8.526563e-08, 
    8.536338e-08, 8.538716e-08, 8.550163e-08, 8.540882e-08, 8.556219e-08, 
    8.543235e-08, 8.565657e-08, 8.525194e-08, 8.542803e-08, 8.510802e-08, 
    8.514256e-08, 8.520522e-08, 8.534803e-08, 8.527073e-08, 8.536099e-08, 
    8.516169e-08, 8.505819e-08, 8.503106e-08, 8.49809e-08, 8.503221e-08, 
    8.502803e-08, 8.507708e-08, 8.50613e-08, 8.517899e-08, 8.511581e-08, 
    8.529497e-08, 8.536022e-08, 8.55436e-08, 8.565573e-08, 8.576914e-08, 
    8.581924e-08, 8.583445e-08, 8.584082e-08,
  2.315453e-10, 2.321432e-10, 2.320267e-10, 2.325093e-10, 2.322412e-10, 
    2.325575e-10, 2.31666e-10, 2.321674e-10, 2.318471e-10, 2.315984e-10, 
    2.334503e-10, 2.325307e-10, 2.344015e-10, 2.338154e-10, 2.35285e-10, 
    2.34311e-10, 2.354809e-10, 2.352556e-10, 2.359302e-10, 2.35737e-10, 
    2.366014e-10, 2.360194e-10, 2.370469e-10, 2.364618e-10, 2.365538e-10, 
    2.360004e-10, 2.327139e-10, 2.333359e-10, 2.326775e-10, 2.327657e-10, 
    2.327258e-10, 2.322472e-10, 2.320066e-10, 2.314988e-10, 2.315908e-10, 
    2.319633e-10, 2.328053e-10, 2.325188e-10, 2.332408e-10, 2.332245e-10, 
    2.34031e-10, 2.336675e-10, 2.350204e-10, 2.346359e-10, 2.35745e-10, 
    2.354665e-10, 2.357322e-10, 2.356515e-10, 2.357332e-10, 2.353246e-10, 
    2.354998e-10, 2.351397e-10, 2.337358e-10, 2.341492e-10, 2.329161e-10, 
    2.321803e-10, 2.316883e-10, 2.313398e-10, 2.313891e-10, 2.314832e-10, 
    2.319655e-10, 2.324175e-10, 2.327621e-10, 2.329935e-10, 2.332221e-10, 
    2.339167e-10, 2.342812e-10, 2.350987e-10, 2.349502e-10, 2.352009e-10, 
    2.354388e-10, 2.358393e-10, 2.357732e-10, 2.359498e-10, 2.351935e-10, 
    2.356967e-10, 2.348659e-10, 2.350934e-10, 2.332884e-10, 2.325959e-10, 
    2.323061e-10, 2.320493e-10, 2.31427e-10, 2.31857e-10, 2.316877e-10, 
    2.320897e-10, 2.323456e-10, 2.322189e-10, 2.329999e-10, 2.32696e-10, 
    2.343029e-10, 2.336107e-10, 2.35411e-10, 2.349806e-10, 2.35514e-10, 
    2.352417e-10, 2.357085e-10, 2.352884e-10, 2.360152e-10, 2.361738e-10, 
    2.360655e-10, 2.3648e-10, 2.352652e-10, 2.357326e-10, 2.322155e-10, 
    2.322362e-10, 2.323321e-10, 2.319104e-10, 2.318844e-10, 2.314964e-10, 
    2.318413e-10, 2.319884e-10, 2.323601e-10, 2.325806e-10, 2.327899e-10, 
    2.332523e-10, 2.337698e-10, 2.344914e-10, 2.350086e-10, 2.353551e-10, 
    2.351424e-10, 2.353303e-10, 2.351204e-10, 2.350218e-10, 2.361147e-10, 
    2.355017e-10, 2.364204e-10, 2.363695e-10, 2.359542e-10, 2.363752e-10, 
    2.322507e-10, 2.321317e-10, 2.317198e-10, 2.320422e-10, 2.314541e-10, 
    2.317839e-10, 2.319737e-10, 2.327032e-10, 2.328624e-10, 2.330122e-10, 
    2.333072e-10, 2.336862e-10, 2.343505e-10, 2.349272e-10, 2.354524e-10, 
    2.354139e-10, 2.354275e-10, 2.355452e-10, 2.352541e-10, 2.355929e-10, 
    2.356501e-10, 2.355011e-10, 2.363627e-10, 2.361166e-10, 2.363684e-10, 
    2.362081e-10, 2.321703e-10, 2.323702e-10, 2.322623e-10, 2.324655e-10, 
    2.323226e-10, 2.329593e-10, 2.331513e-10, 2.340476e-10, 2.336789e-10, 
    2.342644e-10, 2.337381e-10, 2.338316e-10, 2.342853e-10, 2.337663e-10, 
    2.348962e-10, 2.341319e-10, 2.355498e-10, 2.347892e-10, 2.355975e-10, 
    2.354502e-10, 2.356936e-10, 2.35912e-10, 2.361858e-10, 2.366919e-10, 
    2.365746e-10, 2.369969e-10, 2.326678e-10, 2.329276e-10, 2.329038e-10, 
    2.331767e-10, 2.333786e-10, 2.33815e-10, 2.345151e-10, 2.342517e-10, 
    2.347343e-10, 2.348314e-10, 2.340977e-10, 2.34549e-10, 2.331019e-10, 
    2.333368e-10, 2.331964e-10, 2.326887e-10, 2.343135e-10, 2.3348e-10, 
    2.350173e-10, 2.345663e-10, 2.35881e-10, 2.352284e-10, 2.365102e-10, 
    2.370592e-10, 2.375716e-10, 2.381739e-10, 2.330694e-10, 2.328919e-10, 
    2.332089e-10, 2.336487e-10, 2.340542e-10, 2.34594e-10, 2.346488e-10, 
    2.347501e-10, 2.350114e-10, 2.352314e-10, 2.347828e-10, 2.352864e-10, 
    2.333927e-10, 2.343854e-10, 2.328259e-10, 2.332967e-10, 2.336224e-10, 
    2.334788e-10, 2.342214e-10, 2.343965e-10, 2.351079e-10, 2.347398e-10, 
    2.369244e-10, 2.359592e-10, 2.386294e-10, 2.378853e-10, 2.328305e-10, 
    2.330684e-10, 2.338982e-10, 2.335034e-10, 2.346296e-10, 2.349068e-10, 
    2.351314e-10, 2.354195e-10, 2.3545e-10, 2.356206e-10, 2.353412e-10, 
    2.356093e-10, 2.345951e-10, 2.350485e-10, 2.338024e-10, 2.341065e-10, 
    2.339663e-10, 2.338132e-10, 2.342858e-10, 2.347901e-10, 2.347996e-10, 
    2.349614e-10, 2.354194e-10, 2.346341e-10, 2.370512e-10, 2.35562e-10, 
    2.333282e-10, 2.337885e-10, 2.338527e-10, 2.336747e-10, 2.348791e-10, 
    2.344432e-10, 2.356163e-10, 2.352992e-10, 2.358183e-10, 2.355605e-10, 
    2.355227e-10, 2.351911e-10, 2.349849e-10, 2.344634e-10, 2.340383e-10, 
    2.337004e-10, 2.337789e-10, 2.3415e-10, 2.348206e-10, 2.354534e-10, 
    2.35315e-10, 2.357788e-10, 2.345481e-10, 2.350652e-10, 2.348658e-10, 
    2.353853e-10, 2.342449e-10, 2.3522e-10, 2.339959e-10, 2.34103e-10, 
    2.344345e-10, 2.351011e-10, 2.352465e-10, 2.354041e-10, 2.353066e-10, 
    2.348374e-10, 2.3476e-10, 2.344261e-10, 2.343346e-10, 2.340796e-10, 
    2.338691e-10, 2.340618e-10, 2.342643e-10, 2.348371e-10, 2.353534e-10, 
    2.359153e-10, 2.360522e-10, 2.367108e-10, 2.361765e-10, 2.370597e-10, 
    2.363115e-10, 2.376046e-10, 2.352745e-10, 2.36287e-10, 2.344492e-10, 
    2.346472e-10, 2.350065e-10, 2.358269e-10, 2.353828e-10, 2.359015e-10, 
    2.347568e-10, 2.341634e-10, 2.340083e-10, 2.337212e-10, 2.340148e-10, 
    2.339909e-10, 2.342718e-10, 2.341815e-10, 2.348561e-10, 2.344938e-10, 
    2.35522e-10, 2.358971e-10, 2.369531e-10, 2.376001e-10, 2.382557e-10, 
    2.385455e-10, 2.386336e-10, 2.386705e-10,
  1.287137e-13, 1.291628e-13, 1.290753e-13, 1.29438e-13, 1.292365e-13, 
    1.294742e-13, 1.288044e-13, 1.29181e-13, 1.289404e-13, 1.287537e-13, 
    1.301449e-13, 1.29454e-13, 1.308606e-13, 1.304197e-13, 1.315261e-13, 
    1.307925e-13, 1.316764e-13, 1.315042e-13, 1.320248e-13, 1.31875e-13, 
    1.325453e-13, 1.320939e-13, 1.328913e-13, 1.32437e-13, 1.325084e-13, 
    1.320792e-13, 1.295919e-13, 1.30059e-13, 1.295645e-13, 1.296308e-13, 
    1.296009e-13, 1.292409e-13, 1.290601e-13, 1.286789e-13, 1.287479e-13, 
    1.290276e-13, 1.296606e-13, 1.294452e-13, 1.299879e-13, 1.299756e-13, 
    1.305819e-13, 1.303086e-13, 1.313268e-13, 1.310373e-13, 1.318813e-13, 
    1.316654e-13, 1.318712e-13, 1.318087e-13, 1.318721e-13, 1.315561e-13, 
    1.316912e-13, 1.314168e-13, 1.303599e-13, 1.306708e-13, 1.297439e-13, 
    1.291905e-13, 1.288211e-13, 1.285595e-13, 1.285965e-13, 1.286672e-13, 
    1.290293e-13, 1.293691e-13, 1.296282e-13, 1.298021e-13, 1.299739e-13, 
    1.304957e-13, 1.307701e-13, 1.313858e-13, 1.31274e-13, 1.314628e-13, 
    1.316439e-13, 1.319543e-13, 1.319031e-13, 1.3204e-13, 1.314574e-13, 
    1.318437e-13, 1.312105e-13, 1.313819e-13, 1.300232e-13, 1.295032e-13, 
    1.292851e-13, 1.290922e-13, 1.28625e-13, 1.289478e-13, 1.288206e-13, 
    1.291227e-13, 1.29315e-13, 1.292198e-13, 1.298069e-13, 1.295784e-13, 
    1.307864e-13, 1.302658e-13, 1.316224e-13, 1.312969e-13, 1.317022e-13, 
    1.314937e-13, 1.318529e-13, 1.315289e-13, 1.320907e-13, 1.322136e-13, 
    1.321297e-13, 1.324513e-13, 1.315114e-13, 1.318715e-13, 1.292172e-13, 
    1.292328e-13, 1.293049e-13, 1.289879e-13, 1.289684e-13, 1.286771e-13, 
    1.28936e-13, 1.290465e-13, 1.293259e-13, 1.294917e-13, 1.29649e-13, 
    1.299965e-13, 1.303854e-13, 1.309284e-13, 1.31318e-13, 1.315792e-13, 
    1.314188e-13, 1.315604e-13, 1.314022e-13, 1.31328e-13, 1.321678e-13, 
    1.316926e-13, 1.32405e-13, 1.323655e-13, 1.320433e-13, 1.3237e-13, 
    1.292436e-13, 1.291543e-13, 1.288448e-13, 1.29087e-13, 1.286454e-13, 
    1.288929e-13, 1.290354e-13, 1.295838e-13, 1.297036e-13, 1.298161e-13, 
    1.300378e-13, 1.303226e-13, 1.308223e-13, 1.312566e-13, 1.316545e-13, 
    1.316247e-13, 1.316352e-13, 1.317263e-13, 1.315031e-13, 1.317633e-13, 
    1.318076e-13, 1.316922e-13, 1.323602e-13, 1.321694e-13, 1.323647e-13, 
    1.322403e-13, 1.291832e-13, 1.293335e-13, 1.292523e-13, 1.294051e-13, 
    1.292977e-13, 1.297763e-13, 1.299205e-13, 1.305943e-13, 1.303171e-13, 
    1.307575e-13, 1.303617e-13, 1.30432e-13, 1.30773e-13, 1.303829e-13, 
    1.312331e-13, 1.306577e-13, 1.317299e-13, 1.311525e-13, 1.317669e-13, 
    1.316527e-13, 1.318414e-13, 1.320106e-13, 1.32223e-13, 1.326157e-13, 
    1.325247e-13, 1.328526e-13, 1.295573e-13, 1.297526e-13, 1.297348e-13, 
    1.299397e-13, 1.300914e-13, 1.304195e-13, 1.309462e-13, 1.30748e-13, 
    1.311113e-13, 1.311845e-13, 1.306321e-13, 1.309718e-13, 1.298835e-13, 
    1.300598e-13, 1.299545e-13, 1.295729e-13, 1.307944e-13, 1.301675e-13, 
    1.313245e-13, 1.309849e-13, 1.319866e-13, 1.314836e-13, 1.324747e-13, 
    1.329008e-13, 1.332993e-13, 1.337677e-13, 1.298591e-13, 1.297258e-13, 
    1.29964e-13, 1.302943e-13, 1.305994e-13, 1.310057e-13, 1.31047e-13, 
    1.311232e-13, 1.313201e-13, 1.314859e-13, 1.311478e-13, 1.315274e-13, 
    1.301017e-13, 1.308486e-13, 1.296761e-13, 1.300297e-13, 1.302746e-13, 
    1.301667e-13, 1.307252e-13, 1.30857e-13, 1.313927e-13, 1.311155e-13, 
    1.327961e-13, 1.320471e-13, 1.341226e-13, 1.335431e-13, 1.296796e-13, 
    1.298584e-13, 1.30482e-13, 1.301852e-13, 1.310325e-13, 1.312413e-13, 
    1.314105e-13, 1.316289e-13, 1.316527e-13, 1.317848e-13, 1.315687e-13, 
    1.31776e-13, 1.310065e-13, 1.31348e-13, 1.304101e-13, 1.306387e-13, 
    1.305334e-13, 1.304182e-13, 1.307737e-13, 1.311533e-13, 1.311606e-13, 
    1.312824e-13, 1.316283e-13, 1.310359e-13, 1.328943e-13, 1.31739e-13, 
    1.300536e-13, 1.303994e-13, 1.304478e-13, 1.30314e-13, 1.312204e-13, 
    1.308921e-13, 1.317814e-13, 1.31537e-13, 1.31938e-13, 1.317382e-13, 
    1.317089e-13, 1.314555e-13, 1.313001e-13, 1.309073e-13, 1.305874e-13, 
    1.303333e-13, 1.303924e-13, 1.306714e-13, 1.311763e-13, 1.316552e-13, 
    1.315489e-13, 1.319074e-13, 1.309711e-13, 1.313606e-13, 1.312103e-13, 
    1.316025e-13, 1.307429e-13, 1.314769e-13, 1.305556e-13, 1.306362e-13, 
    1.308856e-13, 1.313875e-13, 1.314973e-13, 1.31617e-13, 1.315426e-13, 
    1.31189e-13, 1.311306e-13, 1.308793e-13, 1.308103e-13, 1.306186e-13, 
    1.304602e-13, 1.306051e-13, 1.307575e-13, 1.311888e-13, 1.315778e-13, 
    1.320132e-13, 1.321194e-13, 1.326301e-13, 1.322155e-13, 1.329008e-13, 
    1.323199e-13, 1.333246e-13, 1.315182e-13, 1.323012e-13, 1.308967e-13, 
    1.310458e-13, 1.313163e-13, 1.319445e-13, 1.316006e-13, 1.320024e-13, 
    1.311283e-13, 1.306815e-13, 1.305649e-13, 1.303489e-13, 1.305698e-13, 
    1.305518e-13, 1.307632e-13, 1.306952e-13, 1.312031e-13, 1.309303e-13, 
    1.317084e-13, 1.31999e-13, 1.328185e-13, 1.333213e-13, 1.338316e-13, 
    1.340573e-13, 1.341259e-13, 1.341547e-13,
  1.866553e-17, 1.87402e-17, 1.872566e-17, 1.878598e-17, 1.875247e-17, 
    1.879201e-17, 1.868062e-17, 1.874321e-17, 1.870322e-17, 1.867219e-17, 
    1.89034e-17, 1.878865e-17, 1.902236e-17, 1.89491e-17, 1.913309e-17, 
    1.901102e-17, 1.915876e-17, 1.912946e-17, 1.921898e-17, 1.919309e-17, 
    1.930895e-17, 1.923094e-17, 1.936888e-17, 1.929025e-17, 1.930259e-17, 
    1.922838e-17, 1.881161e-17, 1.888913e-17, 1.880705e-17, 1.881808e-17, 
    1.881311e-17, 1.87532e-17, 1.87231e-17, 1.865976e-17, 1.867123e-17, 
    1.871771e-17, 1.882304e-17, 1.87872e-17, 1.887741e-17, 1.887537e-17, 
    1.897605e-17, 1.893064e-17, 1.909994e-17, 1.905177e-17, 1.919417e-17, 
    1.915688e-17, 1.919244e-17, 1.918164e-17, 1.919258e-17, 1.913811e-17, 
    1.916132e-17, 1.911491e-17, 1.893917e-17, 1.899082e-17, 1.883691e-17, 
    1.874478e-17, 1.868338e-17, 1.863992e-17, 1.864607e-17, 1.86578e-17, 
    1.871799e-17, 1.877453e-17, 1.881767e-17, 1.884658e-17, 1.887508e-17, 
    1.896168e-17, 1.900731e-17, 1.910974e-17, 1.909115e-17, 1.912257e-17, 
    1.915316e-17, 1.920678e-17, 1.919794e-17, 1.922159e-17, 1.912167e-17, 
    1.918767e-17, 1.908059e-17, 1.91091e-17, 1.888319e-17, 1.879685e-17, 
    1.876053e-17, 1.872846e-17, 1.86508e-17, 1.870445e-17, 1.86833e-17, 
    1.873354e-17, 1.876553e-17, 1.874969e-17, 1.884737e-17, 1.880938e-17, 
    1.901002e-17, 1.892352e-17, 1.914945e-17, 1.909496e-17, 1.916323e-17, 
    1.912772e-17, 1.918925e-17, 1.913358e-17, 1.923037e-17, 1.925161e-17, 
    1.92371e-17, 1.929273e-17, 1.913066e-17, 1.919247e-17, 1.874926e-17, 
    1.875185e-17, 1.876385e-17, 1.871111e-17, 1.870787e-17, 1.865946e-17, 
    1.87025e-17, 1.872086e-17, 1.876735e-17, 1.879493e-17, 1.882113e-17, 
    1.887883e-17, 1.894339e-17, 1.903364e-17, 1.909846e-17, 1.914199e-17, 
    1.911526e-17, 1.913883e-17, 1.91125e-17, 1.910014e-17, 1.924368e-17, 
    1.916156e-17, 1.928473e-17, 1.92779e-17, 1.922217e-17, 1.927867e-17, 
    1.875366e-17, 1.873879e-17, 1.868733e-17, 1.87276e-17, 1.865419e-17, 
    1.869532e-17, 1.8719e-17, 1.881025e-17, 1.883022e-17, 1.884889e-17, 
    1.888568e-17, 1.893297e-17, 1.9016e-17, 1.908824e-17, 1.9155e-17, 
    1.914984e-17, 1.915166e-17, 1.91674e-17, 1.912928e-17, 1.917379e-17, 
    1.918144e-17, 1.916151e-17, 1.927698e-17, 1.924397e-17, 1.927775e-17, 
    1.925625e-17, 1.874361e-17, 1.876861e-17, 1.875511e-17, 1.878052e-17, 
    1.876264e-17, 1.884227e-17, 1.886619e-17, 1.897809e-17, 1.893206e-17, 
    1.900523e-17, 1.893946e-17, 1.895113e-17, 1.900777e-17, 1.894299e-17, 
    1.908433e-17, 1.898862e-17, 1.916801e-17, 1.907089e-17, 1.91744e-17, 
    1.91547e-17, 1.918729e-17, 1.921653e-17, 1.925325e-17, 1.932117e-17, 
    1.930542e-17, 1.936219e-17, 1.880585e-17, 1.883834e-17, 1.883541e-17, 
    1.886941e-17, 1.889458e-17, 1.894907e-17, 1.903662e-17, 1.900367e-17, 
    1.906409e-17, 1.907625e-17, 1.898441e-17, 1.904086e-17, 1.886006e-17, 
    1.888932e-17, 1.887185e-17, 1.880845e-17, 1.901135e-17, 1.890719e-17, 
    1.909955e-17, 1.904304e-17, 1.921237e-17, 1.912601e-17, 1.929677e-17, 
    1.937049e-17, 1.943959e-17, 1.952078e-17, 1.885602e-17, 1.883392e-17, 
    1.887343e-17, 1.892825e-17, 1.897895e-17, 1.904651e-17, 1.905338e-17, 
    1.906606e-17, 1.909883e-17, 1.912642e-17, 1.907014e-17, 1.913334e-17, 
    1.889624e-17, 1.902037e-17, 1.882564e-17, 1.888432e-17, 1.892499e-17, 
    1.890708e-17, 1.899988e-17, 1.902179e-17, 1.91109e-17, 1.906479e-17, 
    1.935236e-17, 1.92228e-17, 1.958241e-17, 1.948183e-17, 1.882623e-17, 
    1.885591e-17, 1.895943e-17, 1.891015e-17, 1.905098e-17, 1.90857e-17, 
    1.911388e-17, 1.915057e-17, 1.915468e-17, 1.917749e-17, 1.914021e-17, 
    1.917599e-17, 1.904665e-17, 1.910347e-17, 1.894751e-17, 1.898549e-17, 
    1.896799e-17, 1.894886e-17, 1.900794e-17, 1.907104e-17, 1.907228e-17, 
    1.909254e-17, 1.915038e-17, 1.905155e-17, 1.93693e-17, 1.91695e-17, 
    1.888831e-17, 1.894571e-17, 1.895377e-17, 1.893156e-17, 1.908222e-17, 
    1.902762e-17, 1.917692e-17, 1.913494e-17, 1.920398e-17, 1.916946e-17, 
    1.916439e-17, 1.912137e-17, 1.90955e-17, 1.903014e-17, 1.897697e-17, 
    1.893476e-17, 1.894457e-17, 1.899093e-17, 1.907488e-17, 1.91551e-17, 
    1.913689e-17, 1.919869e-17, 1.904076e-17, 1.910555e-17, 1.908054e-17, 
    1.914601e-17, 1.900281e-17, 1.912485e-17, 1.897169e-17, 1.898508e-17, 
    1.902654e-17, 1.911002e-17, 1.912833e-17, 1.914851e-17, 1.913587e-17, 
    1.907699e-17, 1.906729e-17, 1.90255e-17, 1.901402e-17, 1.898216e-17, 
    1.895584e-17, 1.897991e-17, 1.900522e-17, 1.907697e-17, 1.914175e-17, 
    1.921696e-17, 1.923534e-17, 1.932362e-17, 1.925191e-17, 1.937044e-17, 
    1.926989e-17, 1.944389e-17, 1.913176e-17, 1.926671e-17, 1.902839e-17, 
    1.905318e-17, 1.909816e-17, 1.920506e-17, 1.914568e-17, 1.921507e-17, 
    1.906691e-17, 1.899258e-17, 1.897323e-17, 1.893735e-17, 1.897405e-17, 
    1.897106e-17, 1.900619e-17, 1.899489e-17, 1.907935e-17, 1.903397e-17, 
    1.916429e-17, 1.92145e-17, 1.935628e-17, 1.944337e-17, 1.953191e-17, 
    1.957109e-17, 1.9583e-17, 1.958799e-17,
  7.810657e-22, 7.846024e-22, 7.839133e-22, 7.86772e-22, 7.851841e-22, 
    7.87058e-22, 7.817803e-22, 7.847445e-22, 7.828506e-22, 7.813813e-22, 
    7.923391e-22, 7.868991e-22, 7.979898e-22, 7.945105e-22, 8.032567e-22, 
    7.974503e-22, 8.044773e-22, 8.030847e-22, 8.0734e-22, 8.061096e-22, 
    8.116348e-22, 8.079081e-22, 8.145784e-22, 8.107283e-22, 8.113233e-22, 
    8.077865e-22, 7.879883e-22, 7.916622e-22, 7.877719e-22, 7.882949e-22, 
    7.880593e-22, 7.852183e-22, 7.83791e-22, 7.807929e-22, 7.813361e-22, 
    7.835367e-22, 7.8853e-22, 7.868308e-22, 7.911091e-22, 7.910123e-22, 
    7.957903e-22, 7.936346e-22, 8.0168e-22, 7.99389e-22, 8.061608e-22, 
    8.04389e-22, 8.060783e-22, 8.055654e-22, 8.06085e-22, 8.034966e-22, 
    8.045999e-22, 8.023926e-22, 7.94039e-22, 7.964917e-22, 7.89188e-22, 
    7.848179e-22, 7.81911e-22, 7.798541e-22, 7.801448e-22, 7.806998e-22, 
    7.835497e-22, 7.862297e-22, 7.88276e-22, 7.896469e-22, 7.909984e-22, 
    7.951061e-22, 7.972745e-22, 8.021456e-22, 8.012621e-22, 8.027563e-22, 
    8.042127e-22, 8.067598e-22, 8.063397e-22, 8.074636e-22, 8.027142e-22, 
    8.05851e-22, 8.007598e-22, 8.021161e-22, 7.913802e-22, 7.872884e-22, 
    7.855645e-22, 7.840463e-22, 7.803685e-22, 7.829083e-22, 7.81907e-22, 
    7.84287e-22, 7.85803e-22, 7.850525e-22, 7.896843e-22, 7.878826e-22, 
    7.974032e-22, 7.932961e-22, 8.040362e-22, 8.01443e-22, 8.046909e-22, 
    8.030022e-22, 8.059267e-22, 8.03281e-22, 8.078809e-22, 8.088907e-22, 
    8.082008e-22, 8.108469e-22, 8.031423e-22, 8.060797e-22, 7.850321e-22, 
    7.851546e-22, 7.857236e-22, 7.83224e-22, 7.830704e-22, 7.807787e-22, 
    7.828164e-22, 7.83686e-22, 7.858897e-22, 7.871972e-22, 7.884399e-22, 
    7.91176e-22, 7.94239e-22, 7.985262e-22, 8.016098e-22, 8.036821e-22, 
    8.024094e-22, 8.035312e-22, 8.022777e-22, 8.016898e-22, 8.085132e-22, 
    8.046111e-22, 8.104661e-22, 8.101412e-22, 8.074909e-22, 8.101778e-22, 
    7.852403e-22, 7.845361e-22, 7.820978e-22, 7.840057e-22, 7.805291e-22, 
    7.824761e-22, 7.835975e-22, 7.879233e-22, 7.888717e-22, 7.897562e-22, 
    7.915013e-22, 7.93745e-22, 7.97688e-22, 8.011231e-22, 8.043001e-22, 
    8.040552e-22, 8.041415e-22, 8.048889e-22, 8.030763e-22, 8.051924e-22, 
    8.055553e-22, 8.046089e-22, 8.100977e-22, 8.085279e-22, 8.101342e-22, 
    8.091116e-22, 7.847646e-22, 7.859492e-22, 7.853092e-22, 7.865137e-22, 
    7.856661e-22, 7.894417e-22, 7.905756e-22, 7.958865e-22, 7.937016e-22, 
    7.971761e-22, 7.940531e-22, 7.946069e-22, 7.972956e-22, 7.942208e-22, 
    8.009362e-22, 7.963862e-22, 8.04918e-22, 8.002964e-22, 8.052215e-22, 
    8.042857e-22, 8.058338e-22, 8.072229e-22, 8.089692e-22, 8.122357e-22, 
    8.114631e-22, 8.142501e-22, 7.877153e-22, 7.892557e-22, 7.891174e-22, 
    7.907294e-22, 7.919231e-22, 7.945096e-22, 7.986683e-22, 7.971025e-22, 
    7.99975e-22, 8.005531e-22, 7.961878e-22, 7.988695e-22, 7.902857e-22, 
    7.916727e-22, 7.908448e-22, 7.878382e-22, 7.974669e-22, 7.925207e-22, 
    8.016613e-22, 7.98974e-22, 8.070252e-22, 8.0292e-22, 8.110388e-22, 
    8.146564e-22, 8.180542e-22, 8.220476e-22, 7.900944e-22, 7.89047e-22, 
    7.909204e-22, 7.935204e-22, 7.959283e-22, 7.991383e-22, 7.994655e-22, 
    8.000684e-22, 8.016274e-22, 8.029405e-22, 8.002616e-22, 8.032695e-22, 
    7.919998e-22, 7.978956e-22, 7.886537e-22, 7.914355e-22, 7.933658e-22, 
    7.925161e-22, 7.969229e-22, 7.97964e-22, 8.02201e-22, 8.000081e-22, 
    8.137653e-22, 8.075203e-22, 8.25084e-22, 8.20131e-22, 7.886819e-22, 
    7.900895e-22, 7.950009e-22, 7.92662e-22, 7.993513e-22, 8.010026e-22, 
    8.023436e-22, 8.040892e-22, 8.042846e-22, 8.05368e-22, 8.035967e-22, 
    8.052968e-22, 7.991451e-22, 8.018482e-22, 7.944356e-22, 7.962388e-22, 
    7.954082e-22, 7.944995e-22, 7.973058e-22, 8.003045e-22, 8.003642e-22, 
    8.013275e-22, 8.040766e-22, 7.993783e-22, 8.145954e-22, 8.049852e-22, 
    7.91626e-22, 7.943485e-22, 7.947325e-22, 7.936781e-22, 8.008372e-22, 
    7.982407e-22, 8.053409e-22, 8.03346e-22, 8.066268e-22, 8.049866e-22, 
    8.047457e-22, 8.027e-22, 8.014687e-22, 7.983605e-22, 7.958339e-22, 
    7.938305e-22, 7.942958e-22, 7.96497e-22, 8.00487e-22, 8.043043e-22, 
    8.03438e-22, 8.063757e-22, 7.988657e-22, 8.019464e-22, 8.007565e-22, 
    8.038727e-22, 7.970618e-22, 8.028622e-22, 7.955835e-22, 7.962197e-22, 
    7.981892e-22, 8.021584e-22, 8.030312e-22, 8.039913e-22, 8.033903e-22, 
    8.005876e-22, 8.001269e-22, 7.981402e-22, 7.975942e-22, 7.960808e-22, 
    7.948309e-22, 7.95974e-22, 7.97176e-22, 8.00587e-22, 8.036697e-22, 
    8.072434e-22, 8.081172e-22, 8.12354e-22, 8.089032e-22, 8.14651e-22, 
    8.097562e-22, 8.182624e-22, 8.031924e-22, 8.096067e-22, 7.982774e-22, 
    7.994561e-22, 8.015946e-22, 8.066768e-22, 8.038571e-22, 8.07153e-22, 
    8.001085e-22, 7.965751e-22, 7.956567e-22, 7.93953e-22, 7.956956e-22, 
    7.955537e-22, 7.972228e-22, 7.96686e-22, 8.007003e-22, 7.985428e-22, 
    8.047408e-22, 8.071258e-22, 8.139595e-22, 8.182389e-22, 8.225973e-22, 
    8.245267e-22, 8.251139e-22, 8.253597e-22,
  1.00588e-26, 1.011082e-26, 1.010068e-26, 1.014275e-26, 1.011938e-26, 
    1.014696e-26, 1.006931e-26, 1.01129e-26, 1.008505e-26, 1.006345e-26, 
    1.022478e-26, 1.014463e-26, 1.030824e-26, 1.025685e-26, 1.038616e-26, 
    1.030026e-26, 1.040401e-26, 1.038362e-26, 1.044562e-26, 1.042773e-26, 
    1.050818e-26, 1.045388e-26, 1.055155e-26, 1.049489e-26, 1.05036e-26, 
    1.045211e-26, 1.016068e-26, 1.021479e-26, 1.015749e-26, 1.016519e-26, 
    1.016172e-26, 1.011988e-26, 1.009887e-26, 1.00548e-26, 1.006278e-26, 
    1.009514e-26, 1.016865e-26, 1.014363e-26, 1.020668e-26, 1.020525e-26, 
    1.027575e-26, 1.024393e-26, 1.036283e-26, 1.032894e-26, 1.042848e-26, 
    1.040273e-26, 1.042728e-26, 1.041982e-26, 1.042737e-26, 1.038972e-26, 
    1.040579e-26, 1.037338e-26, 1.024989e-26, 1.028611e-26, 1.017835e-26, 
    1.011397e-26, 1.007123e-26, 1.004101e-26, 1.004528e-26, 1.005343e-26, 
    1.009533e-26, 1.013478e-26, 1.016492e-26, 1.018512e-26, 1.020504e-26, 
    1.026562e-26, 1.029767e-26, 1.036971e-26, 1.035665e-26, 1.037875e-26, 
    1.040017e-26, 1.043718e-26, 1.043108e-26, 1.044741e-26, 1.037814e-26, 
    1.042397e-26, 1.034922e-26, 1.036929e-26, 1.021063e-26, 1.015037e-26, 
    1.012496e-26, 1.010263e-26, 1.004856e-26, 1.008589e-26, 1.007117e-26, 
    1.010618e-26, 1.012849e-26, 1.011745e-26, 1.018567e-26, 1.015912e-26, 
    1.029957e-26, 1.023893e-26, 1.039761e-26, 1.035932e-26, 1.040712e-26, 
    1.038241e-26, 1.042507e-26, 1.038653e-26, 1.045348e-26, 1.046816e-26, 
    1.045813e-26, 1.049663e-26, 1.038448e-26, 1.042729e-26, 1.011715e-26, 
    1.011895e-26, 1.012733e-26, 1.009054e-26, 1.008828e-26, 1.005459e-26, 
    1.008455e-26, 1.009733e-26, 1.012977e-26, 1.014902e-26, 1.016733e-26, 
    1.020766e-26, 1.025284e-26, 1.031617e-26, 1.036179e-26, 1.039247e-26, 
    1.037363e-26, 1.039024e-26, 1.037168e-26, 1.036298e-26, 1.046267e-26, 
    1.040595e-26, 1.049109e-26, 1.048636e-26, 1.044781e-26, 1.048689e-26, 
    1.012021e-26, 1.010985e-26, 1.007398e-26, 1.010204e-26, 1.005092e-26, 
    1.007954e-26, 1.009603e-26, 1.015971e-26, 1.01737e-26, 1.018673e-26, 
    1.021246e-26, 1.024556e-26, 1.030378e-26, 1.035458e-26, 1.040144e-26, 
    1.039789e-26, 1.039914e-26, 1.040999e-26, 1.03835e-26, 1.04144e-26, 
    1.041967e-26, 1.040593e-26, 1.048573e-26, 1.046289e-26, 1.048626e-26, 
    1.047138e-26, 1.011321e-26, 1.013065e-26, 1.012123e-26, 1.013895e-26, 
    1.012648e-26, 1.018208e-26, 1.019879e-26, 1.027716e-26, 1.024491e-26, 
    1.029622e-26, 1.02501e-26, 1.025828e-26, 1.029797e-26, 1.025258e-26, 
    1.035181e-26, 1.028454e-26, 1.041042e-26, 1.034234e-26, 1.041483e-26, 
    1.040123e-26, 1.042373e-26, 1.044391e-26, 1.046931e-26, 1.051704e-26, 
    1.050566e-26, 1.054672e-26, 1.015666e-26, 1.017935e-26, 1.017732e-26, 
    1.020108e-26, 1.021867e-26, 1.025684e-26, 1.031828e-26, 1.029514e-26, 
    1.033761e-26, 1.034615e-26, 1.028163e-26, 1.032125e-26, 1.019453e-26, 
    1.021497e-26, 1.020277e-26, 1.015846e-26, 1.030051e-26, 1.022748e-26, 
    1.036255e-26, 1.03228e-26, 1.044104e-26, 1.038118e-26, 1.049942e-26, 
    1.055269e-26, 1.060411e-26, 1.066479e-26, 1.019171e-26, 1.017628e-26, 
    1.020389e-26, 1.024223e-26, 1.027779e-26, 1.032523e-26, 1.033007e-26, 
    1.033898e-26, 1.036205e-26, 1.038149e-26, 1.034183e-26, 1.038636e-26, 
    1.021978e-26, 1.030685e-26, 1.017048e-26, 1.021147e-26, 1.023995e-26, 
    1.022742e-26, 1.029249e-26, 1.030787e-26, 1.037054e-26, 1.03381e-26, 
    1.053955e-26, 1.044822e-26, 1.071102e-26, 1.063565e-26, 1.01709e-26, 
    1.019164e-26, 1.026409e-26, 1.022958e-26, 1.032838e-26, 1.03528e-26, 
    1.037266e-26, 1.039837e-26, 1.040122e-26, 1.041695e-26, 1.039121e-26, 
    1.041592e-26, 1.032533e-26, 1.036532e-26, 1.025575e-26, 1.028238e-26, 
    1.027011e-26, 1.02567e-26, 1.029814e-26, 1.034247e-26, 1.034336e-26, 
    1.035761e-26, 1.039815e-26, 1.032878e-26, 1.055176e-26, 1.041136e-26, 
    1.02143e-26, 1.025445e-26, 1.026013e-26, 1.024457e-26, 1.035036e-26, 
    1.031196e-26, 1.041656e-26, 1.03875e-26, 1.043525e-26, 1.041142e-26, 
    1.040791e-26, 1.037793e-26, 1.03597e-26, 1.031373e-26, 1.027639e-26, 
    1.024682e-26, 1.025369e-26, 1.028619e-26, 1.034517e-26, 1.04015e-26, 
    1.038885e-26, 1.04316e-26, 1.03212e-26, 1.036677e-26, 1.034916e-26, 
    1.039523e-26, 1.029454e-26, 1.038029e-26, 1.02727e-26, 1.02821e-26, 
    1.03112e-26, 1.03699e-26, 1.038283e-26, 1.039695e-26, 1.038815e-26, 
    1.034666e-26, 1.033985e-26, 1.031048e-26, 1.03024e-26, 1.028005e-26, 
    1.026159e-26, 1.027847e-26, 1.029622e-26, 1.034666e-26, 1.039228e-26, 
    1.044421e-26, 1.045692e-26, 1.051876e-26, 1.046833e-26, 1.055258e-26, 
    1.048071e-26, 1.060723e-26, 1.03852e-26, 1.047855e-26, 1.03125e-26, 
    1.032993e-26, 1.036155e-26, 1.043596e-26, 1.039501e-26, 1.044289e-26, 
    1.033958e-26, 1.028734e-26, 1.027378e-26, 1.024863e-26, 1.027436e-26, 
    1.027226e-26, 1.029692e-26, 1.028899e-26, 1.034833e-26, 1.031643e-26, 
    1.040784e-26, 1.044249e-26, 1.054243e-26, 1.06069e-26, 1.067318e-26, 
    1.070254e-26, 1.071149e-26, 1.071523e-26,
  4.063426e-32, 4.088648e-32, 4.083731e-32, 4.104154e-32, 4.092808e-32, 
    4.106201e-32, 4.068521e-32, 4.089659e-32, 4.07615e-32, 4.065681e-32, 
    4.144518e-32, 4.105065e-32, 4.186438e-32, 4.160626e-32, 4.225689e-32, 
    4.182424e-32, 4.234591e-32, 4.224417e-32, 4.255249e-32, 4.246369e-32, 
    4.286296e-32, 4.259353e-32, 4.307672e-32, 4.279739e-32, 4.284045e-32, 
    4.258473e-32, 4.112869e-32, 4.139514e-32, 4.111319e-32, 4.11506e-32, 
    4.113377e-32, 4.093049e-32, 4.082846e-32, 4.061491e-32, 4.065358e-32, 
    4.08104e-32, 4.116743e-32, 4.104584e-32, 4.135468e-32, 4.134752e-32, 
    4.170116e-32, 4.154142e-32, 4.213931e-32, 4.196864e-32, 4.246739e-32, 
    4.233965e-32, 4.246141e-32, 4.242444e-32, 4.246189e-32, 4.227493e-32, 
    4.235482e-32, 4.219251e-32, 4.157133e-32, 4.175318e-32, 4.121462e-32, 
    4.090172e-32, 4.06945e-32, 4.054809e-32, 4.056877e-32, 4.060823e-32, 
    4.081132e-32, 4.100284e-32, 4.114933e-32, 4.124758e-32, 4.13465e-32, 
    4.165018e-32, 4.181123e-32, 4.217398e-32, 4.210818e-32, 4.221958e-32, 
    4.232695e-32, 4.251057e-32, 4.248028e-32, 4.256137e-32, 4.221652e-32, 
    4.244497e-32, 4.207077e-32, 4.217187e-32, 4.137427e-32, 4.107859e-32, 
    4.095509e-32, 4.084678e-32, 4.058468e-32, 4.076557e-32, 4.06942e-32, 
    4.086403e-32, 4.097232e-32, 4.091871e-32, 4.125027e-32, 4.112113e-32, 
    4.18208e-32, 4.151629e-32, 4.231424e-32, 4.212166e-32, 4.236141e-32, 
    4.223805e-32, 4.245045e-32, 4.225888e-32, 4.259153e-32, 4.266445e-32, 
    4.261462e-32, 4.280606e-32, 4.22485e-32, 4.246147e-32, 4.091723e-32, 
    4.092598e-32, 4.096666e-32, 4.078808e-32, 4.077714e-32, 4.061388e-32, 
    4.075907e-32, 4.082107e-32, 4.097856e-32, 4.107205e-32, 4.116105e-32, 
    4.135957e-32, 4.158609e-32, 4.190434e-32, 4.213409e-32, 4.228876e-32, 
    4.21938e-32, 4.227757e-32, 4.218395e-32, 4.214011e-32, 4.263715e-32, 
    4.23556e-32, 4.277848e-32, 4.275497e-32, 4.256332e-32, 4.275762e-32, 
    4.093211e-32, 4.088183e-32, 4.070782e-32, 4.084394e-32, 4.059613e-32, 
    4.073477e-32, 4.081471e-32, 4.112396e-32, 4.119201e-32, 4.125538e-32, 
    4.138363e-32, 4.154958e-32, 4.184204e-32, 4.209775e-32, 4.233327e-32, 
    4.231564e-32, 4.232186e-32, 4.237566e-32, 4.224356e-32, 4.239754e-32, 
    4.242365e-32, 4.235549e-32, 4.275183e-32, 4.26383e-32, 4.275448e-32, 
    4.268051e-32, 4.089815e-32, 4.098278e-32, 4.093704e-32, 4.102312e-32, 
    4.096251e-32, 4.123274e-32, 4.131511e-32, 4.170819e-32, 4.154635e-32, 
    4.180399e-32, 4.157241e-32, 4.161341e-32, 4.181267e-32, 4.158486e-32, 
    4.208374e-32, 4.174522e-32, 4.237776e-32, 4.203596e-32, 4.239963e-32, 
    4.233223e-32, 4.244381e-32, 4.2544e-32, 4.267019e-32, 4.290665e-32, 
    4.285067e-32, 4.305293e-32, 4.110916e-32, 4.121946e-32, 4.120963e-32, 
    4.132661e-32, 4.141478e-32, 4.160624e-32, 4.191496e-32, 4.179862e-32, 
    4.201228e-32, 4.205531e-32, 4.173072e-32, 4.192989e-32, 4.12938e-32, 
    4.139616e-32, 4.13351e-32, 4.111792e-32, 4.182556e-32, 4.145887e-32, 
    4.213792e-32, 4.193772e-32, 4.252972e-32, 4.223179e-32, 4.281992e-32, 
    4.308227e-32, 4.333833e-32, 4.364129e-32, 4.127971e-32, 4.120459e-32, 
    4.134074e-32, 4.153285e-32, 4.171141e-32, 4.194994e-32, 4.197434e-32, 
    4.20192e-32, 4.213545e-32, 4.223344e-32, 4.203351e-32, 4.225802e-32, 
    4.142016e-32, 4.185746e-32, 4.117635e-32, 4.137861e-32, 4.152145e-32, 
    4.145862e-32, 4.178531e-32, 4.186265e-32, 4.217814e-32, 4.201474e-32, 
    4.301751e-32, 4.256535e-32, 4.38764e-32, 4.349571e-32, 4.117842e-32, 
    4.127939e-32, 4.164257e-32, 4.146943e-32, 4.196584e-32, 4.208881e-32, 
    4.218889e-32, 4.231802e-32, 4.233214e-32, 4.241017e-32, 4.228246e-32, 
    4.240507e-32, 4.195045e-32, 4.215188e-32, 4.160079e-32, 4.173445e-32, 
    4.167288e-32, 4.160551e-32, 4.181373e-32, 4.203668e-32, 4.204126e-32, 
    4.211299e-32, 4.231669e-32, 4.196785e-32, 4.307756e-32, 4.238221e-32, 
    4.139286e-32, 4.159415e-32, 4.162274e-32, 4.154467e-32, 4.207647e-32, 
    4.188318e-32, 4.240824e-32, 4.226373e-32, 4.2501e-32, 4.238272e-32, 
    4.236535e-32, 4.221548e-32, 4.212358e-32, 4.189206e-32, 4.170439e-32, 
    4.155596e-32, 4.159042e-32, 4.17536e-32, 4.20503e-32, 4.233351e-32, 
    4.227051e-32, 4.248289e-32, 4.192969e-32, 4.215915e-32, 4.207041e-32, 
    4.230247e-32, 4.179557e-32, 4.222716e-32, 4.168589e-32, 4.173308e-32, 
    4.187935e-32, 4.217488e-32, 4.224021e-32, 4.231097e-32, 4.226704e-32, 
    4.205782e-32, 4.202354e-32, 4.187574e-32, 4.18351e-32, 4.172279e-32, 
    4.163008e-32, 4.171482e-32, 4.180401e-32, 4.205783e-32, 4.228778e-32, 
    4.254545e-32, 4.260863e-32, 4.291501e-32, 4.26652e-32, 4.308157e-32, 
    4.272657e-32, 4.33537e-32, 4.2252e-32, 4.271602e-32, 4.188595e-32, 
    4.197364e-32, 4.213284e-32, 4.250444e-32, 4.230135e-32, 4.253884e-32, 
    4.202219e-32, 4.175933e-32, 4.169131e-32, 4.156501e-32, 4.16942e-32, 
    4.168367e-32, 4.180758e-32, 4.176772e-32, 4.206628e-32, 4.190568e-32, 
    4.236496e-32, 4.253691e-32, 4.303177e-32, 4.335217e-32, 4.368331e-32, 
    4.383287e-32, 4.387881e-32, 4.389804e-32,
  5.366372e-38, 5.411483e-38, 5.402676e-38, 5.439307e-38, 5.418946e-38, 
    5.442986e-38, 5.375476e-38, 5.413291e-38, 5.389112e-38, 5.370404e-38, 
    5.512234e-38, 5.440945e-38, 5.588809e-38, 5.541613e-38, 5.662753e-38, 
    5.581448e-38, 5.679534e-38, 5.66035e-38, 5.718431e-38, 5.701696e-38, 
    5.777032e-38, 5.726173e-38, 5.817127e-38, 5.764722e-38, 5.772827e-38, 
    5.724512e-38, 5.454983e-38, 5.50313e-38, 5.452192e-38, 5.458922e-38, 
    5.455897e-38, 5.419373e-38, 5.401082e-38, 5.362927e-38, 5.369828e-38, 
    5.397855e-38, 5.461951e-38, 5.440087e-38, 5.49581e-38, 5.494511e-38, 
    5.558946e-38, 5.529791e-38, 5.640457e-38, 5.608171e-38, 5.702393e-38, 
    5.67837e-38, 5.701266e-38, 5.694309e-38, 5.701357e-38, 5.666192e-38, 
    5.681217e-38, 5.650545e-38, 5.535243e-38, 5.568454e-38, 5.470454e-38, 
    5.414201e-38, 5.377132e-38, 5.35101e-38, 5.354694e-38, 5.361731e-38, 
    5.39802e-38, 5.432363e-38, 5.4587e-38, 5.476399e-38, 5.494324e-38, 
    5.549611e-38, 5.579073e-38, 5.647023e-38, 5.634561e-38, 5.655676e-38, 
    5.675985e-38, 5.710524e-38, 5.704819e-38, 5.7201e-38, 5.655104e-38, 
    5.698166e-38, 5.627482e-38, 5.646631e-38, 5.499335e-38, 5.445972e-38, 
    5.423775e-38, 5.40437e-38, 5.357531e-38, 5.389834e-38, 5.377076e-38, 
    5.407466e-38, 5.426883e-38, 5.417267e-38, 5.476884e-38, 5.453625e-38, 
    5.580824e-38, 5.525207e-38, 5.673597e-38, 5.637115e-38, 5.682458e-38, 
    5.659191e-38, 5.699199e-38, 5.663146e-38, 5.725793e-38, 5.739561e-38, 
    5.73015e-38, 5.766372e-38, 5.661175e-38, 5.701274e-38, 5.417002e-38, 
    5.418569e-38, 5.425869e-38, 5.393861e-38, 5.391906e-38, 5.362741e-38, 
    5.388676e-38, 5.399767e-38, 5.428005e-38, 5.444797e-38, 5.460807e-38, 
    5.496696e-38, 5.537929e-38, 5.59614e-38, 5.639468e-38, 5.668816e-38, 
    5.650793e-38, 5.666697e-38, 5.648924e-38, 5.640613e-38, 5.734403e-38, 
    5.681361e-38, 5.761146e-38, 5.756694e-38, 5.720467e-38, 5.757196e-38, 
    5.419669e-38, 5.410656e-38, 5.379514e-38, 5.403869e-38, 5.359574e-38, 
    5.384329e-38, 5.398624e-38, 5.454126e-38, 5.466385e-38, 5.477803e-38, 
    5.501071e-38, 5.53128e-38, 5.584721e-38, 5.632581e-38, 5.677174e-38, 
    5.673864e-38, 5.67503e-38, 5.685135e-38, 5.660236e-38, 5.689248e-38, 
    5.694156e-38, 5.681346e-38, 5.756099e-38, 5.734626e-38, 5.7566e-38, 
    5.742605e-38, 5.413582e-38, 5.428762e-38, 5.420555e-38, 5.436003e-38, 
    5.42512e-38, 5.473714e-38, 5.488608e-38, 5.56022e-38, 5.530687e-38, 
    5.57775e-38, 5.535442e-38, 5.542917e-38, 5.579325e-38, 5.537715e-38, 
    5.629921e-38, 5.566988e-38, 5.685529e-38, 5.620872e-38, 5.689642e-38, 
    5.676978e-38, 5.697954e-38, 5.716825e-38, 5.740653e-38, 5.785225e-38, 
    5.774748e-38, 5.812665e-38, 5.45147e-38, 5.471325e-38, 5.46956e-38, 
    5.49071e-38, 5.506731e-38, 5.541615e-38, 5.598093e-38, 5.576776e-38, 
    5.616417e-38, 5.624554e-38, 5.564354e-38, 5.600847e-38, 5.484748e-38, 
    5.503336e-38, 5.49225e-38, 5.453042e-38, 5.5817e-38, 5.514745e-38, 
    5.640193e-38, 5.602332e-38, 5.714132e-38, 5.65799e-38, 5.768996e-38, 
    5.818159e-38, 5.865906e-38, 5.9232e-38, 5.482195e-38, 5.468652e-38, 
    5.493278e-38, 5.52822e-38, 5.560819e-38, 5.604636e-38, 5.609248e-38, 
    5.617724e-38, 5.639729e-38, 5.658314e-38, 5.620421e-38, 5.662983e-38, 
    5.507685e-38, 5.587547e-38, 5.46356e-38, 5.500144e-38, 5.526147e-38, 
    5.514709e-38, 5.574341e-38, 5.588504e-38, 5.647814e-38, 5.616884e-38, 
    5.805993e-38, 5.720841e-38, 5.968742e-38, 5.895294e-38, 5.463937e-38, 
    5.482139e-38, 5.548239e-38, 5.516678e-38, 5.607642e-38, 5.630892e-38, 
    5.649861e-38, 5.674304e-38, 5.676961e-38, 5.691622e-38, 5.667628e-38, 
    5.690666e-38, 5.604731e-38, 5.642842e-38, 5.540622e-38, 5.565033e-38, 
    5.553784e-38, 5.541484e-38, 5.579544e-38, 5.621019e-38, 5.621898e-38, 
    5.635468e-38, 5.674013e-38, 5.608023e-38, 5.817247e-38, 5.686327e-38, 
    5.502751e-38, 5.539396e-38, 5.544624e-38, 5.530387e-38, 5.628557e-38, 
    5.592265e-38, 5.69126e-38, 5.664067e-38, 5.708724e-38, 5.686462e-38, 
    5.683197e-38, 5.654906e-38, 5.637477e-38, 5.593892e-38, 5.559536e-38, 
    5.532446e-38, 5.53873e-38, 5.568532e-38, 5.623598e-38, 5.677212e-38, 
    5.665348e-38, 5.705312e-38, 5.600817e-38, 5.644215e-38, 5.627403e-38, 
    5.671388e-38, 5.576215e-38, 5.657084e-38, 5.55616e-38, 5.564785e-38, 
    5.591563e-38, 5.647189e-38, 5.659601e-38, 5.67298e-38, 5.664696e-38, 
    5.625022e-38, 5.618543e-38, 5.590905e-38, 5.583452e-38, 5.562904e-38, 
    5.545967e-38, 5.561446e-38, 5.577758e-38, 5.62503e-38, 5.668627e-38, 
    5.717098e-38, 5.729023e-38, 5.78677e-38, 5.739687e-38, 5.817999e-38, 
    5.751265e-38, 5.868739e-38, 5.661816e-38, 5.749292e-38, 5.592777e-38, 
    5.609118e-38, 5.639223e-38, 5.709355e-38, 5.671178e-38, 5.715843e-38, 
    5.618288e-38, 5.569575e-38, 5.557149e-38, 5.534093e-38, 5.557677e-38, 
    5.555754e-38, 5.578418e-38, 5.571122e-38, 5.626628e-38, 5.596396e-38, 
    5.683121e-38, 5.715482e-38, 5.808686e-38, 5.868474e-38, 5.931324e-38, 
    5.960292e-38, 5.969218e-38, 5.972956e-38,
  2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 3.082857e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  5.018213e-06, 4.75359e-06, 4.804705e-06, 4.593667e-06, 4.710366e-06, 
    4.572701e-06, 4.964221e-06, 4.74319e-06, 4.883953e-06, 4.994195e-06, 
    4.192902e-06, 4.584314e-06, 3.79729e-06, 4.036672e-06, 3.446875e-06, 
    3.83419e-06, 3.370993e-06, 3.457745e-06, 3.199686e-06, 3.272633e-06, 
    2.953456e-06, 3.166293e-06, 2.794725e-06, 3.003558e-06, 2.970367e-06, 
    3.173451e-06, 4.504567e-06, 4.241e-06, 4.52036e-06, 4.482408e-06, 
    4.499412e-06, 4.707966e-06, 4.814172e-06, 5.038557e-06, 4.997606e-06, 
    4.832875e-06, 4.465374e-06, 4.589089e-06, 4.279326e-06, 4.286239e-06, 
    3.947762e-06, 4.097855e-06, 3.549808e-06, 3.702263e-06, 3.269571e-06, 
    3.376075e-06, 3.274546e-06, 3.30517e-06, 3.274148e-06, 3.430997e-06, 
    3.363374e-06, 3.502917e-06, 4.069594e-06, 3.899496e-06, 4.417599e-06, 
    4.738097e-06, 4.954479e-06, 5.109648e-06, 5.087637e-06, 5.045755e-06, 
    4.831918e-06, 4.633222e-06, 4.483531e-06, 4.384293e-06, 4.287235e-06, 
    3.995816e-06, 3.846042e-06, 3.519345e-06, 3.577339e-06, 3.479311e-06, 
    3.386757e-06, 3.234062e-06, 3.258956e-06, 3.192526e-06, 3.481852e-06, 
    3.288245e-06, 3.610569e-06, 3.521056e-06, 4.261162e-06, 4.555599e-06, 
    4.682812e-06, 4.794875e-06, 5.070734e-06, 4.87979e-06, 4.954833e-06, 
    4.776787e-06, 4.664657e-06, 4.720008e-06, 4.381589e-06, 4.512217e-06, 
    3.837236e-06, 4.12182e-06, 3.397492e-06, 3.565398e-06, 3.357794e-06, 
    3.463012e-06, 3.283674e-06, 3.444877e-06, 3.167963e-06, 3.109191e-06, 
    3.149298e-06, 2.996624e-06, 3.453923e-06, 3.274562e-06, 4.721571e-06, 
    4.712531e-06, 4.670459e-06, 4.85622e-06, 4.86764e-06, 5.039691e-06, 
    4.886502e-06, 4.821678e-06, 4.658166e-06, 4.562286e-06, 4.471709e-06, 
    4.274668e-06, 4.055766e-06, 3.760722e-06, 3.554406e-06, 3.418986e-06, 
    3.501731e-06, 3.428633e-06, 3.5104e-06, 3.549016e-06, 3.131157e-06, 
    3.362757e-06, 3.018341e-06, 3.036902e-06, 3.190961e-06, 3.034807e-06, 
    4.706183e-06, 4.758262e-06, 4.940405e-06, 4.797696e-06, 5.05852e-06, 
    4.912084e-06, 4.828431e-06, 4.509516e-06, 4.440314e-06, 4.376518e-06, 
    4.251397e-06, 4.090122e-06, 3.817609e-06, 3.586698e-06, 3.381401e-06, 
    3.396251e-06, 3.391021e-06, 3.345877e-06, 3.45824e-06, 3.327595e-06, 
    3.305917e-06, 3.362765e-06, 3.039393e-06, 3.130109e-06, 3.037297e-06, 
    3.096183e-06, 4.74131e-06, 4.653862e-06, 4.701058e-06, 4.612438e-06, 
    4.674834e-06, 4.399468e-06, 4.317975e-06, 3.941412e-06, 4.093231e-06, 
    3.85261e-06, 4.068521e-06, 4.029944e-06, 3.844932e-06, 4.056727e-06, 
    3.599302e-06, 3.907093e-06, 3.344128e-06, 3.642132e-06, 3.325847e-06, 
    3.382277e-06, 3.289077e-06, 3.206687e-06, 3.104479e-06, 2.920413e-06, 
    2.962501e-06, 2.812008e-06, 4.524403e-06, 4.412746e-06, 4.422506e-06, 
    4.30654e-06, 4.221466e-06, 4.036587e-06, 3.750976e-06, 3.857389e-06, 
    3.662944e-06, 3.624431e-06, 3.920166e-06, 3.737482e-06, 4.33851e-06, 
    4.239582e-06, 4.298362e-06, 4.515583e-06, 3.832805e-06, 4.179353e-06, 
    3.551044e-06, 3.730276e-06, 3.218375e-06, 3.46869e-06, 2.985814e-06, 
    2.790849e-06, 2.614006e-06, 2.416257e-06, 4.352159e-06, 4.427589e-06, 
    4.292809e-06, 4.106179e-06, 3.938209e-06, 3.719241e-06, 3.697111e-06, 
    3.656776e-06, 3.553148e-06, 3.467054e-06, 3.644094e-06, 3.445618e-06, 
    4.216823e-06, 3.80349e-06, 4.456252e-06, 4.256537e-06, 4.116918e-06, 
    4.17941e-06, 3.869619e-06, 3.798588e-06, 3.515648e-06, 3.660723e-06, 
    2.838318e-06, 3.189458e-06, 2.272227e-06, 2.509996e-06, 4.454054e-06, 
    4.352402e-06, 4.002604e-06, 4.169048e-06, 3.70479e-06, 3.594586e-06, 
    3.506041e-06, 3.394356e-06, 3.382375e-06, 3.317099e-06, 3.424381e-06, 
    3.321294e-06, 3.718781e-06, 3.538667e-06, 4.041681e-06, 3.916784e-06, 
    3.974042e-06, 4.037241e-06, 3.843445e-06, 3.641285e-06, 3.636964e-06, 
    3.573165e-06, 3.396185e-06, 3.702964e-06, 2.794686e-06, 3.341057e-06, 
    4.24247e-06, 4.048253e-06, 4.021109e-06, 4.094715e-06, 3.605572e-06, 
    3.779896e-06, 3.318675e-06, 3.440657e-06, 3.241875e-06, 3.339957e-06, 
    3.354507e-06, 3.482748e-06, 3.563708e-06, 3.771837e-06, 3.94476e-06, 
    4.084001e-06, 4.051457e-06, 3.899076e-06, 3.629057e-06, 3.381313e-06, 
    3.43491e-06, 3.256782e-06, 3.737529e-06, 3.532348e-06, 3.611075e-06, 
    3.407423e-06, 3.860245e-06, 3.473222e-06, 3.961892e-06, 3.917982e-06, 
    3.78339e-06, 3.518649e-06, 3.461142e-06, 3.400306e-06, 3.437776e-06, 
    3.622298e-06, 3.65291e-06, 3.786626e-06, 3.823922e-06, 3.927521e-06, 
    4.014138e-06, 3.934984e-06, 3.852535e-06, 3.622198e-06, 3.419928e-06, 
    3.205529e-06, 3.154071e-06, 2.914481e-06, 3.10884e-06, 2.791797e-06, 
    3.060286e-06, 2.604195e-06, 3.45127e-06, 3.068285e-06, 3.777294e-06, 
    3.697721e-06, 3.555688e-06, 3.239333e-06, 3.408367e-06, 3.21107e-06, 
    3.654107e-06, 3.893887e-06, 3.956857e-06, 4.075494e-06, 3.954161e-06, 
    3.963974e-06, 3.849097e-06, 3.885864e-06, 3.614653e-06, 3.759322e-06, 
    3.354887e-06, 3.212594e-06, 2.827593e-06, 2.604924e-06, 2.389415e-06, 
    2.29806e-06, 2.270721e-06, 2.25936e-06,
  7.830568e-06, 7.669986e-06, 7.700953e-06, 7.573319e-06, 7.643845e-06, 
    7.560671e-06, 7.797758e-06, 7.663677e-06, 7.749013e-06, 7.815985e-06, 
    7.332453e-06, 7.567678e-06, 6.816638e-06, 6.927026e-06, 6.657101e-06, 
    6.833568e-06, 6.622889e-06, 6.662035e-06, 6.546119e-06, 6.57874e-06, 
    6.436879e-06, 6.531226e-06, 6.367298e-06, 6.459001e-06, 6.444343e-06, 
    6.534414e-06, 7.519624e-06, 7.361233e-06, 7.529136e-06, 7.506265e-06, 
    7.516519e-06, 7.642381e-06, 7.706652e-06, 7.842972e-06, 7.818058e-06, 
    7.718014e-06, 7.496008e-06, 7.570584e-06, 7.384305e-06, 7.388449e-06, 
    6.885909e-06, 6.955417e-06, 6.703731e-06, 6.773163e-06, 6.577369e-06, 
    6.625196e-06, 6.579594e-06, 6.593328e-06, 6.579416e-06, 6.649952e-06, 
    6.619476e-06, 6.682475e-06, 6.942292e-06, 6.863643e-06, 7.467282e-06, 
    7.660557e-06, 7.79183e-06, 7.886254e-06, 7.872844e-06, 7.847335e-06, 
    7.717433e-06, 7.597225e-06, 7.506968e-06, 7.447285e-06, 7.389046e-06, 
    6.908068e-06, 6.839027e-06, 6.689902e-06, 6.716239e-06, 6.671777e-06, 
    6.630008e-06, 6.561471e-06, 6.572613e-06, 6.542915e-06, 6.672941e-06, 
    6.585724e-06, 6.731355e-06, 6.690693e-06, 7.3733e-06, 7.550383e-06, 
    7.627128e-06, 7.69499e-06, 7.862547e-06, 7.746471e-06, 7.792039e-06, 
    7.684053e-06, 7.616214e-06, 7.649689e-06, 7.445661e-06, 7.524238e-06, 
    6.834981e-06, 6.966539e-06, 6.634843e-06, 6.710812e-06, 6.616971e-06, 
    6.664423e-06, 6.583679e-06, 6.656227e-06, 6.531965e-06, 6.505803e-06, 
    6.523646e-06, 6.455951e-06, 6.660313e-06, 6.579594e-06, 7.650629e-06, 
    7.645158e-06, 7.619725e-06, 7.73217e-06, 7.739102e-06, 7.843655e-06, 
    7.750561e-06, 7.711235e-06, 7.612301e-06, 7.554414e-06, 7.499842e-06, 
    7.381502e-06, 6.935866e-06, 6.799889e-06, 6.70582e-06, 6.64454e-06, 
    6.681944e-06, 6.648893e-06, 6.685868e-06, 6.703382e-06, 6.515567e-06, 
    6.619193e-06, 6.465546e-06, 6.473759e-06, 6.542214e-06, 6.472832e-06, 
    7.641319e-06, 7.672839e-06, 7.783284e-06, 7.69672e-06, 7.855118e-06, 
    7.76608e-06, 7.71531e-06, 7.522583e-06, 7.480959e-06, 7.442603e-06, 
    7.367567e-06, 6.951825e-06, 6.825979e-06, 6.720481e-06, 6.627599e-06, 
    6.63429e-06, 6.631933e-06, 6.611609e-06, 6.662262e-06, 6.603394e-06, 
    6.593653e-06, 6.619206e-06, 6.474861e-06, 6.515115e-06, 6.473934e-06, 
    6.50004e-06, 7.662579e-06, 7.609693e-06, 7.638223e-06, 7.584667e-06, 
    7.622355e-06, 7.456364e-06, 7.407429e-06, 6.882956e-06, 6.953264e-06, 
    6.842058e-06, 6.9418e-06, 6.923909e-06, 6.838492e-06, 6.936335e-06, 
    6.726198e-06, 6.867119e-06, 6.610822e-06, 6.745678e-06, 6.602609e-06, 
    6.627994e-06, 6.586112e-06, 6.549238e-06, 6.503721e-06, 6.422356e-06, 
    6.44089e-06, 6.374853e-06, 7.531581e-06, 7.46436e-06, 7.470253e-06, 
    7.400614e-06, 7.34964e-06, 6.926998e-06, 6.795435e-06, 6.844275e-06, 
    6.755215e-06, 6.737658e-06, 6.873188e-06, 6.789251e-06, 7.419776e-06, 
    7.360452e-06, 7.395702e-06, 7.526251e-06, 6.83295e-06, 7.32442e-06, 
    6.704292e-06, 6.785965e-06, 6.554458e-06, 6.666968e-06, 6.451172e-06, 
    6.365588e-06, 6.288929e-06, 6.204322e-06, 7.427979e-06, 7.47331e-06, 
    7.392387e-06, 6.959262e-06, 6.881501e-06, 6.780916e-06, 6.77081e-06, 
    6.752397e-06, 6.705256e-06, 6.66625e-06, 6.746599e-06, 6.656563e-06, 
    7.346777e-06, 6.819498e-06, 7.490533e-06, 7.3706e-06, 6.964261e-06, 
    7.324483e-06, 6.849906e-06, 6.817266e-06, 6.688231e-06, 6.754202e-06, 
    6.386322e-06, 6.541527e-06, 6.143648e-06, 6.244255e-06, 7.489226e-06, 
    7.428136e-06, 6.911247e-06, 7.318293e-06, 6.774318e-06, 6.724075e-06, 
    6.683896e-06, 6.633424e-06, 6.628035e-06, 6.598676e-06, 6.646975e-06, 
    6.600565e-06, 6.780705e-06, 6.698679e-06, 6.929363e-06, 6.871619e-06, 
    6.89806e-06, 6.927305e-06, 6.837867e-06, 6.745315e-06, 6.74337e-06, 
    6.714331e-06, 6.63417e-06, 6.773484e-06, 6.367219e-06, 6.60937e-06, 
    7.362226e-06, 6.932373e-06, 6.919825e-06, 6.953965e-06, 6.729072e-06, 
    6.808687e-06, 6.599387e-06, 6.654322e-06, 6.564971e-06, 6.60895e-06, 
    6.615491e-06, 6.673349e-06, 6.710044e-06, 6.804989e-06, 6.884523e-06, 
    6.948993e-06, 6.933894e-06, 6.863454e-06, 6.739748e-06, 6.627547e-06, 
    6.65171e-06, 6.571642e-06, 6.789287e-06, 6.695803e-06, 6.731565e-06, 
    6.63932e-06, 6.845583e-06, 6.668963e-06, 6.892447e-06, 6.87218e-06, 
    6.810289e-06, 6.689576e-06, 6.663577e-06, 6.636105e-06, 6.653021e-06, 
    6.736675e-06, 6.75063e-06, 6.811779e-06, 6.828885e-06, 6.876582e-06, 
    6.916606e-06, 6.880019e-06, 6.84203e-06, 6.73664e-06, 6.644952e-06, 
    6.548717e-06, 6.52578e-06, 6.419713e-06, 6.50562e-06, 6.365955e-06, 
    6.484023e-06, 6.284649e-06, 6.659071e-06, 6.487613e-06, 6.807502e-06, 
    6.77109e-06, 6.706382e-06, 6.563803e-06, 6.639747e-06, 6.551177e-06, 
    6.751179e-06, 6.861049e-06, 6.890119e-06, 6.945038e-06, 6.888874e-06, 
    6.893407e-06, 6.840467e-06, 6.857385e-06, 6.733205e-06, 6.799267e-06, 
    6.615655e-06, 6.551863e-06, 6.381656e-06, 6.284994e-06, 6.192974e-06, 
    6.154477e-06, 6.143026e-06, 6.138275e-06,
  9.692789e-06, 9.704461e-06, 9.702402e-06, 9.710255e-06, 9.706125e-06, 
    9.710939e-06, 9.69537e-06, 9.704868e-06, 9.699022e-06, 9.693948e-06, 
    9.720047e-06, 9.710562e-06, 1.004597e-05, 1.008924e-05, 9.97865e-06, 
    1.005276e-05, 9.963364e-06, 9.980834e-06, 9.927802e-06, 9.943139e-06, 
    9.873744e-06, 9.920685e-06, 9.83684e-06, 9.885055e-06, 9.877584e-06, 
    9.922214e-06, 9.713038e-06, 9.719257e-06, 9.712568e-06, 9.713679e-06, 
    9.713189e-06, 9.706215e-06, 9.702012e-06, 9.691789e-06, 9.693785e-06, 
    9.701227e-06, 9.714157e-06, 9.710405e-06, 9.718552e-06, 9.718417e-06, 
    1.007341e-05, 1.009999e-05, 9.99898e-06, 1.002823e-05, 9.942501e-06, 
    9.964411e-06, 9.943535e-06, 9.949888e-06, 9.943452e-06, 9.975489e-06, 
    9.961825e-06, 9.989787e-06, 1.009504e-05, 1.00647e-05, 9.715432e-06, 
    9.705066e-06, 9.695825e-06, 9.688193e-06, 9.689325e-06, 9.691434e-06, 
    9.701268e-06, 9.708915e-06, 9.713647e-06, 9.716263e-06, 9.718397e-06, 
    1.008197e-05, 1.005494e-05, 9.993009e-06, 1.000434e-05, 9.985112e-06, 
    9.966578e-06, 9.935061e-06, 9.940283e-06, 9.926275e-06, 9.985625e-06, 
    9.946375e-06, 1.001076e-05, 9.993356e-06, 9.718893e-06, 9.711483e-06, 
    9.707149e-06, 9.702806e-06, 9.690182e-06, 9.699205e-06, 9.695809e-06, 
    9.703539e-06, 9.707805e-06, 9.705759e-06, 9.716327e-06, 9.712812e-06, 
    1.005333e-05, 1.010416e-05, 9.968749e-06, 1.000202e-05, 9.960691e-06, 
    9.981888e-06, 9.945429e-06, 9.978272e-06, 9.921038e-06, 9.908355e-06, 
    9.91703e-06, 9.883512e-06, 9.980075e-06, 9.943533e-06, 9.7057e-06, 
    9.706043e-06, 9.707597e-06, 9.700231e-06, 9.699736e-06, 9.691733e-06, 
    9.69891e-06, 9.701698e-06, 9.708038e-06, 9.711272e-06, 9.713981e-06, 
    9.718641e-06, 1.00926e-05, 1.003918e-05, 9.999878e-06, 9.973083e-06, 
    9.989558e-06, 9.97502e-06, 9.991263e-06, 9.998832e-06, 9.913116e-06, 
    9.961695e-06, 9.888367e-06, 9.892495e-06, 9.92594e-06, 9.89203e-06, 
    9.706282e-06, 9.704277e-06, 9.696477e-06, 9.70269e-06, 9.690796e-06, 
    9.697767e-06, 9.701415e-06, 9.712892e-06, 9.714839e-06, 9.716449e-06, 
    9.719075e-06, 1.009864e-05, 1.004973e-05, 1.000614e-05, 9.965494e-06, 
    9.968502e-06, 9.967443e-06, 9.958256e-06, 9.980935e-06, 9.954508e-06, 
    9.950036e-06, 9.961704e-06, 9.893047e-06, 9.912899e-06, 9.892582e-06, 
    9.905533e-06, 9.704941e-06, 9.708191e-06, 9.706473e-06, 9.709626e-06, 
    9.707439e-06, 9.71589e-06, 9.717766e-06, 1.007226e-05, 1.009918e-05, 
    1.005615e-05, 1.009486e-05, 1.008805e-05, 1.005473e-05, 1.009279e-05, 
    1.000857e-05, 1.006606e-05, 9.957897e-06, 1.001678e-05, 9.954148e-06, 
    9.965673e-06, 9.946558e-06, 9.929282e-06, 9.90734e-06, 9.866219e-06, 
    9.875815e-06, 9.840955e-06, 9.712447e-06, 9.715556e-06, 9.715306e-06, 
    9.718006e-06, 9.719594e-06, 1.008923e-05, 1.003737e-05, 1.005704e-05, 
    1.002078e-05, 1.001342e-05, 1.006845e-05, 1.003484e-05, 9.717322e-06, 
    9.719284e-06, 9.718174e-06, 9.712711e-06, 1.005252e-05, 9.720252e-06, 
    9.999221e-06, 1.00335e-05, 9.931753e-06, 9.983001e-06, 9.881078e-06, 
    9.8359e-06, 9.792494e-06, 9.740605e-06, 9.717017e-06, 9.715174e-06, 
    9.718286e-06, 1.010143e-05, 1.007169e-05, 1.003142e-05, 1.002726e-05, 
    1.00196e-05, 9.999637e-06, 9.98269e-06, 1.001717e-05, 9.97842e-06, 
    9.719669e-06, 1.004712e-05, 9.714408e-06, 9.71898e-06, 1.010331e-05, 
    9.720252e-06, 1.005928e-05, 1.004623e-05, 9.992285e-06, 1.002036e-05, 
    9.847138e-06, 9.925608e-06, 9.700265e-06, 9.765668e-06, 9.714468e-06, 
    9.717011e-06, 1.00832e-05, 9.7204e-06, 1.002871e-05, 1.000767e-05, 
    9.990407e-06, 9.96811e-06, 9.965691e-06, 9.952345e-06, 9.974167e-06, 
    9.953214e-06, 1.003134e-05, 9.996807e-06, 1.009014e-05, 1.006783e-05, 
    1.007813e-05, 1.008935e-05, 1.005449e-05, 1.001663e-05, 1.001582e-05, 
    1.000352e-05, 9.968427e-06, 1.002836e-05, 9.836778e-06, 9.957218e-06, 
    9.719234e-06, 1.009127e-05, 1.008649e-05, 1.009945e-05, 1.000979e-05, 
    1.004276e-05, 9.952672e-06, 9.977428e-06, 9.936706e-06, 9.957044e-06, 
    9.960019e-06, 9.985804e-06, 1.000169e-05, 1.004126e-05, 1.007287e-05, 
    1.009757e-05, 1.009186e-05, 1.006462e-05, 1.001429e-05, 9.965469e-06, 
    9.976266e-06, 9.93983e-06, 1.003486e-05, 9.995563e-06, 1.001084e-05, 
    9.970753e-06, 1.005756e-05, 9.983865e-06, 1.007595e-05, 1.006805e-05, 
    1.004341e-05, 9.992866e-06, 9.981515e-06, 9.969312e-06, 9.976852e-06, 
    1.0013e-05, 1.001886e-05, 1.004401e-05, 1.00509e-05, 1.006977e-05, 
    1.008526e-05, 1.007112e-05, 1.005614e-05, 1.001299e-05, 9.973264e-06, 
    9.929034e-06, 9.918062e-06, 9.864829e-06, 9.908259e-06, 9.836087e-06, 
    9.897593e-06, 9.789959e-06, 9.979518e-06, 9.899387e-06, 1.004228e-05, 
    1.002737e-05, 1.000011e-05, 9.93615e-06, 9.970943e-06, 9.930196e-06, 
    1.001909e-05, 1.006367e-05, 1.007505e-05, 1.009608e-05, 1.007456e-05, 
    1.007632e-05, 1.005552e-05, 1.006223e-05, 1.001154e-05, 1.003893e-05, 
    9.960093e-06, 9.930523e-06, 9.844633e-06, 9.790174e-06, 9.733287e-06, 
    9.707688e-06, 9.699838e-06, 9.696548e-06,
  4.369422e-06, 4.283264e-06, 4.300002e-06, 4.230608e-06, 4.269091e-06, 
    4.223671e-06, 4.351944e-06, 4.279844e-06, 4.32586e-06, 4.361664e-06, 
    4.096308e-06, 4.227516e-06, 3.960917e-06, 4.044181e-06, 3.835542e-06, 
    3.973852e-06, 3.807754e-06, 3.83953e-06, 3.744054e-06, 3.771363e-06, 
    3.649707e-06, 3.731462e-06, 3.586964e-06, 3.669205e-06, 3.656311e-06, 
    3.734164e-06, 4.20108e-06, 4.112612e-06, 4.206327e-06, 4.193696e-06, 
    4.199364e-06, 4.268292e-06, 4.303069e-06, 4.37602e-06, 4.362768e-06, 
    4.309195e-06, 4.188018e-06, 4.229114e-06, 4.125651e-06, 4.127984e-06, 
    4.013469e-06, 4.065196e-06, 3.872883e-06, 3.927399e-06, 3.770223e-06, 
    3.809646e-06, 3.772071e-06, 3.783459e-06, 3.771923e-06, 3.829772e-06, 
    3.804967e-06, 3.855942e-06, 4.055499e-06, 3.996691e-06, 4.172078e-06, 
    4.278147e-06, 4.348778e-06, 4.398961e-06, 4.391863e-06, 4.378334e-06, 
    4.308882e-06, 4.243695e-06, 4.194089e-06, 4.160945e-06, 4.12832e-06, 
    4.030047e-06, 3.978014e-06, 3.86187e-06, 3.882798e-06, 3.847362e-06, 
    3.813572e-06, 3.756949e-06, 3.76626e-06, 3.741348e-06, 3.848302e-06, 
    3.777158e-06, 3.894724e-06, 3.862508e-06, 4.119425e-06, 4.218024e-06, 
    4.25999e-06, 4.296783e-06, 4.386406e-06, 4.324493e-06, 4.348889e-06, 
    4.290879e-06, 4.254056e-06, 4.272265e-06, 4.160039e-06, 4.203627e-06, 
    3.974933e-06, 4.073381e-06, 3.817511e-06, 3.878502e-06, 3.802918e-06, 
    3.841456e-06, 3.775462e-06, 3.834848e-06, 3.732087e-06, 3.709775e-06, 
    3.725019e-06, 3.666536e-06, 3.838144e-06, 3.772069e-06, 4.272774e-06, 
    4.269803e-06, 4.255971e-06, 4.316811e-06, 4.320537e-06, 4.376382e-06, 
    4.32669e-06, 4.305545e-06, 4.251925e-06, 4.220239e-06, 4.190145e-06, 
    4.12407e-06, 4.050737e-06, 3.948056e-06, 3.874542e-06, 3.825391e-06, 
    3.855519e-06, 3.828918e-06, 3.858656e-06, 3.872609e-06, 3.71813e-06, 
    3.804734e-06, 3.674937e-06, 3.682098e-06, 3.740755e-06, 3.681291e-06, 
    4.267718e-06, 4.284814e-06, 4.344213e-06, 4.29772e-06, 4.382468e-06, 
    4.335006e-06, 4.307738e-06, 4.202709e-06, 4.17968e-06, 4.15833e-06, 
    4.116212e-06, 4.062546e-06, 3.96807e-06, 3.886147e-06, 3.81161e-06, 
    3.817063e-06, 3.815142e-06, 3.798519e-06, 3.839715e-06, 3.791764e-06, 
    3.783724e-06, 3.804748e-06, 3.683057e-06, 3.717749e-06, 3.68225e-06, 
    3.704831e-06, 4.279257e-06, 4.250501e-06, 4.266036e-06, 4.236826e-06, 
    4.257401e-06, 4.165998e-06, 4.13864e-06, 4.011243e-06, 4.063606e-06, 
    3.980325e-06, 4.055138e-06, 4.041865e-06, 3.9776e-06, 4.051092e-06, 
    3.890651e-06, 3.999308e-06, 3.797874e-06, 3.90595e-06, 3.791118e-06, 
    3.811931e-06, 3.777485e-06, 3.746678e-06, 3.707993e-06, 3.636805e-06, 
    3.653267e-06, 3.593895e-06, 4.207676e-06, 4.170452e-06, 4.173733e-06, 
    4.134822e-06, 4.106073e-06, 4.044164e-06, 3.944628e-06, 3.982017e-06, 
    3.913425e-06, 3.899675e-06, 4.003901e-06, 3.939853e-06, 4.145567e-06, 
    4.112184e-06, 4.13206e-06, 4.204735e-06, 3.973388e-06, 4.091758e-06, 
    3.873328e-06, 3.937317e-06, 3.751067e-06, 3.843496e-06, 3.662334e-06, 
    3.585385e-06, 3.5133e-06, 3.429433e-06, 4.15016e-06, 4.175433e-06, 
    4.1302e-06, 4.068022e-06, 4.010157e-06, 3.933408e-06, 3.925571e-06, 
    3.911221e-06, 3.874097e-06, 3.842926e-06, 3.90668e-06, 3.835119e-06, 
    4.104436e-06, 3.963113e-06, 4.184987e-06, 4.117915e-06, 4.071706e-06, 
    4.091798e-06, 3.986294e-06, 3.96141e-06, 3.860538e-06, 3.912634e-06, 
    3.604341e-06, 3.740168e-06, 3.365906e-06, 3.469636e-06, 4.184266e-06, 
    4.150249e-06, 4.032433e-06, 4.088277e-06, 3.928295e-06, 3.888985e-06, 
    3.857081e-06, 3.816353e-06, 3.811964e-06, 3.787874e-06, 3.827364e-06, 
    3.789435e-06, 3.933244e-06, 3.86887e-06, 4.045921e-06, 4.002715e-06, 
    4.022585e-06, 4.044393e-06, 3.977143e-06, 3.905674e-06, 3.904158e-06, 
    3.881285e-06, 3.816932e-06, 3.927648e-06, 3.586865e-06, 3.796654e-06, 
    4.113196e-06, 4.048143e-06, 4.038828e-06, 4.064127e-06, 3.892923e-06, 
    3.954827e-06, 3.788462e-06, 3.833309e-06, 3.75988e-06, 3.796336e-06, 
    3.801704e-06, 3.848631e-06, 3.877893e-06, 3.951983e-06, 4.012428e-06, 
    4.060458e-06, 4.049283e-06, 3.996548e-06, 3.901311e-06, 3.811563e-06, 
    3.831191e-06, 3.765451e-06, 3.939886e-06, 3.866577e-06, 3.894882e-06, 
    3.821152e-06, 3.983009e-06, 3.845081e-06, 4.01838e-06, 4.003141e-06, 
    3.956057e-06, 3.861606e-06, 3.840774e-06, 3.818535e-06, 3.832257e-06, 
    3.898899e-06, 3.90984e-06, 3.957203e-06, 3.97029e-06, 4.006459e-06, 
    4.036435e-06, 4.009044e-06, 3.980305e-06, 3.898875e-06, 3.82572e-06, 
    3.746238e-06, 3.726837e-06, 3.63443e-06, 3.709607e-06, 3.585702e-06, 
    3.690973e-06, 3.50915e-06, 3.837126e-06, 3.694096e-06, 3.95392e-06, 
    3.92579e-06, 3.874981e-06, 3.758891e-06, 3.821498e-06, 3.748302e-06, 
    3.910269e-06, 3.994726e-06, 4.016634e-06, 4.057534e-06, 4.015699e-06, 
    4.0191e-06, 3.979122e-06, 3.991963e-06, 3.896176e-06, 3.947584e-06, 
    3.801837e-06, 3.748882e-06, 3.600104e-06, 3.509498e-06, 3.417799e-06, 
    3.377488e-06, 3.365241e-06, 3.360124e-06,
  4.506543e-07, 4.337497e-07, 4.370064e-07, 4.235899e-07, 4.310022e-07, 
    4.222611e-07, 4.471969e-07, 4.330859e-07, 4.420635e-07, 4.491178e-07, 
    3.982628e-07, 4.229974e-07, 3.73526e-07, 3.886024e-07, 3.514235e-07, 
    3.758472e-07, 3.466216e-07, 3.521154e-07, 3.357462e-07, 3.403862e-07, 
    3.199751e-07, 3.336181e-07, 3.097085e-07, 3.232015e-07, 3.210661e-07, 
    3.340741e-07, 4.179492e-07, 4.012929e-07, 4.189485e-07, 4.16545e-07, 
    4.176228e-07, 4.308477e-07, 4.376045e-07, 4.519633e-07, 4.493364e-07, 
    4.388008e-07, 4.15467e-07, 4.233036e-07, 4.037248e-07, 4.041609e-07, 
    3.830044e-07, 3.924579e-07, 3.579314e-07, 3.675466e-07, 3.401917e-07, 
    3.469475e-07, 3.405069e-07, 3.424522e-07, 3.404816e-07, 3.504234e-07, 
    3.46142e-07, 3.54971e-07, 3.906764e-07, 3.799643e-07, 4.124487e-07, 
    4.327566e-07, 4.465721e-07, 4.565306e-07, 4.551148e-07, 4.524229e-07, 
    4.387396e-07, 4.261028e-07, 4.166198e-07, 4.103476e-07, 4.042236e-07, 
    3.860208e-07, 3.765957e-07, 3.560055e-07, 3.5967e-07, 3.534767e-07, 
    3.476242e-07, 3.379329e-07, 3.395165e-07, 3.352883e-07, 3.536402e-07, 
    3.413751e-07, 3.617674e-07, 3.561167e-07, 4.025626e-07, 4.211811e-07, 
    4.29243e-07, 4.363791e-07, 4.54028e-07, 4.417954e-07, 4.465939e-07, 
    4.352297e-07, 4.280981e-07, 4.316167e-07, 4.101769e-07, 4.184342e-07, 
    3.760416e-07, 3.939652e-07, 3.483037e-07, 3.589161e-07, 3.457896e-07, 
    3.5245e-07, 3.410856e-07, 3.513031e-07, 3.337236e-07, 3.299697e-07, 
    3.32532e-07, 3.227589e-07, 3.518748e-07, 3.405065e-07, 4.317153e-07, 
    4.311402e-07, 4.284673e-07, 4.402902e-07, 4.4102e-07, 4.520352e-07, 
    4.422265e-07, 4.380878e-07, 4.276873e-07, 4.216045e-07, 4.158707e-07, 
    4.034295e-07, 3.898029e-07, 3.712256e-07, 3.582221e-07, 3.496652e-07, 
    3.548973e-07, 3.502756e-07, 3.554444e-07, 3.578835e-07, 3.313728e-07, 
    3.461019e-07, 3.241533e-07, 3.253444e-07, 3.35188e-07, 3.252101e-07, 
    4.307367e-07, 4.340506e-07, 4.45672e-07, 4.365617e-07, 4.532445e-07, 
    4.438599e-07, 4.38516e-07, 4.182593e-07, 4.138867e-07, 4.09855e-07, 
    4.019634e-07, 3.919706e-07, 3.748085e-07, 3.602583e-07, 3.472858e-07, 
    3.482264e-07, 3.47895e-07, 3.450337e-07, 3.521476e-07, 3.438745e-07, 
    3.424975e-07, 3.461043e-07, 3.255041e-07, 3.313087e-07, 3.253698e-07, 
    3.29141e-07, 4.329719e-07, 4.274129e-07, 4.304114e-07, 4.24783e-07, 
    4.287432e-07, 4.113005e-07, 4.061554e-07, 3.826003e-07, 3.921655e-07, 
    3.770116e-07, 3.9061e-07, 3.881787e-07, 3.765211e-07, 3.89868e-07, 
    3.610503e-07, 3.804377e-07, 3.449228e-07, 3.637474e-07, 3.437636e-07, 
    3.473413e-07, 3.414309e-07, 3.361906e-07, 3.296709e-07, 3.178495e-07, 
    3.205629e-07, 3.108338e-07, 4.192057e-07, 4.121415e-07, 4.127616e-07, 
    4.054402e-07, 4.000761e-07, 3.885992e-07, 3.706137e-07, 3.773162e-07, 
    3.650691e-07, 3.6264e-07, 3.812692e-07, 3.697623e-07, 4.074548e-07, 
    4.012131e-07, 4.049232e-07, 4.186452e-07, 3.757637e-07, 3.974193e-07, 
    3.580094e-07, 3.693105e-07, 3.369345e-07, 3.528043e-07, 3.220626e-07, 
    3.094524e-07, 2.978794e-07, 2.84706e-07, 4.083177e-07, 4.13083e-07, 
    4.045751e-07, 3.92978e-07, 3.824032e-07, 3.686148e-07, 3.672221e-07, 
    3.646792e-07, 3.58144e-07, 3.527053e-07, 3.638764e-07, 3.513501e-07, 
    3.997717e-07, 3.739194e-07, 4.148922e-07, 4.022809e-07, 3.936564e-07, 
    3.974268e-07, 3.780872e-07, 3.736142e-07, 3.557728e-07, 3.649292e-07, 
    3.125342e-07, 3.350888e-07, 2.749348e-07, 2.909818e-07, 4.147555e-07, 
    4.083346e-07, 3.864558e-07, 3.967748e-07, 3.67706e-07, 3.607573e-07, 
    3.551696e-07, 3.481038e-07, 3.47347e-07, 3.432078e-07, 3.500066e-07, 
    3.434752e-07, 3.685858e-07, 3.572289e-07, 3.889209e-07, 3.810544e-07, 
    3.846615e-07, 3.886411e-07, 3.764389e-07, 3.636986e-07, 3.63431e-07, 
    3.594044e-07, 3.482038e-07, 3.67591e-07, 3.096925e-07, 3.447133e-07, 
    4.014015e-07, 3.893278e-07, 3.876235e-07, 3.922613e-07, 3.614502e-07, 
    3.724357e-07, 3.433086e-07, 3.510362e-07, 3.38431e-07, 3.446587e-07, 
    3.455809e-07, 3.536974e-07, 3.588093e-07, 3.719272e-07, 3.828152e-07, 
    3.915868e-07, 3.895365e-07, 3.799387e-07, 3.629284e-07, 3.472777e-07, 
    3.506693e-07, 3.393789e-07, 3.697682e-07, 3.568278e-07, 3.617951e-07, 
    3.489325e-07, 3.77495e-07, 3.530799e-07, 3.838965e-07, 3.811315e-07, 
    3.726558e-07, 3.559593e-07, 3.523316e-07, 3.484806e-07, 3.508541e-07, 
    3.625031e-07, 3.644348e-07, 3.728608e-07, 3.752073e-07, 3.817326e-07, 
    3.871863e-07, 3.822012e-07, 3.77008e-07, 3.624988e-07, 3.497222e-07, 
    3.361161e-07, 3.328383e-07, 3.174591e-07, 3.299416e-07, 3.095037e-07, 
    3.268238e-07, 2.972201e-07, 3.516983e-07, 3.273454e-07, 3.722734e-07, 
    3.672609e-07, 3.582989e-07, 3.38263e-07, 3.489923e-07, 3.364659e-07, 
    3.645107e-07, 3.796092e-07, 3.835791e-07, 3.910498e-07, 3.834093e-07, 
    3.840274e-07, 3.76795e-07, 3.791101e-07, 3.620231e-07, 3.711414e-07, 
    3.456036e-07, 3.365641e-07, 3.11844e-07, 2.972754e-07, 2.829032e-07, 
    2.767029e-07, 2.748335e-07, 2.740544e-07,
  1.268738e-08, 1.195778e-08, 1.209717e-08, 1.152654e-08, 1.184061e-08, 
    1.147054e-08, 1.253694e-08, 1.192943e-08, 1.231473e-08, 1.262045e-08, 
    1.047571e-08, 1.150156e-08, 9.483518e-09, 1.008415e-08, 8.626416e-09, 
    9.575158e-09, 8.443965e-09, 8.652821e-09, 8.035793e-09, 8.209077e-09, 
    7.45652e-09, 7.956751e-09, 7.092817e-09, 7.573793e-09, 7.496102e-09, 
    7.973664e-09, 1.128949e-08, 1.059958e-08, 1.133136e-08, 1.123075e-08, 
    1.127583e-08, 1.183404e-08, 1.212283e-08, 1.27445e-08, 1.262997e-08, 
    1.217421e-08, 1.118573e-08, 1.151446e-08, 1.069937e-08, 1.07173e-08, 
    9.859639e-09, 1.02398e-08, 8.875847e-09, 9.24887e-09, 8.20179e-09, 
    8.456305e-09, 8.213606e-09, 8.286646e-09, 8.212657e-09, 8.588308e-09, 
    8.425816e-09, 8.762076e-09, 1.016778e-08, 9.738453e-09, 1.106e-08, 
    1.191538e-08, 1.250982e-08, 1.29445e-08, 1.288239e-08, 1.276458e-08, 
    1.217158e-08, 1.163269e-08, 1.123388e-08, 1.097276e-08, 1.071988e-08, 
    9.980399e-09, 9.604775e-09, 8.801774e-09, 8.942899e-09, 8.704844e-09, 
    8.481948e-09, 8.117299e-09, 8.176501e-09, 8.018763e-09, 8.711101e-09, 
    8.246177e-09, 9.024023e-09, 8.806047e-09, 1.065165e-08, 1.14251e-08, 
    1.176581e-08, 1.207027e-08, 1.283478e-08, 1.230316e-08, 1.251077e-08, 
    1.202105e-08, 1.171721e-08, 1.186679e-08, 1.096568e-08, 1.130981e-08, 
    9.582846e-09, 1.030088e-08, 8.507723e-09, 8.9138e-09, 8.412488e-09, 
    8.665597e-09, 8.235308e-09, 8.621825e-09, 7.960661e-09, 7.82187e-09, 
    7.916512e-09, 7.557666e-09, 8.643636e-09, 8.213587e-09, 1.187099e-08, 
    1.184649e-08, 1.173288e-08, 1.223829e-08, 1.226973e-08, 1.274764e-08, 
    1.232176e-08, 1.214358e-08, 1.169979e-08, 1.144291e-08, 1.120258e-08, 
    1.068724e-08, 1.013253e-08, 9.393004e-09, 8.887046e-09, 8.559454e-09, 
    8.759252e-09, 8.582678e-09, 8.780236e-09, 8.874e-09, 7.873647e-09, 
    8.4243e-09, 7.608509e-09, 7.652036e-09, 8.015033e-09, 7.647122e-09, 
    1.182931e-08, 1.197063e-08, 1.247079e-08, 1.20781e-08, 1.280049e-08, 
    1.239233e-08, 1.216197e-08, 1.130248e-08, 1.111984e-08, 1.095235e-08, 
    1.062707e-08, 1.022009e-08, 9.534115e-09, 8.965629e-09, 8.469121e-09, 
    8.504789e-09, 8.492218e-09, 8.383929e-09, 8.654046e-09, 8.340196e-09, 
    8.28835e-09, 8.42439e-09, 7.657879e-09, 7.871281e-09, 7.652963e-09, 
    7.791346e-09, 1.192457e-08, 1.168816e-08, 1.181547e-08, 1.157689e-08, 
    1.174458e-08, 1.10123e-08, 1.079943e-08, 9.843503e-09, 1.022797e-08, 
    9.621244e-09, 1.01651e-08, 1.00671e-08, 9.601822e-09, 1.013516e-08, 
    8.99626e-09, 9.757287e-09, 8.379741e-09, 9.100843e-09, 8.33602e-09, 
    8.471223e-09, 8.248271e-09, 8.052333e-09, 7.810858e-09, 7.379607e-09, 
    7.477837e-09, 7.127738e-09, 1.134215e-08, 1.104723e-08, 1.107301e-08, 
    1.076996e-08, 1.054978e-08, 1.008403e-08, 9.368977e-09, 9.633313e-09, 
    9.152244e-09, 9.05785e-09, 9.790407e-09, 9.335581e-09, 1.085306e-08, 
    1.059632e-08, 1.074867e-08, 1.131865e-08, 9.571858e-09, 1.044131e-08, 
    8.878851e-09, 9.317879e-09, 8.08005e-09, 8.679134e-09, 7.532322e-09, 
    7.08367e-09, 6.674739e-09, 6.219874e-09, 1.088871e-08, 1.108638e-08, 
    1.073434e-08, 1.026086e-08, 9.835634e-09, 9.290639e-09, 9.236195e-09, 
    9.137069e-09, 8.884038e-09, 8.67535e-09, 9.105854e-09, 8.623619e-09, 
    1.053733e-08, 9.499027e-09, 1.116175e-08, 1.064009e-08, 1.028836e-08, 
    1.044162e-08, 9.663883e-09, 9.486997e-09, 8.792839e-09, 9.146798e-09, 
    7.188501e-09, 8.011346e-09, 5.889937e-09, 6.435147e-09, 1.115604e-08, 
    1.088941e-08, 9.997857e-09, 1.041506e-08, 9.255096e-09, 8.984923e-09, 
    8.769693e-09, 8.500137e-09, 8.471439e-09, 8.315083e-09, 8.57244e-09, 
    8.325152e-09, 9.289503e-09, 8.848803e-09, 1.009698e-08, 9.781848e-09, 
    9.925918e-09, 1.008572e-08, 9.598567e-09, 9.098945e-09, 9.088549e-09, 
    8.932644e-09, 8.503933e-09, 9.250603e-09, 7.092246e-09, 8.371835e-09, 
    1.060403e-08, 1.011338e-08, 1.004477e-08, 1.023185e-08, 9.011739e-09, 
    9.440578e-09, 8.318876e-09, 8.611653e-09, 8.135903e-09, 8.369775e-09, 
    8.404601e-09, 8.713288e-09, 8.909685e-09, 9.420577e-09, 9.852085e-09, 
    1.020457e-08, 1.012179e-08, 9.73743e-09, 9.06904e-09, 8.468815e-09, 
    8.597671e-09, 8.171351e-09, 9.335814e-09, 8.833377e-09, 9.025097e-09, 
    8.531599e-09, 9.640397e-09, 8.689667e-09, 9.895304e-09, 9.78492e-09, 
    9.449242e-09, 8.800003e-09, 8.661073e-09, 8.514436e-09, 8.604711e-09, 
    9.052541e-09, 9.127563e-09, 9.457314e-09, 9.549864e-09, 9.80888e-09, 
    1.00272e-08, 9.827572e-09, 9.621102e-09, 9.052375e-09, 8.561621e-09, 
    8.04956e-09, 7.927852e-09, 7.365511e-09, 7.820833e-09, 7.085505e-09, 
    7.706216e-09, 6.651702e-09, 8.636899e-09, 7.725349e-09, 9.434196e-09, 
    9.23771e-09, 8.890007e-09, 8.129624e-09, 8.533872e-09, 8.062584e-09, 
    9.130517e-09, 9.724332e-09, 9.88261e-09, 1.018286e-08, 9.875824e-09, 
    9.900539e-09, 9.612667e-09, 9.704493e-09, 9.033934e-09, 9.389693e-09, 
    8.405461e-09, 8.066244e-09, 7.163815e-09, 6.653634e-09, 6.158519e-09, 
    5.949164e-09, 5.886551e-09, 5.860525e-09,
  8.754804e-11, 7.986251e-11, 8.131317e-11, 7.542875e-11, 7.864975e-11, 
    7.485915e-11, 8.594481e-11, 7.956854e-11, 8.359414e-11, 8.683356e-11, 
    6.498139e-11, 7.517446e-11, 5.561129e-11, 6.122406e-11, 4.793569e-11, 
    5.645553e-11, 4.635503e-11, 4.816603e-11, 4.288976e-11, 4.434876e-11, 
    3.814695e-11, 4.223029e-11, 3.207231e-11, 3.909004e-11, 3.846428e-11, 
    4.237108e-11, 7.302719e-11, 6.618578e-11, 7.344951e-11, 7.243601e-11, 
    7.288954e-11, 7.858187e-11, 8.158113e-11, 8.815922e-11, 8.693501e-11, 
    8.211856e-11, 7.198395e-11, 7.53058e-11, 6.71614e-11, 6.733716e-11, 
    5.910428e-11, 6.270855e-11, 5.012743e-11, 5.346995e-11, 4.428704e-11, 
    4.646133e-11, 4.438713e-11, 4.50077e-11, 4.437909e-11, 4.760395e-11, 
    4.619886e-11, 4.912336e-11, 6.202014e-11, 5.797079e-11, 7.072661e-11, 
    7.942295e-11, 8.565678e-11, 9.030991e-11, 8.964024e-11, 8.837434e-11, 
    8.2091e-11, 7.651241e-11, 7.246743e-11, 6.985854e-11, 6.736246e-11, 
    6.024125e-11, 5.672932e-11, 4.947288e-11, 5.07226e-11, 4.862103e-11, 
    4.66825e-11, 4.357376e-11, 4.40731e-11, 4.274735e-11, 4.867586e-11, 
    4.466347e-11, 5.144601e-11, 4.951056e-11, 6.669417e-11, 7.439791e-11, 
    7.787859e-11, 8.103261e-11, 8.912798e-11, 8.347236e-11, 8.566684e-11, 
    8.051995e-11, 7.737896e-11, 7.892013e-11, 6.978828e-11, 7.323198e-11, 
    5.652654e-11, 6.329436e-11, 4.690521e-11, 5.046401e-11, 4.60843e-11, 
    4.827763e-11, 4.457119e-11, 4.789568e-11, 4.226283e-11, 4.111382e-11, 
    4.189605e-11, 3.895983e-11, 4.808586e-11, 4.438698e-11, 7.896354e-11, 
    7.871041e-11, 7.75399e-11, 8.279038e-11, 8.312064e-11, 8.819283e-11, 
    8.366824e-11, 8.179801e-11, 7.720013e-11, 7.457853e-11, 7.215305e-11, 
    6.704249e-11, 6.168418e-11, 5.478179e-11, 5.022666e-11, 4.735332e-11, 
    4.909853e-11, 4.755501e-11, 4.928314e-11, 5.011109e-11, 4.154107e-11, 
    4.618582e-11, 3.937091e-11, 3.972414e-11, 4.271618e-11, 3.968421e-11, 
    7.853309e-11, 7.999593e-11, 8.524281e-11, 8.111425e-11, 8.875967e-11, 
    8.44127e-11, 8.199044e-11, 7.31581e-11, 7.132411e-11, 6.965593e-11, 
    6.6454e-11, 6.251982e-11, 5.607687e-11, 5.092492e-11, 4.657182e-11, 
    4.687983e-11, 4.677119e-11, 4.583914e-11, 4.817673e-11, 4.546468e-11, 
    4.502222e-11, 4.61866e-11, 3.977165e-11, 4.152151e-11, 3.973168e-11, 
    4.086273e-11, 7.951814e-11, 7.708079e-11, 7.839029e-11, 7.59422e-11, 
    7.766024e-11, 7.025149e-11, 6.814441e-11, 5.895291e-11, 6.259528e-11, 
    5.688176e-11, 6.199456e-11, 6.106216e-11, 5.670199e-11, 6.170916e-11, 
    5.119802e-11, 5.814645e-11, 4.580324e-11, 5.213438e-11, 4.542898e-11, 
    4.658995e-11, 4.468126e-11, 4.302824e-11, 4.102317e-11, 3.753327e-11, 
    3.831773e-11, 3.555078e-11, 7.355844e-11, 7.059931e-11, 7.085638e-11, 
    6.785433e-11, 6.570067e-11, 6.122287e-11, 5.456233e-11, 5.699356e-11, 
    5.25968e-11, 5.174874e-11, 5.84558e-11, 5.425782e-11, 6.867321e-11, 
    6.615394e-11, 6.764506e-11, 7.332119e-11, 5.642505e-11, 6.464831e-11, 
    5.015404e-11, 5.409665e-11, 4.326066e-11, 4.839597e-11, 3.875554e-11, 
    3.201886e-11, 2.964212e-11, 2.70291e-11, 6.902559e-11, 7.09898e-11, 
    6.750437e-11, 6.291034e-11, 5.887914e-11, 5.384897e-11, 5.335513e-11, 
    5.246013e-11, 5.020001e-11, 4.836288e-11, 5.21794e-11, 4.791131e-11, 
    6.557962e-11, 5.575386e-11, 7.174358e-11, 6.658121e-11, 6.31741e-11, 
    6.46513e-11, 5.727711e-11, 5.564325e-11, 4.939414e-11, 5.254774e-11, 
    3.60252e-11, 4.268539e-11, 2.515546e-11, 2.826158e-11, 7.168646e-11, 
    6.903249e-11, 6.040624e-11, 6.439448e-11, 5.35264e-11, 5.109689e-11, 
    4.919036e-11, 4.683963e-11, 4.659182e-11, 4.525016e-11, 4.746607e-11, 
    4.533613e-11, 5.383866e-11, 4.98881e-11, 6.134595e-11, 5.837581e-11, 
    5.972738e-11, 6.12389e-11, 5.667189e-11, 5.211734e-11, 5.202401e-11, 
    5.063142e-11, 4.687243e-11, 5.348566e-11, 3.206897e-11, 4.573548e-11, 
    6.622919e-11, 6.150184e-11, 6.085037e-11, 6.263239e-11, 5.133624e-11, 
    5.521723e-11, 4.528255e-11, 4.780707e-11, 4.373044e-11, 4.571783e-11, 
    4.601654e-11, 4.869502e-11, 5.042747e-11, 5.503402e-11, 5.90334e-11, 
    6.237141e-11, 6.158191e-11, 5.796126e-11, 5.184901e-11, 4.656919e-11, 
    4.768538e-11, 4.402958e-11, 5.425994e-11, 4.975177e-11, 5.145561e-11, 
    4.711185e-11, 5.705923e-11, 4.848813e-11, 5.943929e-11, 5.840452e-11, 
    5.529666e-11, 4.945726e-11, 4.82381e-11, 4.696327e-11, 4.774664e-11, 
    5.170118e-11, 5.237459e-11, 5.537069e-11, 5.622206e-11, 5.862859e-11, 
    6.068385e-11, 5.88036e-11, 5.688044e-11, 5.169969e-11, 4.737213e-11, 
    4.300501e-11, 4.199014e-11, 3.742121e-11, 4.110528e-11, 3.202958e-11, 
    4.01655e-11, 2.950899e-11, 4.802709e-11, 4.032181e-11, 5.515874e-11, 
    5.336885e-11, 5.025292e-11, 4.367754e-11, 4.713153e-11, 4.311415e-11, 
    5.240116e-11, 5.783921e-11, 5.931997e-11, 6.216407e-11, 5.925622e-11, 
    5.948852e-11, 5.680235e-11, 5.765453e-11, 5.153463e-11, 5.475154e-11, 
    4.602392e-11, 4.314483e-11, 3.583216e-11, 2.952015e-11, 2.667925e-11, 
    2.549039e-11, 2.513633e-11, 2.498936e-11,
  8.438737e-14, 7.197421e-14, 7.428549e-14, 6.50088e-14, 7.005396e-14, 
    6.412518e-14, 8.176464e-14, 7.150774e-14, 7.795022e-14, 8.321648e-14, 
    4.925327e-14, 6.4614e-14, 3.606518e-14, 4.38453e-14, 2.610349e-14, 
    3.721082e-14, 2.416485e-14, 2.638948e-14, 2.006977e-14, 2.176687e-14, 
    1.485465e-14, 1.931626e-14, 1.189426e-14, 1.58523e-14, 1.518802e-14, 
    1.947639e-14, 6.130148e-14, 5.101776e-14, 6.194994e-14, 6.039628e-14, 
    6.109045e-14, 6.99468e-14, 7.471409e-14, 8.539161e-14, 8.338253e-14, 
    7.557525e-14, 5.970614e-14, 6.481785e-14, 5.245762e-14, 5.2718e-14, 
    4.08628e-14, 4.596395e-14, 2.88591e-14, 3.320134e-14, 2.169426e-14, 
    2.429389e-14, 2.181205e-14, 2.254647e-14, 2.180258e-14, 2.569315e-14, 
    2.397561e-14, 2.758727e-14, 4.497846e-14, 3.928954e-14, 5.779597e-14, 
    7.127694e-14, 8.129526e-14, 8.894426e-14, 8.783494e-14, 8.574565e-14, 
    7.553105e-14, 6.669708e-14, 6.044432e-14, 5.648537e-14, 5.27555e-14, 
    4.24561e-14, 3.75843e-14, 2.802822e-14, 2.962027e-14, 2.695694e-14, 
    2.4563e-14, 2.086032e-14, 2.144313e-14, 1.990632e-14, 2.702555e-14, 
    2.213821e-14, 3.055262e-14, 2.807587e-14, 5.17669e-14, 6.341164e-14, 
    6.88387e-14, 7.383729e-14, 8.698826e-14, 7.775363e-14, 8.131164e-14, 
    7.301979e-14, 6.80538e-14, 7.04811e-14, 5.637959e-14, 6.161573e-14, 
    3.73076e-14, 4.680657e-14, 2.483483e-14, 2.928889e-14, 2.383707e-14, 
    2.652836e-14, 2.202913e-14, 2.605391e-14, 1.935322e-14, 1.806065e-14, 
    1.893767e-14, 1.571333e-14, 2.628985e-14, 2.181187e-14, 7.054975e-14, 
    7.014974e-14, 6.830642e-14, 7.665466e-14, 7.718646e-14, 8.544692e-14, 
    7.806989e-14, 7.506136e-14, 6.777332e-14, 6.369085e-14, 5.996408e-14, 
    5.228164e-14, 4.449939e-14, 3.494855e-14, 2.898563e-14, 2.538435e-14, 
    2.755602e-14, 2.563276e-14, 2.778861e-14, 2.883826e-14, 1.853811e-14, 
    2.395984e-14, 1.615337e-14, 1.653454e-14, 1.98706e-14, 1.649131e-14, 
    6.986982e-14, 7.218615e-14, 8.062159e-14, 7.396765e-14, 8.638055e-14, 
    7.927423e-14, 7.536976e-14, 6.150233e-14, 5.870197e-14, 5.618046e-14, 
    5.141268e-14, 4.569327e-14, 3.669585e-14, 2.988025e-14, 2.442823e-14, 
    2.480382e-14, 2.467115e-14, 2.354138e-14, 2.640279e-14, 2.309176e-14, 
    2.256373e-14, 2.396078e-14, 1.658602e-14, 1.851617e-14, 1.65427e-14, 
    1.778184e-14, 7.142782e-14, 6.758629e-14, 6.964457e-14, 6.580754e-14, 
    6.849544e-14, 5.70778e-14, 5.391768e-14, 4.065181e-14, 4.580145e-14, 
    3.779267e-14, 4.494194e-14, 4.36157e-14, 3.754699e-14, 4.453497e-14, 
    3.023213e-14, 3.953233e-14, 2.349816e-14, 3.144692e-14, 2.304903e-14, 
    2.445029e-14, 2.215926e-14, 2.022908e-14, 1.795984e-14, 1.421674e-14, 
    1.503377e-14, 1.221993e-14, 6.211744e-14, 5.760334e-14, 5.799247e-14, 
    5.348587e-14, 5.030531e-14, 4.38436e-14, 3.465464e-14, 3.794566e-14, 
    3.205152e-14, 3.094506e-14, 3.996084e-14, 3.424789e-14, 5.470689e-14, 
    5.097093e-14, 5.317485e-14, 6.175275e-14, 3.71693e-14, 4.876787e-14, 
    2.889301e-14, 3.403311e-14, 2.049732e-14, 2.667584e-14, 1.549608e-14, 
    1.182557e-14, 8.950261e-15, 6.213805e-15, 5.523426e-14, 5.819465e-14, 
    5.296599e-14, 4.625378e-14, 4.054909e-14, 3.370375e-14, 3.304952e-14, 
    3.18725e-14, 2.895162e-14, 2.663458e-14, 3.150565e-14, 2.607328e-14, 
    5.012789e-14, 3.6258e-14, 5.933989e-14, 5.160023e-14, 4.663329e-14, 
    4.877222e-14, 3.833438e-14, 3.610839e-14, 2.792872e-14, 3.198722e-14, 
    1.268861e-14, 1.983533e-14, 4.543957e-15, 7.44705e-15, 5.925293e-14, 
    5.524459e-14, 4.268855e-14, 4.839873e-14, 3.327603e-14, 3.010169e-14, 
    2.767166e-14, 2.47547e-14, 2.445256e-14, 2.283532e-14, 2.552313e-14, 
    2.293798e-14, 3.369004e-14, 2.855453e-14, 4.401835e-14, 3.984993e-14, 
    4.173414e-14, 4.386635e-14, 3.750588e-14, 3.14247e-14, 3.130307e-14, 
    2.95033e-14, 2.479477e-14, 3.322212e-14, 1.188996e-14, 2.341665e-14, 
    5.108164e-14, 4.42399e-14, 4.331581e-14, 4.585466e-14, 3.041064e-14, 
    3.553359e-14, 2.287397e-14, 2.594419e-14, 2.104269e-14, 2.339544e-14, 
    2.375524e-14, 2.704953e-14, 2.924215e-14, 3.528713e-14, 4.076397e-14, 
    4.548069e-14, 4.435381e-14, 3.927637e-14, 3.107535e-14, 2.442502e-14, 
    2.579371e-14, 2.139214e-14, 3.425072e-14, 2.838142e-14, 3.056504e-14, 
    2.508781e-14, 3.803559e-14, 2.679084e-14, 4.133072e-14, 3.988972e-14, 
    3.564058e-14, 2.800848e-14, 2.647914e-14, 2.490585e-14, 2.586942e-14, 
    3.088332e-14, 3.17606e-14, 3.574038e-14, 3.689309e-14, 4.020068e-14, 
    4.308037e-14, 4.044398e-14, 3.779086e-14, 3.088139e-14, 2.540748e-14, 
    2.020234e-14, 1.904402e-14, 1.410125e-14, 1.805114e-14, 1.183933e-14, 
    1.701469e-14, 8.799819e-15, 2.621687e-14, 1.718576e-14, 3.545486e-14, 
    3.306766e-14, 2.901913e-14, 2.098106e-14, 2.511195e-14, 2.032811e-14, 
    3.179535e-14, 3.91079e-14, 4.116391e-14, 4.518407e-14, 4.107485e-14, 
    4.139958e-14, 3.768409e-14, 3.885333e-14, 3.066736e-14, 3.4908e-14, 
    2.376416e-14, 2.036351e-14, 1.24972e-14, 8.812388e-15, 5.882963e-15, 
    4.823848e-15, 4.528222e-15, 4.408221e-15,
  2.852239e-19, 2.437973e-19, 2.515189e-19, 2.20503e-19, 2.373792e-19, 
    2.175452e-19, 2.764797e-19, 2.422385e-19, 2.637543e-19, 2.813207e-19, 
    1.676608e-19, 2.191816e-19, 1.232317e-19, 1.494668e-19, 8.952008e-20, 
    1.270998e-19, 8.29395e-20, 9.049022e-20, 6.901307e-20, 7.478908e-20, 
    5.121714e-20, 6.644631e-20, 4.111687e-20, 5.462748e-20, 5.235708e-20, 
    6.69919e-20, 2.08089e-19, 1.735903e-19, 2.102612e-19, 2.050561e-19, 
    2.07382e-19, 2.37021e-19, 2.529503e-19, 2.885709e-19, 2.818743e-19, 
    2.558261e-19, 2.027434e-19, 2.198639e-19, 1.784266e-19, 1.793009e-19, 
    1.394186e-19, 1.565984e-19, 9.886152e-20, 1.135553e-19, 7.454209e-20, 
    8.337776e-20, 7.494273e-20, 7.744018e-20, 7.491054e-20, 8.812782e-20, 
    8.229677e-20, 9.455178e-20, 1.532818e-19, 1.341138e-19, 1.963399e-19, 
    2.414672e-19, 2.749143e-19, 3.004064e-19, 2.967116e-19, 2.897507e-19, 
    2.556785e-19, 2.261526e-19, 2.052171e-19, 1.919446e-19, 1.794268e-19, 
    1.447878e-19, 1.283604e-19, 9.604631e-20, 1.014395e-19, 9.241472e-20, 
    8.429162e-20, 7.170451e-20, 7.368774e-20, 6.845643e-20, 9.264736e-20, 
    7.605202e-20, 1.045959e-19, 9.620778e-20, 1.761068e-19, 2.151563e-19, 
    2.333159e-19, 2.500218e-19, 2.938911e-19, 2.630982e-19, 2.749689e-19, 
    2.472909e-19, 2.30691e-19, 2.388071e-19, 1.915898e-19, 2.091417e-19, 
    1.274265e-19, 1.594333e-19, 8.521455e-20, 1.003173e-19, 8.182616e-20, 
    9.096127e-20, 7.568107e-20, 8.935186e-20, 6.657227e-20, 6.216604e-20, 
    6.515618e-20, 5.415262e-20, 9.015227e-20, 7.494212e-20, 2.390365e-19, 
    2.376993e-19, 2.315358e-19, 2.594299e-19, 2.612051e-19, 2.887552e-19, 
    2.641537e-19, 2.541101e-19, 2.297529e-19, 2.160912e-19, 2.036078e-19, 
    1.778356e-19, 1.516691e-19, 1.194598e-19, 9.929013e-20, 8.707985e-20, 
    9.444583e-20, 8.79229e-20, 9.523423e-20, 9.879094e-20, 6.379415e-20, 
    8.224318e-20, 5.565607e-20, 5.695791e-20, 6.833476e-20, 5.681027e-20, 
    2.367636e-19, 2.445056e-19, 2.726674e-19, 2.504573e-19, 2.918663e-19, 
    2.681724e-19, 2.551399e-19, 2.087618e-19, 1.993775e-19, 1.909217e-19, 
    1.74917e-19, 1.556875e-19, 1.253613e-19, 1.023198e-19, 8.383396e-20, 
    8.510927e-20, 8.465883e-20, 8.082159e-20, 9.053537e-20, 7.929373e-20, 
    7.749886e-20, 8.224637e-20, 5.713369e-20, 6.371933e-20, 5.698578e-20, 
    6.121501e-20, 2.419714e-19, 2.291273e-19, 2.360105e-19, 2.231762e-19, 
    2.32168e-19, 1.939316e-19, 1.833286e-19, 1.387073e-19, 1.560516e-19, 
    1.290636e-19, 1.531588e-19, 1.486937e-19, 1.282345e-19, 1.517889e-19, 
    1.035111e-19, 1.349327e-19, 8.067474e-20, 1.076222e-19, 7.914849e-20, 
    8.390888e-20, 7.612359e-20, 6.955557e-20, 6.182218e-20, 4.903486e-20, 
    5.182965e-20, 4.219469e-20, 2.108222e-19, 1.95694e-19, 1.969988e-19, 
    1.818791e-19, 1.711965e-19, 1.494611e-19, 1.184667e-19, 1.295799e-19, 
    1.096673e-19, 1.059241e-19, 1.363777e-19, 1.170923e-19, 1.859775e-19, 
    1.734329e-19, 1.808349e-19, 2.096007e-19, 1.269596e-19, 1.66029e-19, 
    9.897641e-20, 1.163665e-19, 7.046886e-20, 9.146147e-20, 5.341015e-20, 
    4.088101e-20, 3.099039e-20, 2.153799e-20, 1.877472e-19, 1.976767e-19, 
    1.801336e-19, 1.575736e-19, 1.383611e-19, 1.152534e-19, 1.130421e-19, 
    1.090619e-19, 9.917496e-20, 9.132153e-20, 1.078208e-19, 8.941757e-20, 
    1.706003e-19, 1.238829e-19, 2.015158e-19, 1.75547e-19, 1.588504e-19, 
    1.660437e-19, 1.308916e-19, 1.233776e-19, 9.570908e-20, 1.094499e-19, 
    4.380149e-20, 6.821461e-20, 1.574461e-20, 2.58033e-20, 2.012244e-19, 
    1.877819e-19, 1.455709e-19, 1.647879e-19, 1.138078e-19, 1.030695e-19, 
    9.483781e-20, 8.494251e-20, 8.39166e-20, 7.842212e-20, 8.755085e-20, 
    7.877108e-20, 1.152071e-19, 9.782971e-20, 1.500495e-19, 1.360037e-19, 
    1.423553e-19, 1.495377e-19, 1.280957e-19, 1.07547e-19, 1.071355e-19, 
    1.010434e-19, 8.507854e-20, 1.136255e-19, 4.11021e-20, 8.039779e-20, 
    1.738049e-19, 1.507955e-19, 1.476837e-19, 1.562306e-19, 1.041153e-19, 
    1.214363e-19, 7.855351e-20, 8.897961e-20, 7.232516e-20, 8.032572e-20, 
    8.154816e-20, 9.272869e-20, 1.00159e-19, 1.206037e-19, 1.390854e-19, 
    1.549721e-19, 1.51179e-19, 1.340694e-19, 1.063649e-19, 8.382308e-20, 
    8.846902e-20, 7.351426e-20, 1.171018e-19, 9.724318e-20, 1.04638e-19, 
    8.607334e-20, 1.298834e-19, 9.185147e-20, 1.409957e-19, 1.361379e-19, 
    1.217977e-19, 9.59794e-20, 9.079434e-20, 8.545565e-20, 8.872594e-20, 
    1.057151e-19, 1.086833e-19, 1.221347e-19, 1.260272e-19, 1.371864e-19, 
    1.468907e-19, 1.380067e-19, 1.290575e-19, 1.057086e-19, 8.715837e-20, 
    6.94645e-20, 6.551862e-20, 4.86396e-20, 6.213361e-20, 4.092825e-20, 
    5.859721e-20, 3.047182e-20, 8.99047e-20, 5.91811e-20, 1.211704e-19, 
    1.131034e-19, 9.940361e-20, 7.211545e-20, 8.615529e-20, 6.989277e-20, 
    1.088009e-19, 1.335011e-19, 1.404335e-19, 1.539738e-19, 1.401334e-19, 
    1.412278e-19, 1.286972e-19, 1.326424e-19, 1.049843e-19, 1.193228e-19, 
    8.157846e-20, 7.001328e-20, 4.314536e-20, 3.051515e-20, 2.039195e-20, 
    1.671733e-20, 1.56899e-20, 1.527261e-20,
  2.093585e-25, 1.790998e-25, 1.847414e-25, 1.620751e-25, 1.744099e-25, 
    1.599128e-25, 2.029733e-25, 1.779608e-25, 1.936794e-25, 2.065084e-25, 
    1.234213e-25, 1.611091e-25, 9.087389e-26, 1.100992e-25, 6.613277e-26, 
    9.370971e-26, 6.12976e-26, 6.684542e-26, 5.105743e-26, 5.53059e-26, 
    3.79534e-26, 4.916881e-26, 3.051395e-26, 4.046652e-26, 3.879354e-26, 
    4.957029e-26, 1.529988e-25, 1.277614e-25, 1.545872e-25, 1.50781e-25, 
    1.524818e-25, 1.741481e-25, 1.857872e-25, 2.118023e-25, 2.069127e-25, 
    1.878881e-25, 1.490897e-25, 1.616079e-25, 1.313008e-25, 1.319406e-25, 
    1.027381e-25, 1.153221e-25, 7.29931e-26, 8.377708e-26, 5.512427e-26, 
    6.161969e-26, 5.541889e-26, 5.725523e-26, 5.539521e-26, 6.510995e-26, 
    6.082523e-26, 6.982851e-26, 1.128933e-25, 9.885077e-26, 1.444063e-25, 
    1.773972e-25, 2.018302e-25, 2.204429e-25, 2.177457e-25, 2.126637e-25, 
    1.877802e-25, 1.662048e-25, 1.508987e-25, 1.411912e-25, 1.320327e-25, 
    1.066718e-25, 9.463381e-26, 7.092601e-26, 7.488572e-26, 6.825899e-26, 
    6.229126e-26, 5.303733e-26, 5.449597e-26, 5.064788e-26, 6.842986e-26, 
    5.623458e-26, 7.720262e-26, 7.104458e-26, 1.296031e-25, 1.581662e-25, 
    1.714404e-25, 1.836477e-25, 2.156865e-25, 1.932002e-25, 2.018701e-25, 
    1.816524e-25, 1.69522e-25, 1.754534e-25, 1.409316e-25, 1.537686e-25, 
    9.39492e-26, 1.173979e-25, 6.296946e-26, 7.40619e-26, 6.047935e-26, 
    6.719142e-26, 5.596181e-26, 6.600919e-26, 4.92615e-26, 4.601841e-26, 
    4.821937e-26, 4.011665e-26, 6.659717e-26, 5.541844e-26, 1.75621e-25, 
    1.746439e-25, 1.701395e-25, 1.905206e-25, 1.918174e-25, 2.119369e-25, 
    1.939711e-25, 1.866345e-25, 1.688363e-25, 1.588497e-25, 1.497219e-25, 
    1.308683e-25, 1.117122e-25, 8.810809e-26, 7.330778e-26, 6.434002e-26, 
    6.975071e-26, 6.49594e-26, 7.032967e-26, 7.294128e-26, 4.721689e-26, 
    6.078584e-26, 4.122431e-26, 4.218328e-26, 5.055837e-26, 4.207453e-26, 
    1.7396e-25, 1.796173e-25, 2.001892e-25, 1.839658e-25, 2.142083e-25, 
    1.969064e-25, 1.873868e-25, 1.534908e-25, 1.46628e-25, 1.40443e-25, 
    1.287324e-25, 1.146551e-25, 9.243521e-26, 7.553191e-26, 6.195494e-26, 
    6.28921e-26, 6.256111e-26, 5.974098e-26, 6.687858e-26, 5.86179e-26, 
    5.729837e-26, 6.078819e-26, 4.231275e-26, 4.716182e-26, 4.220381e-26, 
    4.531825e-26, 1.777656e-25, 1.683791e-25, 1.734097e-25, 1.640292e-25, 
    1.706015e-25, 1.426447e-25, 1.348878e-25, 1.022169e-25, 1.149216e-25, 
    9.514929e-26, 1.128032e-25, 1.095329e-25, 9.45415e-26, 1.117999e-25, 
    7.640636e-26, 9.945088e-26, 5.963304e-26, 7.942364e-26, 5.851113e-26, 
    6.201e-26, 5.62872e-26, 5.145654e-26, 4.576526e-26, 3.63447e-26, 
    3.840484e-26, 3.129928e-26, 1.549974e-25, 1.439339e-25, 1.448882e-25, 
    1.338271e-25, 1.260093e-25, 1.10095e-25, 8.737982e-26, 9.552776e-26, 
    8.092442e-26, 7.817742e-26, 1.005098e-25, 8.637176e-26, 1.368258e-25, 
    1.276462e-25, 1.330631e-25, 1.541042e-25, 9.360696e-26, 1.222268e-25, 
    7.307745e-26, 8.583939e-26, 5.21284e-26, 6.755884e-26, 3.956957e-26, 
    3.033981e-26, 2.303062e-26, 1.602985e-26, 1.381206e-25, 1.453841e-25, 
    1.325499e-25, 1.160362e-25, 1.019632e-25, 8.502287e-26, 8.340054e-26, 
    8.048013e-26, 7.322322e-26, 6.745604e-26, 7.956944e-26, 6.605746e-26, 
    1.25573e-25, 9.135131e-26, 1.481919e-25, 1.291934e-25, 1.169711e-25, 
    1.222375e-25, 9.648918e-26, 9.098088e-26, 7.067837e-26, 8.076485e-26, 
    3.248493e-26, 5.046997e-26, 1.172844e-26, 1.919123e-26, 1.479788e-25, 
    1.38146e-25, 1.072454e-25, 1.213182e-25, 8.39623e-26, 7.608224e-26, 
    7.003856e-26, 6.276956e-26, 6.201567e-26, 5.797714e-26, 6.468607e-26, 
    5.823368e-26, 8.49889e-26, 7.223552e-26, 1.10526e-25, 1.002358e-25, 
    1.048897e-25, 1.101511e-25, 9.443981e-26, 7.936847e-26, 7.906647e-26, 
    7.459496e-26, 6.286951e-26, 8.382861e-26, 3.050304e-26, 5.942947e-26, 
    1.279185e-25, 1.110723e-25, 1.087931e-25, 1.150528e-25, 7.684989e-26, 
    8.955742e-26, 5.807373e-26, 6.573572e-26, 5.349384e-26, 5.937649e-26, 
    6.027503e-26, 6.848959e-26, 7.394566e-26, 8.894692e-26, 1.02494e-25, 
    1.141312e-25, 1.113532e-25, 9.881823e-26, 7.850097e-26, 6.194695e-26, 
    6.536063e-26, 5.436839e-26, 8.637877e-26, 7.180487e-26, 7.723348e-26, 
    6.360049e-26, 9.57502e-26, 6.784529e-26, 1.038936e-25, 1.003341e-25, 
    8.98224e-26, 7.087688e-26, 6.70688e-26, 6.314663e-26, 6.554937e-26, 
    7.802408e-26, 8.020235e-26, 9.006956e-26, 9.292341e-26, 1.011024e-25, 
    1.082123e-25, 1.017035e-25, 9.514483e-26, 7.801928e-26, 6.439771e-26, 
    5.138954e-26, 4.848611e-26, 3.605327e-26, 4.599454e-26, 3.037469e-26, 
    4.339064e-26, 2.264699e-26, 6.641531e-26, 4.382063e-26, 8.936241e-26, 
    8.344551e-26, 7.339109e-26, 5.333959e-26, 6.366071e-26, 5.170461e-26, 
    8.028861e-26, 9.840176e-26, 1.034817e-25, 1.134001e-25, 1.032618e-25, 
    1.040637e-25, 9.48807e-26, 9.77724e-26, 7.748766e-26, 8.800762e-26, 
    6.029729e-26, 5.179326e-26, 3.20008e-26, 2.267905e-26, 1.517969e-26, 
    1.245136e-26, 1.168777e-26, 1.137754e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.0112758, 0.01128991, 0.01128716, 0.01129854, 0.01129222, 0.01129968, 
    0.01127865, 0.01129049, 0.01128293, 0.01127705, 0.0113206, 0.01129905, 
    0.01134276, 0.01132911, 0.01136331, 0.01134066, 0.01136786, 0.01136262, 
    0.01137828, 0.0113738, 0.01139384, 0.01138035, 0.01140415, 0.0113906, 
    0.01139274, 0.01137991, 0.01130336, 0.01131793, 0.0113025, 0.01130458, 
    0.01130364, 0.01129237, 0.01128669, 0.0112747, 0.01127687, 0.01128567, 
    0.01130552, 0.01129877, 0.0113157, 0.01131532, 0.01133413, 0.01132566, 
    0.01135716, 0.01134822, 0.01137398, 0.01136752, 0.01137369, 0.01137181, 
    0.01137371, 0.01136423, 0.01136829, 0.01135993, 0.01132725, 0.01133689, 
    0.01130812, 0.01129079, 0.01127918, 0.01127094, 0.01127211, 0.01127433, 
    0.01128572, 0.01129638, 0.0113045, 0.01130993, 0.01131526, 0.01133148, 
    0.01133997, 0.01135898, 0.01135553, 0.01136135, 0.01136688, 0.01137617, 
    0.01137464, 0.01137874, 0.01136118, 0.01137287, 0.01135356, 0.01135885, 
    0.01131682, 0.01130058, 0.01129376, 0.0112877, 0.01127301, 0.01128316, 
    0.01127916, 0.01128865, 0.01129468, 0.0112917, 0.01131007, 0.01130294, 
    0.01134047, 0.01132434, 0.01136623, 0.01135623, 0.01136862, 0.0113623, 
    0.01137314, 0.01136338, 0.01138025, 0.01138393, 0.01138142, 0.01139102, 
    0.01136284, 0.0113737, 0.01129162, 0.0112921, 0.01129437, 0.01128442, 
    0.01128381, 0.01127465, 0.01128279, 0.01128626, 0.01129503, 0.01130022, 
    0.01130515, 0.01131597, 0.01132805, 0.01134486, 0.01135688, 0.01136493, 
    0.01135999, 0.01136436, 0.01135948, 0.01135719, 0.01138256, 0.01136834, 
    0.01138964, 0.01138846, 0.01137884, 0.0113886, 0.01129245, 0.01128964, 
    0.01127992, 0.01128753, 0.01127365, 0.01128143, 0.01128592, 0.01130311, 
    0.01130686, 0.01131036, 0.01131725, 0.01132609, 0.01134157, 0.01135499, 
    0.01136719, 0.0113663, 0.01136661, 0.01136935, 0.01136259, 0.01137045, 
    0.01137178, 0.01136832, 0.01138831, 0.0113826, 0.01138844, 0.01138472, 
    0.01129055, 0.01129526, 0.01129272, 0.01129751, 0.01129414, 0.01130913, 
    0.01131362, 0.01133452, 0.01132593, 0.01133957, 0.01132731, 0.01132949, 
    0.01134006, 0.01132796, 0.01135427, 0.01133649, 0.01136945, 0.01135179, 
    0.01137056, 0.01136714, 0.01137279, 0.01137786, 0.01138421, 0.01139593, 
    0.01139322, 0.01140299, 0.01130228, 0.01130839, 0.01130783, 0.01131421, 
    0.01131892, 0.0113291, 0.01134541, 0.01133927, 0.0113505, 0.01135276, 
    0.01133568, 0.0113462, 0.01131246, 0.01131795, 0.01131466, 0.01130277, 
    0.01134071, 0.01132129, 0.01135708, 0.0113466, 0.01137714, 0.01136199, 
    0.01139173, 0.01140444, 0.01141628, 0.01143019, 0.0113117, 0.01130755, 
    0.01131496, 0.01132522, 0.01133467, 0.01134724, 0.01134851, 0.01135087, 
    0.01135695, 0.01136206, 0.01135164, 0.01136334, 0.01131926, 0.01134239, 
    0.011306, 0.01131701, 0.01132461, 0.01132126, 0.01133857, 0.01134264, 
    0.01135919, 0.01135063, 0.01140132, 0.01137896, 0.01144069, 0.01142352, 
    0.01130611, 0.01131168, 0.01133104, 0.01132183, 0.01134807, 0.01135452, 
    0.01135973, 0.01136643, 0.01136714, 0.0113711, 0.01136461, 0.01137083, 
    0.01134727, 0.01135781, 0.01132881, 0.01133589, 0.01133263, 0.01132906, 
    0.01134007, 0.01135181, 0.01135202, 0.01135579, 0.01136644, 0.01134817, 
    0.01140426, 0.01136975, 0.01131774, 0.01132848, 0.01132998, 0.01132583, 
    0.01135387, 0.01134373, 0.011371, 0.01136363, 0.01137568, 0.0113697, 
    0.01136882, 0.01136112, 0.01135633, 0.0113442, 0.0113343, 0.01132642, 
    0.01132826, 0.01133691, 0.01135251, 0.01136722, 0.011364, 0.01137477, 
    0.01134617, 0.0113582, 0.01135356, 0.01136563, 0.01133912, 0.0113618, 
    0.01133331, 0.01133581, 0.01134353, 0.01135904, 0.01136241, 0.01136607, 
    0.01136381, 0.01135291, 0.0113511, 0.01134333, 0.0113412, 0.01133526, 
    0.01133036, 0.01133485, 0.01133957, 0.0113529, 0.0113649, 0.01137794, 
    0.01138111, 0.01139638, 0.011384, 0.01140446, 0.01138713, 0.01141705, 
    0.01136307, 0.01138656, 0.01134387, 0.01134848, 0.01135684, 0.01137589, 
    0.01136558, 0.01137762, 0.01135103, 0.01133722, 0.0113336, 0.01132691, 
    0.01133375, 0.0113332, 0.01133974, 0.01133764, 0.01135334, 0.01134491, 
    0.01136881, 0.01137752, 0.01140198, 0.01141694, 0.01143207, 0.01143875, 
    0.01144078, 0.01144163,
  3.675845e-05, 3.68498e-05, 3.683201e-05, 3.690573e-05, 3.686477e-05, 
    3.691308e-05, 3.67769e-05, 3.68535e-05, 3.680456e-05, 3.676657e-05, 
    3.70495e-05, 3.690899e-05, 3.719479e-05, 3.710526e-05, 3.732969e-05, 
    3.718098e-05, 3.73596e-05, 3.732521e-05, 3.742819e-05, 3.739869e-05, 
    3.753063e-05, 3.744179e-05, 3.75986e-05, 3.750932e-05, 3.752337e-05, 
    3.743889e-05, 3.693697e-05, 3.703203e-05, 3.693141e-05, 3.694489e-05, 
    3.69388e-05, 3.686568e-05, 3.682894e-05, 3.675134e-05, 3.67654e-05, 
    3.682232e-05, 3.695094e-05, 3.690718e-05, 3.701748e-05, 3.701497e-05, 
    3.713819e-05, 3.708266e-05, 3.728929e-05, 3.723058e-05, 3.739992e-05, 
    3.73574e-05, 3.739796e-05, 3.738564e-05, 3.739812e-05, 3.733574e-05, 
    3.736248e-05, 3.730751e-05, 3.70931e-05, 3.715625e-05, 3.696786e-05, 
    3.685548e-05, 3.67803e-05, 3.672704e-05, 3.673457e-05, 3.674897e-05, 
    3.682265e-05, 3.689171e-05, 3.694434e-05, 3.697969e-05, 3.701462e-05, 
    3.712074e-05, 3.717642e-05, 3.730125e-05, 3.727857e-05, 3.731685e-05, 
    3.735317e-05, 3.741431e-05, 3.740422e-05, 3.743119e-05, 3.731572e-05, 
    3.739254e-05, 3.726569e-05, 3.730043e-05, 3.702476e-05, 3.691896e-05, 
    3.68747e-05, 3.683546e-05, 3.674038e-05, 3.680609e-05, 3.678021e-05, 
    3.684163e-05, 3.688072e-05, 3.686136e-05, 3.698066e-05, 3.693424e-05, 
    3.717972e-05, 3.707398e-05, 3.734893e-05, 3.728321e-05, 3.736465e-05, 
    3.732308e-05, 3.739434e-05, 3.73302e-05, 3.744116e-05, 3.746537e-05, 
    3.744884e-05, 3.75121e-05, 3.732666e-05, 3.739802e-05, 3.686085e-05, 
    3.686401e-05, 3.687866e-05, 3.681424e-05, 3.681027e-05, 3.675099e-05, 
    3.680367e-05, 3.682615e-05, 3.688293e-05, 3.691662e-05, 3.694858e-05, 
    3.701924e-05, 3.70983e-05, 3.720852e-05, 3.728748e-05, 3.73404e-05, 
    3.730791e-05, 3.733659e-05, 3.730456e-05, 3.72895e-05, 3.745635e-05, 
    3.736277e-05, 3.7503e-05, 3.749523e-05, 3.743185e-05, 3.749611e-05, 
    3.686622e-05, 3.684804e-05, 3.678512e-05, 3.683436e-05, 3.674452e-05, 
    3.679491e-05, 3.682391e-05, 3.693535e-05, 3.695965e-05, 3.698254e-05, 
    3.702762e-05, 3.708551e-05, 3.718699e-05, 3.727505e-05, 3.735525e-05, 
    3.734936e-05, 3.735144e-05, 3.736941e-05, 3.732498e-05, 3.73767e-05, 
    3.738543e-05, 3.736268e-05, 3.749419e-05, 3.745664e-05, 3.749507e-05, 
    3.74706e-05, 3.685393e-05, 3.688448e-05, 3.686799e-05, 3.689903e-05, 
    3.687721e-05, 3.697447e-05, 3.70038e-05, 3.714074e-05, 3.708441e-05, 
    3.717385e-05, 3.709345e-05, 3.710774e-05, 3.717704e-05, 3.709775e-05, 
    3.727033e-05, 3.715362e-05, 3.737011e-05, 3.725401e-05, 3.737739e-05, 
    3.73549e-05, 3.739207e-05, 3.742541e-05, 3.746721e-05, 3.754444e-05, 
    3.752654e-05, 3.759097e-05, 3.692993e-05, 3.696962e-05, 3.696598e-05, 
    3.700768e-05, 3.703853e-05, 3.710519e-05, 3.721212e-05, 3.717189e-05, 
    3.72456e-05, 3.726043e-05, 3.714837e-05, 3.721731e-05, 3.699625e-05, 
    3.703214e-05, 3.701068e-05, 3.693313e-05, 3.718134e-05, 3.705402e-05, 
    3.728881e-05, 3.721995e-05, 3.742067e-05, 3.732106e-05, 3.751671e-05, 
    3.760049e-05, 3.767865e-05, 3.777053e-05, 3.699128e-05, 3.696416e-05, 
    3.70126e-05, 3.707979e-05, 3.714173e-05, 3.722418e-05, 3.723254e-05, 
    3.724801e-05, 3.728791e-05, 3.73215e-05, 3.725302e-05, 3.732991e-05, 
    3.704071e-05, 3.719232e-05, 3.695409e-05, 3.702603e-05, 3.707578e-05, 
    3.705384e-05, 3.716726e-05, 3.719402e-05, 3.730265e-05, 3.724644e-05, 
    3.757993e-05, 3.743262e-05, 3.783999e-05, 3.772651e-05, 3.695477e-05, 
    3.699113e-05, 3.71179e-05, 3.705759e-05, 3.722961e-05, 3.727194e-05, 
    3.730623e-05, 3.735023e-05, 3.735489e-05, 3.738092e-05, 3.733827e-05, 
    3.737919e-05, 3.722436e-05, 3.729358e-05, 3.710328e-05, 3.714972e-05, 
    3.712831e-05, 3.710492e-05, 3.717711e-05, 3.725413e-05, 3.725558e-05, 
    3.728029e-05, 3.735023e-05, 3.72303e-05, 3.759928e-05, 3.737201e-05, 
    3.703083e-05, 3.710115e-05, 3.711095e-05, 3.708376e-05, 3.726771e-05, 
    3.720114e-05, 3.738026e-05, 3.733186e-05, 3.74111e-05, 3.737175e-05, 
    3.736597e-05, 3.731535e-05, 3.728387e-05, 3.720423e-05, 3.713931e-05, 
    3.708768e-05, 3.709967e-05, 3.715637e-05, 3.725879e-05, 3.73554e-05, 
    3.733428e-05, 3.740508e-05, 3.721716e-05, 3.729613e-05, 3.726568e-05, 
    3.7345e-05, 3.717087e-05, 3.731978e-05, 3.713282e-05, 3.71492e-05, 
    3.719982e-05, 3.730162e-05, 3.732382e-05, 3.734788e-05, 3.733299e-05, 
    3.726135e-05, 3.724952e-05, 3.719854e-05, 3.718456e-05, 3.714562e-05, 
    3.711345e-05, 3.714289e-05, 3.717383e-05, 3.72613e-05, 3.734014e-05, 
    3.742591e-05, 3.744681e-05, 3.754734e-05, 3.746579e-05, 3.760058e-05, 
    3.748641e-05, 3.768371e-05, 3.73281e-05, 3.748265e-05, 3.720205e-05, 
    3.723229e-05, 3.728717e-05, 3.741242e-05, 3.734462e-05, 3.742381e-05, 
    3.724904e-05, 3.715842e-05, 3.713471e-05, 3.709086e-05, 3.713572e-05, 
    3.713206e-05, 3.717497e-05, 3.716117e-05, 3.72642e-05, 3.720887e-05, 
    3.736588e-05, 3.742313e-05, 3.758429e-05, 3.768301e-05, 3.7783e-05, 
    3.78272e-05, 3.784063e-05, 3.784625e-05,
  8.749195e-10, 8.776447e-10, 8.771137e-10, 8.793142e-10, 8.780916e-10, 
    8.795339e-10, 8.754697e-10, 8.777549e-10, 8.762948e-10, 8.751617e-10, 
    8.836153e-10, 8.794117e-10, 8.879733e-10, 8.852877e-10, 8.920253e-10, 
    8.875585e-10, 8.929429e-10, 8.918909e-10, 8.950742e-10, 8.941576e-10, 
    8.982592e-10, 8.954971e-10, 9.003755e-10, 8.975967e-10, 8.980336e-10, 
    8.954069e-10, 8.802477e-10, 8.830919e-10, 8.800816e-10, 8.80484e-10, 
    8.803023e-10, 8.781187e-10, 8.770216e-10, 8.747075e-10, 8.751267e-10, 
    8.768243e-10, 8.806649e-10, 8.793579e-10, 8.826571e-10, 8.825821e-10, 
    8.862754e-10, 8.846104e-10, 8.908115e-10, 8.890483e-10, 8.941958e-10, 
    8.928751e-10, 8.941347e-10, 8.937521e-10, 8.941397e-10, 8.922075e-10, 
    8.930328e-10, 8.913589e-10, 8.849234e-10, 8.86817e-10, 8.811709e-10, 
    8.778134e-10, 8.755709e-10, 8.739832e-10, 8.742077e-10, 8.746366e-10, 
    8.768343e-10, 8.788958e-10, 8.80468e-10, 8.815253e-10, 8.825713e-10, 
    8.857513e-10, 8.87422e-10, 8.911706e-10, 8.904896e-10, 8.916396e-10, 
    8.927435e-10, 8.946427e-10, 8.943294e-10, 8.951672e-10, 8.916058e-10, 
    8.939663e-10, 8.901028e-10, 8.911464e-10, 8.828741e-10, 8.797096e-10, 
    8.783875e-10, 8.772164e-10, 8.743806e-10, 8.763401e-10, 8.755681e-10, 
    8.774008e-10, 8.785676e-10, 8.779897e-10, 8.815543e-10, 8.801662e-10, 
    8.875211e-10, 8.843501e-10, 8.92612e-10, 8.90629e-10, 8.931001e-10, 
    8.918269e-10, 8.940224e-10, 8.920412e-10, 8.954774e-10, 8.962299e-10, 
    8.957161e-10, 8.976834e-10, 8.919347e-10, 8.941365e-10, 8.779744e-10, 
    8.780688e-10, 8.785063e-10, 8.765834e-10, 8.764648e-10, 8.746969e-10, 
    8.762683e-10, 8.769389e-10, 8.786338e-10, 8.796396e-10, 8.805944e-10, 
    8.827096e-10, 8.850788e-10, 8.883855e-10, 8.907573e-10, 8.923475e-10, 
    8.913713e-10, 8.922333e-10, 8.912703e-10, 8.908181e-10, 8.959492e-10, 
    8.930416e-10, 8.974004e-10, 8.971587e-10, 8.951878e-10, 8.971859e-10, 
    8.781347e-10, 8.775923e-10, 8.757147e-10, 8.771841e-10, 8.745042e-10, 
    8.760066e-10, 8.768716e-10, 8.80199e-10, 8.809256e-10, 8.816106e-10, 
    8.829609e-10, 8.846958e-10, 8.877394e-10, 8.903838e-10, 8.928083e-10, 
    8.926256e-10, 8.926901e-10, 8.93248e-10, 8.918841e-10, 8.934744e-10, 
    8.937456e-10, 8.930391e-10, 8.971264e-10, 8.959586e-10, 8.971536e-10, 
    8.963927e-10, 8.777681e-10, 8.7868e-10, 8.781876e-10, 8.791145e-10, 
    8.784629e-10, 8.813686e-10, 8.822471e-10, 8.863514e-10, 8.846626e-10, 
    8.873451e-10, 8.849337e-10, 8.853621e-10, 8.874403e-10, 8.850629e-10, 
    8.902415e-10, 8.867378e-10, 8.932697e-10, 8.897509e-10, 8.934959e-10, 
    8.927976e-10, 8.93952e-10, 8.949878e-10, 8.962871e-10, 8.986896e-10, 
    8.981326e-10, 9.001382e-10, 8.800375e-10, 8.812236e-10, 8.81115e-10, 
    8.823636e-10, 8.832877e-10, 8.85286e-10, 8.884941e-10, 8.872867e-10, 
    8.894992e-10, 8.899445e-10, 8.865811e-10, 8.886497e-10, 8.820211e-10, 
    8.830959e-10, 8.824534e-10, 8.801329e-10, 8.875697e-10, 8.837516e-10, 
    8.907972e-10, 8.887291e-10, 8.948405e-10, 8.917659e-10, 8.978268e-10, 
    9.004338e-10, 9.028701e-10, 9.057352e-10, 8.818724e-10, 8.810603e-10, 
    8.825111e-10, 8.845241e-10, 8.863816e-10, 8.88856e-10, 8.891072e-10, 
    8.895716e-10, 8.907702e-10, 8.917796e-10, 8.897218e-10, 8.920323e-10, 
    8.83352e-10, 8.878995e-10, 8.80759e-10, 8.829127e-10, 8.844039e-10, 
    8.837463e-10, 8.871479e-10, 8.879505e-10, 8.912128e-10, 8.895246e-10, 
    8.997935e-10, 8.952114e-10, 9.07904e-10, 9.043618e-10, 8.807798e-10, 
    8.818679e-10, 8.856668e-10, 8.838589e-10, 8.890192e-10, 8.902905e-10, 
    8.913207e-10, 8.926522e-10, 8.92797e-10, 8.936056e-10, 8.922836e-10, 
    8.935519e-10, 8.888612e-10, 8.909404e-10, 8.852286e-10, 8.866212e-10, 
    8.859794e-10, 8.852779e-10, 8.874432e-10, 8.897551e-10, 8.897989e-10, 
    8.90541e-10, 8.926505e-10, 8.8904e-10, 9.003952e-10, 8.933271e-10, 
    8.830571e-10, 8.851643e-10, 8.854585e-10, 8.846435e-10, 8.901633e-10, 
    8.881644e-10, 8.935851e-10, 8.92091e-10, 8.945431e-10, 8.933208e-10, 
    8.931412e-10, 8.915948e-10, 8.906488e-10, 8.882571e-10, 8.86309e-10, 
    8.84761e-10, 8.851206e-10, 8.868208e-10, 8.898952e-10, 8.928127e-10, 
    8.921633e-10, 8.94356e-10, 8.886454e-10, 8.910169e-10, 8.901022e-10, 
    8.9249e-10, 8.872558e-10, 8.917266e-10, 8.861146e-10, 8.866057e-10, 
    8.881247e-10, 8.911815e-10, 8.918493e-10, 8.925792e-10, 8.92125e-10, 
    8.899722e-10, 8.896169e-10, 8.880864e-10, 8.876666e-10, 8.864984e-10, 
    8.855337e-10, 8.864165e-10, 8.873445e-10, 8.899708e-10, 8.923396e-10, 
    8.950033e-10, 8.95653e-10, 8.987789e-10, 8.962421e-10, 9.004357e-10, 
    8.968822e-10, 9.030263e-10, 8.919773e-10, 8.967664e-10, 8.881919e-10, 
    8.890997e-10, 8.907474e-10, 8.945836e-10, 8.924783e-10, 8.949376e-10, 
    8.896026e-10, 8.868822e-10, 8.861713e-10, 8.848561e-10, 8.862013e-10, 
    8.860917e-10, 8.873791e-10, 8.869651e-10, 8.900579e-10, 8.883965e-10, 
    8.931382e-10, 8.949167e-10, 8.999301e-10, 9.030053e-10, 9.06125e-10, 
    9.075048e-10, 9.079242e-10, 9.080998e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.5863606, 0.5554544, 0.5614216, 0.5367937, 0.5504095, 0.5343481, 
    0.5800518, 0.5542405, 0.5706755, 0.583554, 0.4900863, 0.5357026, 
    0.4439954, 0.4718316, 0.4032978, 0.4482845, 0.3944923, 0.4045593, 
    0.3746237, 0.3830826, 0.3460884, 0.3707522, 0.3277075, 0.3518925, 
    0.3480474, 0.371582, 0.5264026, 0.4956877, 0.5282441, 0.5238189, 
    0.5258014, 0.5501295, 0.5625269, 0.5887381, 0.5839525, 0.5647107, 
    0.521833, 0.5362597, 0.5001519, 0.5009573, 0.4614896, 0.4789506, 
    0.4152465, 0.432953, 0.3827275, 0.395082, 0.3833045, 0.3868564, 
    0.3832583, 0.4014551, 0.3936084, 0.4098027, 0.4756621, 0.4558769, 
    0.516264, 0.553646, 0.5789137, 0.5970479, 0.5944747, 0.5895793, 
    0.5645988, 0.541408, 0.5239499, 0.5123821, 0.5010732, 0.4670787, 
    0.4496622, 0.4117098, 0.4184432, 0.4070625, 0.3963214, 0.3786096, 
    0.3814964, 0.3737936, 0.4073574, 0.3848933, 0.4223021, 0.4119084, 
    0.4980361, 0.5323536, 0.5471941, 0.5602739, 0.5924988, 0.5701893, 
    0.5789549, 0.5581622, 0.5450757, 0.5515348, 0.5120671, 0.5272946, 
    0.4486385, 0.4817396, 0.397567, 0.4170566, 0.3929611, 0.4051707, 
    0.3843631, 0.4030659, 0.3709458, 0.3641331, 0.368782, 0.3510891, 
    0.4041157, 0.3833063, 0.5517173, 0.5506622, 0.5457526, 0.5674367, 
    0.5687703, 0.5888706, 0.5709732, 0.5634033, 0.5443183, 0.5331334, 
    0.5225716, 0.4996094, 0.4740531, 0.4397457, 0.4157803, 0.4000612, 
    0.409665, 0.4011807, 0.4106714, 0.4151545, 0.3666793, 0.3935368, 
    0.3536052, 0.3557558, 0.3736121, 0.3555131, 0.5499213, 0.5559998, 
    0.5772694, 0.5606033, 0.5910713, 0.5739613, 0.5641918, 0.5269796, 
    0.5189116, 0.511476, 0.4968987, 0.4780508, 0.4463571, 0.41953, 0.3956999, 
    0.3974231, 0.3968163, 0.3915785, 0.4046168, 0.3894577, 0.386943, 
    0.3935378, 0.3560445, 0.3665578, 0.3558016, 0.3626255, 0.554021, 
    0.543816, 0.5493233, 0.5389833, 0.5462631, 0.5141506, 0.5046545, 
    0.4607511, 0.4784127, 0.4504257, 0.4755372, 0.4710489, 0.4495332, 
    0.4741649, 0.4209937, 0.4567602, 0.3913756, 0.4259679, 0.389255, 
    0.3958016, 0.3849898, 0.3754354, 0.3635871, 0.3422612, 0.3471361, 
    0.3297083, 0.5287155, 0.5156983, 0.5168358, 0.5033222, 0.4934128, 
    0.4718218, 0.4386131, 0.4509813, 0.4283854, 0.423912, 0.4582804, 
    0.4370451, 0.5070471, 0.4955226, 0.5023695, 0.5276871, 0.4481235, 
    0.4885086, 0.41539, 0.4362077, 0.3767907, 0.4058296, 0.3498368, 
    0.3272588, 0.3067935, 0.2839237, 0.5086375, 0.5174284, 0.5017226, 
    0.4799194, 0.4603786, 0.4349257, 0.4323545, 0.427669, 0.4156342, 
    0.4056398, 0.4261958, 0.4031519, 0.492872, 0.444716, 0.5207695, 
    0.4974974, 0.4811692, 0.4885153, 0.4524032, 0.4441463, 0.4112806, 
    0.4281273, 0.3327545, 0.3734378, 0.2672762, 0.2947627, 0.5205134, 
    0.5086658, 0.4678684, 0.4873089, 0.4332467, 0.420446, 0.4101653, 
    0.3972031, 0.395813, 0.3882401, 0.4006872, 0.3887267, 0.4348722, 
    0.4139529, 0.4724143, 0.4578872, 0.4645461, 0.4718978, 0.4493604, 
    0.4258695, 0.4253677, 0.4179586, 0.3974153, 0.4330345, 0.3277029, 
    0.3910193, 0.495859, 0.473179, 0.470021, 0.4785852, 0.4217218, 0.4419738, 
    0.388423, 0.4025761, 0.3795156, 0.3908917, 0.3925797, 0.4074615, 
    0.4168604, 0.4410373, 0.4611405, 0.4773386, 0.4735518, 0.4558281, 
    0.4244493, 0.3956897, 0.4019091, 0.3812444, 0.4370506, 0.4132194, 
    0.4223608, 0.3987194, 0.4513134, 0.4063556, 0.4631329, 0.4580264, 
    0.44238, 0.4116289, 0.4049536, 0.3978936, 0.4022418, 0.4236644, 
    0.4272198, 0.442756, 0.4470909, 0.4591357, 0.4692101, 0.4600036, 
    0.450417, 0.4236527, 0.4001705, 0.3753011, 0.3693354, 0.3415741, 
    0.3640924, 0.3273686, 0.3584654, 0.3056584, 0.4038079, 0.3593924, 
    0.4416714, 0.4324254, 0.4159291, 0.3792208, 0.398829, 0.3759436, 
    0.4273589, 0.4552246, 0.4625473, 0.4763487, 0.4622337, 0.4633751, 
    0.4500174, 0.4542919, 0.4227764, 0.4395829, 0.3926238, 0.3761203, 
    0.3315127, 0.3057427, 0.2808206, 0.2702615, 0.2671022, 0.2657894,
  0.9312716, 0.9125664, 0.9161705, 0.9013243, 0.9095249, 0.8998544, 
    0.9274469, 0.9118322, 0.9217671, 0.9295714, 0.8733776, 0.9006687, 
    0.8115082, 0.8240206, 0.7935101, 0.8134243, 0.7896653, 0.7940651, 
    0.7810593, 0.7847124, 0.7688704, 0.7793934, 0.7611469, 0.7713328, 
    0.7697009, 0.7797499, 0.895086, 0.8767115, 0.8961908, 0.8935347, 
    0.8947253, 0.9093544, 0.916834, 0.932718, 0.9298131, 0.918157, 0.8923436, 
    0.9010065, 0.8793854, 0.8798658, 0.8193549, 0.8272456, 0.7987593, 
    0.806593, 0.7845588, 0.7899245, 0.7848081, 0.7863479, 0.7847881, 
    0.7927063, 0.7892821, 0.7963653, 0.8257544, 0.8168308, 0.8890093, 
    0.9114692, 0.926756, 0.9377666, 0.9362021, 0.9332268, 0.9180892, 
    0.9041032, 0.8936163, 0.8866889, 0.8799349, 0.8218686, 0.8140423, 
    0.7972016, 0.800169, 0.7951611, 0.7904649, 0.7827778, 0.7840258, 
    0.7807008, 0.7952921, 0.7854953, 0.8018736, 0.7972907, 0.87811, 0.898659, 
    0.9075803, 0.9154764, 0.935001, 0.9214711, 0.9267803, 0.9142035, 
    0.906311, 0.9102046, 0.8865005, 0.8956218, 0.8135843, 0.8285099, 
    0.7910081, 0.7995573, 0.7890008, 0.7943338, 0.785266, 0.7934119, 
    0.779476, 0.7765526, 0.778546, 0.7709932, 0.7938714, 0.7848081, 0.910314, 
    0.9096775, 0.9067194, 0.9198054, 0.9206128, 0.9327977, 0.9219475, 
    0.9173675, 0.9058561, 0.8991273, 0.8927888, 0.8790605, 0.8250245, 
    0.8096137, 0.7989947, 0.7920979, 0.7963055, 0.7925872, 0.7967473, 
    0.7987199, 0.7776432, 0.7892503, 0.772062, 0.7729772, 0.7806223, 
    0.7728739, 0.9092309, 0.9128984, 0.92576, 0.9156778, 0.9341345, 
    0.9237553, 0.9178421, 0.8954297, 0.8905967, 0.8861458, 0.8774456, 
    0.8268375, 0.8125653, 0.8006474, 0.7901943, 0.790946, 0.7906811, 
    0.7883989, 0.7940907, 0.787477, 0.7863843, 0.7892518, 0.7731001, 
    0.7775927, 0.7729968, 0.7759091, 0.9117044, 0.9055527, 0.9088708, 
    0.9026433, 0.9070252, 0.8877423, 0.8820662, 0.81902, 0.827001, 0.8143856, 
    0.8256986, 0.8236668, 0.8139819, 0.8250777, 0.8012919, 0.8172246, 
    0.7883106, 0.8034896, 0.7873889, 0.7902386, 0.7855387, 0.7814083, 
    0.7763201, 0.7672556, 0.7693166, 0.7619838, 0.8964747, 0.8886703, 
    0.8893541, 0.881276, 0.8753684, 0.8240174, 0.8091101, 0.8146366, 
    0.8045661, 0.8025846, 0.8179126, 0.8084111, 0.8834981, 0.8766211, 
    0.8807065, 0.8958557, 0.8133544, 0.8724473, 0.7988225, 0.8080396, 
    0.7819926, 0.79462, 0.770461, 0.7609575, 0.7524919, 0.7432099, 0.8844494, 
    0.8897089, 0.8803223, 0.8276826, 0.818855, 0.807469, 0.8063272, 
    0.8042479, 0.7989311, 0.7945392, 0.8035935, 0.7934496, 0.8750368, 
    0.8118318, 0.8917081, 0.877797, 0.8282509, 0.8724546, 0.8152744, 
    0.8115793, 0.7970133, 0.8044518, 0.7632552, 0.7805455, 0.7366009, 
    0.747582, 0.8915564, 0.8844676, 0.8222293, 0.8717377, 0.8067235, 
    0.8010525, 0.7965253, 0.7908486, 0.7902433, 0.7869477, 0.7923715, 
    0.7871597, 0.8074452, 0.7981902, 0.8242859, 0.8177348, 0.8207331, 
    0.8240522, 0.813911, 0.8034486, 0.8032291, 0.7999539, 0.7909326, 
    0.8066293, 0.7611382, 0.7881477, 0.8768266, 0.8246278, 0.823203, 
    0.8270806, 0.801616, 0.8106087, 0.7870275, 0.7931976, 0.7831697, 
    0.7881005, 0.7888346, 0.795338, 0.7994707, 0.8101904, 0.8191977, 
    0.8265156, 0.8248005, 0.8168092, 0.8028204, 0.7901886, 0.792904, 
    0.7839171, 0.8084152, 0.7978662, 0.8018972, 0.7915112, 0.8147848, 
    0.7948446, 0.8200963, 0.8177983, 0.81079, 0.7971649, 0.7942385, 0.79115, 
    0.7930514, 0.8024737, 0.8040485, 0.8109585, 0.8128941, 0.8182973, 
    0.8228376, 0.8186869, 0.8143824, 0.8024697, 0.7921442, 0.78135, 
    0.7787845, 0.7669619, 0.7765321, 0.7609982, 0.7741219, 0.7520207, 
    0.7937317, 0.7745223, 0.8104748, 0.8063589, 0.799058, 0.783039, 
    0.7915592, 0.7816253, 0.8041104, 0.8165368, 0.8198323, 0.8260664, 
    0.8196911, 0.8202053, 0.8142053, 0.8161216, 0.8020822, 0.8095434, 
    0.7888531, 0.7817022, 0.7627379, 0.7520587, 0.7419705, 0.7377772, 
    0.7365333, 0.7360179,
  1.172312, 1.17309, 1.172964, 1.173403, 1.173187, 1.173434, 1.172496, 
    1.173114, 1.172746, 1.172396, 1.173595, 1.173417, 1.212339, 1.218188, 
    1.203267, 1.213257, 1.201211, 1.20356, 1.196433, 1.198493, 1.189186, 
    1.195478, 1.18425, 1.190701, 1.1897, 1.195683, 1.173521, 1.17362, 
    1.173503, 1.173544, 1.173527, 1.173192, 1.17294, 1.17224, 1.172384, 
    1.17289, 1.17356, 1.17341, 1.173631, 1.173632, 1.216046, 1.219642, 
    1.206003, 1.209946, 1.198407, 1.201351, 1.198546, 1.199399, 1.198534, 
    1.202841, 1.201004, 1.204766, 1.218972, 1.214869, 1.173597, 1.173126, 
    1.172528, 1.171973, 1.172058, 1.172214, 1.172893, 1.173337, 1.173543, 
    1.173615, 1.173632, 1.217204, 1.213551, 1.205199, 1.206725, 1.204136, 
    1.201643, 1.197408, 1.198109, 1.196228, 1.204205, 1.198927, 1.20759, 
    1.205246, 1.173626, 1.173458, 1.173244, 1.17299, 1.172122, 1.172758, 
    1.172527, 1.173035, 1.173279, 1.173166, 1.173616, 1.173513, 1.213333, 
    1.220207, 1.201935, 1.206413, 1.200851, 1.203702, 1.1988, 1.203216, 
    1.195525, 1.193824, 1.194988, 1.190494, 1.203459, 1.198545, 1.173163, 
    1.173182, 1.173268, 1.172826, 1.172793, 1.172236, 1.172738, 1.17292, 
    1.173292, 1.173449, 1.173555, 1.17363, 1.218642, 1.211424, 1.206124, 
    1.202518, 1.204735, 1.202778, 1.204964, 1.205984, 1.194462, 1.200986, 
    1.191145, 1.191698, 1.196183, 1.191635, 1.173196, 1.173079, 1.172573, 
    1.172982, 1.172167, 1.172662, 1.172902, 1.173516, 1.173581, 1.173618, 
    1.173625, 1.219459, 1.212847, 1.206968, 1.201497, 1.201901, 1.201759, 
    1.200524, 1.203574, 1.20002, 1.199419, 1.200987, 1.191772, 1.194433, 
    1.19171, 1.193446, 1.173119, 1.1733, 1.173207, 1.173373, 1.17326, 
    1.173607, 1.173632, 1.215891, 1.219533, 1.213715, 1.218947, 1.218027, 
    1.213522, 1.218667, 1.207295, 1.215053, 1.200476, 1.208402, 1.199972, 
    1.201521, 1.198952, 1.196632, 1.193688, 1.188179, 1.189463, 1.1848, 
    1.173498, 1.1736, 1.173594, 1.173633, 1.173613, 1.218186, 1.211179, 
    1.213834, 1.208941, 1.207949, 1.215376, 1.210838, 1.17363, 1.17362, 
    1.173633, 1.173509, 1.213224, 1.173586, 1.206036, 1.210657, 1.196964, 
    1.203852, 1.190168, 1.184124, 1.178329, 1.171416, 1.173626, 1.17359, 
    1.173633, 1.219837, 1.215814, 1.210377, 1.209815, 1.208782, 1.206092, 
    1.20381, 1.208455, 1.203236, 1.173609, 1.212495, 1.173568, 1.173626, 
    1.220091, 1.173587, 1.214136, 1.212374, 1.205102, 1.208884, 1.185626, 
    1.196139, 1.166052, 1.174753, 1.17357, 1.173626, 1.217371, 1.173579, 
    1.21001, 1.207174, 1.204849, 1.201849, 1.201523, 1.199729, 1.202664, 
    1.199846, 1.210365, 1.205711, 1.218309, 1.215292, 1.216684, 1.218202, 
    1.21349, 1.208382, 1.208273, 1.206615, 1.201891, 1.209964, 1.184241, 
    1.200384, 1.173622, 1.218463, 1.217816, 1.219569, 1.20746, 1.211906, 
    1.199773, 1.203102, 1.197629, 1.200361, 1.200761, 1.204229, 1.206368, 
    1.211704, 1.215973, 1.219315, 1.218542, 1.214859, 1.208067, 1.201494, 
    1.202946, 1.198048, 1.21084, 1.205543, 1.207602, 1.202204, 1.213905, 
    1.203969, 1.21639, 1.215322, 1.211994, 1.20518, 1.203652, 1.202011, 
    1.203025, 1.207893, 1.208683, 1.212075, 1.213005, 1.215555, 1.217649, 
    1.215736, 1.213713, 1.207891, 1.202542, 1.196598, 1.195126, 1.187993, 
    1.193811, 1.184149, 1.192381, 1.177991, 1.203383, 1.192622, 1.211842, 
    1.209831, 1.206156, 1.197554, 1.20223, 1.196754, 1.208714, 1.214731, 
    1.216268, 1.219113, 1.216203, 1.21644, 1.21363, 1.214536, 1.207696, 
    1.21139, 1.200771, 1.196798, 1.185291, 1.178019, 1.170442, 1.167039, 
    1.165996, 1.165559,
  0.5064242, 0.4962063, 0.4981907, 0.4899655, 0.4945262, 0.4891436, 
    0.5043508, 0.4958009, 0.5012569, 0.5055038, 0.4740617, 0.4895992, 
    0.4580591, 0.4679053, 0.4432473, 0.4595882, 0.4399667, 0.4437181, 
    0.4324498, 0.4356719, 0.4213248, 0.4309645, 0.4139318, 0.4236231, 
    0.4221032, 0.4312831, 0.4864671, 0.4759914, 0.4870886, 0.4855924, 
    0.4862639, 0.4944316, 0.4985543, 0.507207, 0.5056349, 0.4992808, 
    0.4849198, 0.4897885, 0.4775348, 0.477811, 0.4642727, 0.4703916, 
    0.4476569, 0.4540975, 0.4355373, 0.4401901, 0.4357555, 0.4370993, 
    0.435738, 0.442566, 0.4396378, 0.4456561, 0.4692444, 0.4622885, 0.483032, 
    0.4955997, 0.5039753, 0.5099292, 0.509087, 0.5074816, 0.4992436, 
    0.4915162, 0.485639, 0.4817135, 0.4778507, 0.4662335, 0.4600803, 
    0.4463563, 0.448828, 0.444643, 0.4406536, 0.4339711, 0.4350697, 
    0.4321307, 0.444754, 0.4363557, 0.4502369, 0.4464315, 0.4767978, 
    0.4884745, 0.4934475, 0.4978091, 0.5084394, 0.5010949, 0.5039884, 
    0.4971091, 0.4927442, 0.4949025, 0.4816062, 0.4867688, 0.459716, 
    0.4713602, 0.4411185, 0.4483205, 0.4393959, 0.4439456, 0.4361556, 
    0.4431653, 0.4310382, 0.4284066, 0.4302045, 0.4233084, 0.4435544, 
    0.4357551, 0.4949628, 0.4946107, 0.4929711, 0.5001839, 0.5006257, 
    0.50725, 0.5013555, 0.4988479, 0.4924917, 0.4887369, 0.4851718, 
    0.4773476, 0.4686809, 0.4565389, 0.4478529, 0.4420488, 0.4456062, 
    0.4424651, 0.4459767, 0.4476246, 0.429392, 0.4396103, 0.4242988, 
    0.4251431, 0.4320607, 0.4250479, 0.4943635, 0.49639, 0.5034337, 
    0.4979202, 0.5079721, 0.5023417, 0.4991079, 0.48666, 0.4839323, 
    0.4814039, 0.4764175, 0.4700781, 0.4589046, 0.4492236, 0.4404218, 
    0.4410656, 0.4408389, 0.4388767, 0.44374, 0.4380794, 0.4371306, 
    0.4396119, 0.4252562, 0.4293471, 0.425161, 0.4278236, 0.4957313, 
    0.4923229, 0.4941641, 0.4907024, 0.4931406, 0.4823119, 0.4790725, 
    0.4640094, 0.4702035, 0.4603534, 0.4692016, 0.4676314, 0.4600312, 
    0.4687229, 0.4497557, 0.462598, 0.4388005, 0.4515631, 0.4380032, 
    0.4404598, 0.4363943, 0.4327594, 0.4281965, 0.4198042, 0.4217443, 
    0.4147483, 0.4872485, 0.4828394, 0.483228, 0.4786205, 0.4752175, 
    0.4679033, 0.4561337, 0.4605534, 0.4524463, 0.4508218, 0.4631412, 
    0.4555693, 0.4798926, 0.4759407, 0.4782935, 0.4869, 0.4595333, 0.4735232, 
    0.4477095, 0.4552696, 0.4332772, 0.4441864, 0.4228131, 0.4137458, 
    0.4052577, 0.3953897, 0.4804364, 0.4834293, 0.4780733, 0.470726, 
    0.463881, 0.4548076, 0.4538816, 0.4521859, 0.4478003, 0.4441191, 
    0.4516494, 0.4431973, 0.4750236, 0.4583186, 0.4845609, 0.4766191, 
    0.4711619, 0.473528, 0.4610592, 0.4581173, 0.4461989, 0.4523529, 
    0.4159789, 0.4319915, 0.3879201, 0.400119, 0.4844754, 0.4804471, 
    0.4665156, 0.4731113, 0.4542035, 0.4495589, 0.4457906, 0.4409818, 
    0.4404638, 0.4376203, 0.4422817, 0.4378045, 0.4547884, 0.4471829, 
    0.4681112, 0.4630009, 0.4653509, 0.4679304, 0.4599772, 0.4515305, 
    0.4513514, 0.4486493, 0.4410502, 0.454127, 0.4139202, 0.4386565, 
    0.4760605, 0.4683741, 0.4672721, 0.4702652, 0.4500241, 0.4573391, 
    0.4376898, 0.4429836, 0.4343169, 0.438619, 0.4392526, 0.4447927, 
    0.4482487, 0.457003, 0.4641495, 0.469831, 0.4685089, 0.4622717, 0.451015, 
    0.4404163, 0.4427336, 0.4349743, 0.4555732, 0.4469121, 0.4502555, 
    0.4415483, 0.4606707, 0.4443735, 0.4648535, 0.4630513, 0.4574846, 
    0.4463251, 0.4438651, 0.4412394, 0.4428595, 0.4507301, 0.4520227, 
    0.45762, 0.4591671, 0.4634436, 0.466989, 0.4637493, 0.4603511, 0.4507273, 
    0.4420876, 0.4327075, 0.4304189, 0.4195243, 0.4283868, 0.4137831, 
    0.4261895, 0.4047692, 0.4434343, 0.4265578, 0.4572319, 0.4539074, 
    0.4479047, 0.4342003, 0.4415892, 0.4329511, 0.4520734, 0.4620562, 
    0.4646469, 0.469485, 0.4645364, 0.4649386, 0.4602112, 0.4617295, 
    0.4504084, 0.4564831, 0.4392683, 0.4330194, 0.4154798, 0.4048102, 
    0.3940214, 0.3892816, 0.387842, 0.3872406,
  0.0499117, 0.0480224, 0.04838631, 0.04688734, 0.04771541, 0.04673891, 
    0.04952522, 0.04794822, 0.04895146, 0.04973995, 0.04405922, 0.04682115, 
    0.04129904, 0.04298105, 0.03883455, 0.04155796, 0.03829936, 0.03891169, 
    0.03708753, 0.0376045, 0.03533095, 0.03685046, 0.03418794, 0.03569023, 
    0.03545243, 0.03690125, 0.0462573, 0.04439745, 0.04636891, 0.04610047, 
    0.04622085, 0.04769816, 0.04845314, 0.05005803, 0.04976438, 0.04858683, 
    0.04598008, 0.04685535, 0.04466895, 0.04471763, 0.04235641, 0.04341131, 
    0.03956003, 0.04063216, 0.03758284, 0.03833568, 0.03761796, 0.03783471, 
    0.03761514, 0.03872309, 0.03824591, 0.03923, 0.0432125, 0.04201725, 
    0.04564302, 0.04791143, 0.04945538, 0.05056866, 0.05041037, 0.05010941, 
    0.04857998, 0.04716805, 0.04610883, 0.04540839, 0.04472463, 0.04269297, 
    0.04164146, 0.03934532, 0.03975386, 0.03906342, 0.0384111, 0.03733116, 
    0.0375076, 0.03703652, 0.03908166, 0.0377147, 0.03998772, 0.03935772, 
    0.04453921, 0.04661827, 0.04751887, 0.04831621, 0.05028886, 0.0489215, 
    0.04945782, 0.04818777, 0.04739096, 0.04778408, 0.04538933, 0.04631146, 
    0.04157964, 0.04357954, 0.03848683, 0.0396698, 0.03820663, 0.03894898, 
    0.03768243, 0.03882113, 0.03686221, 0.03644404, 0.03672946, 0.03564094, 
    0.03888487, 0.03761791, 0.04779509, 0.04773083, 0.04743221, 0.04875328, 
    0.04883484, 0.05006607, 0.04896968, 0.04850715, 0.04734507, 0.04666556, 
    0.04602516, 0.04463598, 0.04311502, 0.04104247, 0.03959243, 0.03863858, 
    0.03922179, 0.0387066, 0.03928277, 0.03955469, 0.03660033, 0.03824144, 
    0.03579622, 0.03592888, 0.03702534, 0.03591391, 0.04768575, 0.04805602, 
    0.04935477, 0.04833662, 0.05020126, 0.04915224, 0.048555, 0.04629194, 
    0.0458036, 0.04535339, 0.04447231, 0.04335693, 0.0414421, 0.03981946, 
    0.03837338, 0.03847821, 0.03844128, 0.03812239, 0.03891527, 0.03799321, 
    0.03783976, 0.03824171, 0.03594666, 0.0365932, 0.0359317, 0.03635174, 
    0.04793549, 0.04731441, 0.0476494, 0.04702061, 0.04746302, 0.0455148, 
    0.04494032, 0.04231133, 0.04337868, 0.04168785, 0.04320509, 0.04293377, 
    0.04163314, 0.04312228, 0.03990776, 0.04207005, 0.03811003, 0.0402085, 
    0.03798086, 0.03837956, 0.03772091, 0.03713704, 0.03641075, 0.03509426, 
    0.0353964, 0.03431321, 0.04639763, 0.04560871, 0.04567796, 0.04486046, 
    0.04426163, 0.0429807, 0.04097422, 0.04172183, 0.04035588, 0.04008501, 
    0.04216282, 0.04087926, 0.0450854, 0.04438855, 0.04480274, 0.04633503, 
    0.04154865, 0.04396506, 0.03956872, 0.04082888, 0.03721992, 0.03898847, 
    0.0355634, 0.03415943, 0.03287147, 0.03140602, 0.04518174, 0.04571385, 
    0.04476388, 0.04346936, 0.04228934, 0.04075129, 0.04059597, 0.04031239, 
    0.03958374, 0.03897744, 0.04022288, 0.03882638, 0.04422765, 0.04134292, 
    0.04591589, 0.04450776, 0.04354507, 0.04396591, 0.04180784, 0.04130888, 
    0.03931938, 0.04034027, 0.03450249, 0.03701429, 0.03031948, 0.03210407, 
    0.04590062, 0.04518362, 0.04274151, 0.04389313, 0.04064993, 0.03987509, 
    0.03925214, 0.03846455, 0.0383802, 0.03791892, 0.03867663, 0.03794872, 
    0.04074805, 0.03948171, 0.04301659, 0.04213886, 0.04254131, 0.04298538, 
    0.04162396, 0.04020305, 0.04017321, 0.03972425, 0.0384757, 0.04063711, 
    0.03418616, 0.03808669, 0.04440958, 0.043062, 0.04287182, 0.04338938, 
    0.03995235, 0.04117743, 0.03793015, 0.03879139, 0.03738666, 0.03808061, 
    0.03818337, 0.03908802, 0.03965791, 0.04112072, 0.04233531, 0.0433141, 
    0.0430853, 0.04201438, 0.04011717, 0.03837248, 0.03875049, 0.03749227, 
    0.04087992, 0.039437, 0.03999081, 0.03855691, 0.04174177, 0.03901919, 
    0.04245596, 0.04214747, 0.04120198, 0.03934018, 0.03893578, 0.03850654, 
    0.03877109, 0.04006975, 0.04028515, 0.04122484, 0.04148658, 0.04221452, 
    0.04282303, 0.0422668, 0.04168745, 0.04006927, 0.03864493, 0.03712874, 
    0.03676358, 0.0350508, 0.03644091, 0.03416515, 0.03609364, 0.03279811, 
    0.03886519, 0.03615173, 0.04115933, 0.0406003, 0.03960101, 0.03736793, 
    0.03856358, 0.03716771, 0.04029361, 0.04197763, 0.04242054, 0.04325416, 
    0.0424016, 0.04247056, 0.04166369, 0.04192195, 0.04001623, 0.04103307, 
    0.03818591, 0.03717865, 0.03442566, 0.03280426, 0.03120552, 0.03051606, 
    0.03030822, 0.03022159,
  0.001340993, 0.001263546, 0.00127834, 0.00121778, 0.001251111, 0.001211839, 
    0.001325022, 0.001260537, 0.001301433, 0.001333887, 0.001106295, 
    0.00121513, 0.001001077, 0.001064767, 0.0009102243, 0.001010794, 
    0.0008908893, 0.0009130226, 0.0008476403, 0.000866, 0.0007862778, 
    0.0008392662, 0.0007477449, 0.000798699, 0.0007904702, 0.000841058, 
    0.001192628, 0.001119435, 0.00119707, 0.001186395, 0.001191178, 
    0.001250413, 0.001281064, 0.001347057, 0.001334897, 0.001286518, 
    0.001181617, 0.001216499, 0.00113002, 0.001131922, 0.001040958, 
    0.001081274, 0.0009366602, 0.000976201, 0.0008652278, 0.0008921969, 
    0.0008664798, 0.0008742191, 0.0008663793, 0.0009061857, 0.000888966, 
    0.0009246017, 0.001073636, 0.001028108, 0.001168278, 0.001259046, 
    0.001322143, 0.001368291, 0.001361696, 0.001349188, 0.001286238, 
    0.001229045, 0.001186726, 0.001159023, 0.001132195, 0.001053764, 
    0.001013934, 0.0009288092, 0.0009437672, 0.0009185361, 0.0008949142, 
    0.0008562757, 0.0008625484, 0.0008458361, 0.0009191993, 0.000869931, 
    0.0009523662, 0.0009292621, 0.001124957, 0.001207016, 0.001243172, 
    0.001275486, 0.001356641, 0.001300205, 0.001322243, 0.001270261, 
    0.001238015, 0.001253889, 0.001158272, 0.001194783, 0.001011609, 
    0.001087752, 0.0008976457, 0.0009406829, 0.0008875538, 0.0009143766, 
    0.0008687793, 0.0009097377, 0.0008396804, 0.0008249772, 0.0008350033, 
    0.0007969909, 0.0009120492, 0.0008664779, 0.001254334, 0.001251735, 
    0.001239677, 0.001293319, 0.001296656, 0.00134739, 0.00130218, 
    0.001283266, 0.001236166, 0.001208906, 0.001183406, 0.001128733, 
    0.001069898, 0.0009914811, 0.0009378471, 0.0009031278, 0.0009243024, 
    0.0009055889, 0.0009265264, 0.0009364645, 0.0008304621, 0.0008888054, 
    0.0008023762, 0.0008069867, 0.0008454408, 0.0008064663, 0.001249912, 
    0.00126491, 0.001317999, 0.001276317, 0.001353002, 0.001309671, 
    0.001285219, 0.001194006, 0.001174627, 0.001156857, 0.00112235, 
    0.001079183, 0.001006442, 0.0009461765, 0.000893555, 0.0008973347, 
    0.0008960025, 0.0008845274, 0.0009131525, 0.0008798933, 0.0008743996, 
    0.000888815, 0.0008076056, 0.0008302115, 0.0008070849, 0.0008217437, 
    0.001260021, 0.001234932, 0.001248443, 0.001223124, 0.00124092, 
    0.001163217, 0.001140635, 0.001039247, 0.001080019, 0.00101568, 
    0.001073351, 0.001062959, 0.001013621, 0.001070176, 0.0009494232, 
    0.001030105, 0.0008840836, 0.0009605091, 0.0008794507, 0.0008937777, 
    0.0008701528, 0.0008493926, 0.0008238106, 0.0007781319, 0.0007885356, 
    0.0007514586, 0.001198215, 0.001166923, 0.001169658, 0.001137508, 
    0.001114152, 0.001064754, 0.0009889338, 0.00101696, 0.0009659579, 
    0.0009559519, 0.001033617, 0.0009853934, 0.001146323, 0.001119088, 
    0.001135249, 0.001195721, 0.001010444, 0.001102647, 0.0009369785, 
    0.0009835167, 0.0008523291, 0.0009158113, 0.0007943065, 0.0007467764, 
    0.0007034835, 0.0006553396, 0.001150106, 0.001171077, 0.001133729, 
    0.001083508, 0.001038412, 0.000980629, 0.0009748572, 0.0009643492, 
    0.0009375284, 0.0009154102, 0.0009610403, 0.0009099278, 0.001112832, 
    0.001002722, 0.001179073, 0.001123731, 0.001086424, 0.00110268, 
    0.001020201, 0.001001446, 0.0009278622, 0.0009653805, 0.0007578932, 
    0.0008450503, 0.0006204266, 0.000678123, 0.001178468, 0.00115018, 
    0.001055615, 0.001099863, 0.000976861, 0.0009482217, 0.0009254091, 
    0.0008968419, 0.0008938006, 0.0008772322, 0.000904504, 0.0008782992, 
    0.0009805086, 0.0009337938, 0.001066127, 0.001032709, 0.001047986, 
    0.001064933, 0.001013275, 0.0009603079, 0.000959206, 0.0009426803, 
    0.000897244, 0.0009763847, 0.0007476844, 0.0008832458, 0.001119907, 
    0.001067866, 0.00106059, 0.001080431, 0.0009510641, 0.0009965249, 
    0.0008776342, 0.0009086597, 0.0008582468, 0.0008830276, 0.0008867179, 
    0.0009194309, 0.0009402467, 0.0009944044, 0.001040157, 0.001077537, 
    0.001068759, 0.001027999, 0.000957138, 0.0008935226, 0.0009071779, 
    0.0008620027, 0.0009854181, 0.0009321587, 0.00095248, 0.000900176, 
    0.001017711, 0.0009169276, 0.00104474, 0.001033035, 0.0009974435, 
    0.0009286214, 0.0009138971, 0.0008983572, 0.000907924, 0.0009553891, 
    0.0009633416, 0.0009982992, 0.001008112, 0.001035576, 0.001058726, 
    0.001037558, 0.001015665, 0.0009553715, 0.0009033574, 0.0008490989, 
    0.0008362046, 0.000776639, 0.0008248673, 0.0007469706, 0.0008127258, 
    0.0007010449, 0.0009113352, 0.0008147525, 0.0009958482, 0.0009750179, 
    0.000938161, 0.0008575816, 0.0009004169, 0.0008504788, 0.0009636546, 
    0.00102661, 0.001043394, 0.001075235, 0.001042674, 0.001045295, 
    0.001014771, 0.001024507, 0.0009534166, 0.0009911302, 0.000886809, 
    0.0008508664, 0.000755279, 0.0007012494, 0.0006488466, 0.0006266933, 
    0.0006200684, 0.0006173147,
  8.818055e-06, 8.041776e-06, 8.18829e-06, 7.59401e-06, 7.919295e-06, 
    7.536489e-06, 8.656109e-06, 8.012087e-06, 8.418673e-06, 8.745884e-06, 
    6.539152e-06, 7.568332e-06, 5.593384e-06, 6.159866e-06, 4.818944e-06, 
    5.678582e-06, 4.659502e-06, 4.84218e-06, 4.310015e-06, 4.457151e-06, 
    3.831833e-06, 4.243515e-06, 3.213127e-06, 3.926902e-06, 3.86382e-06, 
    4.257711e-06, 7.351498e-06, 6.660739e-06, 7.394144e-06, 7.291803e-06, 
    7.337599e-06, 7.912439e-06, 8.215355e-06, 8.879793e-06, 8.756131e-06, 
    8.269634e-06, 7.246156e-06, 7.581594e-06, 6.759237e-06, 6.776981e-06, 
    5.945907e-06, 6.309713e-06, 5.040052e-06, 5.377301e-06, 4.450927e-06, 
    4.670224e-06, 4.461021e-06, 4.523608e-06, 4.46021e-06, 4.78548e-06, 
    4.643749e-06, 4.938755e-06, 6.240222e-06, 5.831507e-06, 7.119199e-06, 
    7.997382e-06, 8.627016e-06, 9.097052e-06, 9.029402e-06, 8.901525e-06, 
    8.266851e-06, 7.703446e-06, 7.294975e-06, 7.03155e-06, 6.779535e-06, 
    6.060664e-06, 5.706213e-06, 4.974016e-06, 5.100097e-06, 4.88808e-06, 
    4.692533e-06, 4.378992e-06, 4.429351e-06, 4.295655e-06, 4.893611e-06, 
    4.488891e-06, 5.173085e-06, 4.977817e-06, 6.712065e-06, 7.489914e-06, 
    7.841413e-06, 8.159954e-06, 8.977654e-06, 8.406373e-06, 8.628032e-06, 
    8.108176e-06, 7.790956e-06, 7.946601e-06, 7.024456e-06, 7.372177e-06, 
    5.685749e-06, 6.368848e-06, 4.714997e-06, 5.074009e-06, 4.632194e-06, 
    4.853438e-06, 4.479583e-06, 4.814908e-06, 4.246795e-06, 4.130939e-06, 
    4.209811e-06, 3.913775e-06, 4.834093e-06, 4.461006e-06, 7.950985e-06, 
    7.925421e-06, 7.807209e-06, 8.33749e-06, 8.370848e-06, 8.883189e-06, 
    8.426158e-06, 8.237259e-06, 7.772896e-06, 7.508153e-06, 7.26323e-06, 
    6.747232e-06, 6.20631e-06, 5.509677e-06, 5.050063e-06, 4.760199e-06, 
    4.93625e-06, 4.780543e-06, 4.954874e-06, 5.038402e-06, 4.174018e-06, 
    4.642435e-06, 3.955217e-06, 3.990828e-06, 4.292512e-06, 3.986802e-06, 
    7.907513e-06, 8.055252e-06, 8.585201e-06, 8.168199e-06, 8.940449e-06, 
    8.501353e-06, 8.256694e-06, 7.364718e-06, 7.17953e-06, 7.011093e-06, 
    6.687818e-06, 6.290662e-06, 5.640369e-06, 5.12051e-06, 4.681369e-06, 
    4.712437e-06, 4.701479e-06, 4.607468e-06, 4.843259e-06, 4.569699e-06, 
    4.525072e-06, 4.642513e-06, 3.995618e-06, 4.172045e-06, 3.991588e-06, 
    4.105621e-06, 8.006996e-06, 7.760844e-06, 7.893091e-06, 7.64586e-06, 
    7.819363e-06, 7.071226e-06, 6.858482e-06, 5.930629e-06, 6.298279e-06, 
    5.721598e-06, 6.237641e-06, 6.143523e-06, 5.703455e-06, 6.208832e-06, 
    5.148064e-06, 5.849235e-06, 4.603846e-06, 5.242539e-06, 4.566098e-06, 
    4.683197e-06, 4.490685e-06, 4.323979e-06, 4.121798e-06, 3.769974e-06, 
    3.849048e-06, 3.570167e-06, 7.405143e-06, 7.106345e-06, 7.132302e-06, 
    6.829195e-06, 6.611765e-06, 6.159745e-06, 5.487531e-06, 5.732881e-06, 
    5.289197e-06, 5.203629e-06, 5.880457e-06, 5.456803e-06, 6.911871e-06, 
    6.657525e-06, 6.808067e-06, 7.381186e-06, 5.675506e-06, 6.505526e-06, 
    5.042736e-06, 5.440539e-06, 4.347418e-06, 4.865376e-06, 3.893181e-06, 
    3.207773e-06, 2.969702e-06, 2.707985e-06, 6.94745e-06, 7.145773e-06, 
    6.793863e-06, 6.330082e-06, 5.923184e-06, 5.415546e-06, 5.365715e-06, 
    5.275407e-06, 5.047373e-06, 4.862038e-06, 5.247082e-06, 4.816485e-06, 
    6.599545e-06, 5.607772e-06, 7.221885e-06, 6.700661e-06, 6.356707e-06, 
    6.505828e-06, 5.761497e-06, 5.59661e-06, 4.966073e-06, 5.284247e-06, 
    3.617979e-06, 4.289406e-06, 2.520337e-06, 2.831426e-06, 7.216117e-06, 
    6.948147e-06, 6.077317e-06, 6.479902e-06, 5.382996e-06, 5.137861e-06, 
    4.945515e-06, 4.708382e-06, 4.683386e-06, 4.548063e-06, 4.771571e-06, 
    4.556733e-06, 5.414505e-06, 5.015906e-06, 6.17217e-06, 5.872383e-06, 
    6.008798e-06, 6.161363e-06, 5.700417e-06, 5.24082e-06, 5.231404e-06, 
    5.090898e-06, 4.711691e-06, 5.378886e-06, 3.212793e-06, 4.597011e-06, 
    6.665122e-06, 6.187905e-06, 6.122147e-06, 6.302024e-06, 5.162009e-06, 
    5.553618e-06, 4.551328e-06, 4.80597e-06, 4.394793e-06, 4.595231e-06, 
    4.62536e-06, 4.895544e-06, 5.070322e-06, 5.53513e-06, 5.938753e-06, 
    6.275681e-06, 6.195987e-06, 5.830545e-06, 5.213746e-06, 4.681103e-06, 
    4.793694e-06, 4.424961e-06, 5.457017e-06, 5.002151e-06, 5.174054e-06, 
    4.73584e-06, 5.739508e-06, 4.874672e-06, 5.97972e-06, 5.875281e-06, 
    5.561633e-06, 4.972441e-06, 4.84945e-06, 4.720854e-06, 4.799873e-06, 
    5.19883e-06, 5.266776e-06, 5.569105e-06, 5.655021e-06, 5.897896e-06, 
    6.105339e-06, 5.91556e-06, 5.721465e-06, 5.19868e-06, 4.762096e-06, 
    4.321637e-06, 4.219299e-06, 3.758679e-06, 4.130077e-06, 3.208847e-06, 
    4.035325e-06, 2.956367e-06, 4.828164e-06, 4.051084e-06, 5.547716e-06, 
    5.367099e-06, 5.052711e-06, 4.389459e-06, 4.737827e-06, 4.332644e-06, 
    5.269457e-06, 5.818226e-06, 5.967677e-06, 6.254751e-06, 5.961242e-06, 
    5.984689e-06, 5.713584e-06, 5.799587e-06, 5.182026e-06, 5.506624e-06, 
    4.626105e-06, 4.335737e-06, 3.598524e-06, 2.957485e-06, 2.672947e-06, 
    2.55388e-06, 2.518421e-06, 2.503703e-06,
  8.089846e-09, 6.902192e-09, 7.123347e-09, 6.235646e-09, 6.718446e-09, 
    6.151083e-09, 7.83893e-09, 6.857557e-09, 7.473989e-09, 7.977829e-09, 
    4.727549e-09, 6.197864e-09, 3.464642e-09, 4.209749e-09, 2.510204e-09, 
    3.574376e-09, 2.324393e-09, 2.537613e-09, 1.931808e-09, 2.094521e-09, 
    1.431628e-09, 1.859556e-09, 1.147179e-09, 1.527335e-09, 1.46361e-09, 
    1.874911e-09, 5.880839e-09, 4.896475e-09, 5.942903e-09, 5.794204e-09, 
    5.860642e-09, 6.708191e-09, 7.164357e-09, 8.185918e-09, 7.993714e-09, 
    7.246754e-09, 5.728149e-09, 6.217372e-09, 5.034317e-09, 5.059241e-09, 
    3.924141e-09, 4.412616e-09, 2.774274e-09, 3.190307e-09, 2.087561e-09, 
    2.336762e-09, 2.098852e-09, 2.169259e-09, 2.097945e-09, 2.470876e-09, 
    2.306255e-09, 2.652401e-09, 4.318255e-09, 3.77347e-09, 5.545318e-09, 
    6.835472e-09, 7.794024e-09, 8.525777e-09, 8.419659e-09, 8.219788e-09, 
    7.242525e-09, 6.397213e-09, 5.798801e-09, 5.419872e-09, 5.062831e-09, 
    4.076722e-09, 3.610148e-09, 2.694656e-09, 2.84721e-09, 2.591995e-09, 
    2.362557e-09, 2.007607e-09, 2.063484e-09, 1.916136e-09, 2.59857e-09, 
    2.130121e-09, 2.936544e-09, 2.699222e-09, 4.968193e-09, 6.082794e-09, 
    6.602155e-09, 7.080462e-09, 8.338662e-09, 7.45518e-09, 7.795592e-09, 
    7.00224e-09, 6.527045e-09, 6.759319e-09, 5.409746e-09, 5.910916e-09, 
    3.583646e-09, 4.493295e-09, 2.388611e-09, 2.815458e-09, 2.292975e-09, 
    2.550922e-09, 2.119664e-09, 2.505452e-09, 1.863101e-09, 1.739148e-09, 
    1.823253e-09, 1.514004e-09, 2.528064e-09, 2.098835e-09, 6.765887e-09, 
    6.72761e-09, 6.551219e-09, 7.350032e-09, 7.400915e-09, 8.191209e-09, 
    7.485439e-09, 7.197585e-09, 6.500205e-09, 6.109517e-09, 5.752837e-09, 
    5.017469e-09, 4.272382e-09, 3.357681e-09, 2.786399e-09, 2.44128e-09, 
    2.649406e-09, 2.465089e-09, 2.671695e-09, 2.772278e-09, 1.784936e-09, 
    2.304743e-09, 1.556215e-09, 1.592777e-09, 1.912711e-09, 1.58863e-09, 
    6.700825e-09, 6.922472e-09, 7.729573e-09, 7.092935e-09, 8.280526e-09, 
    7.600665e-09, 7.227093e-09, 5.900063e-09, 5.632037e-09, 5.390685e-09, 
    4.934283e-09, 4.386699e-09, 3.52505e-09, 2.87212e-09, 2.349638e-09, 
    2.385639e-09, 2.372923e-09, 2.264631e-09, 2.538888e-09, 2.221532e-09, 
    2.170913e-09, 2.304833e-09, 1.597715e-09, 1.782832e-09, 1.59356e-09, 
    1.712408e-09, 6.84991e-09, 6.482307e-09, 6.679271e-09, 6.312086e-09, 
    6.569308e-09, 5.476578e-09, 5.174084e-09, 3.903935e-09, 4.397056e-09, 
    3.630105e-09, 4.314758e-09, 4.187764e-09, 3.606574e-09, 4.275789e-09, 
    2.905836e-09, 3.796723e-09, 2.260488e-09, 3.022227e-09, 2.217435e-09, 
    2.351753e-09, 2.132139e-09, 1.947084e-09, 1.729479e-09, 1.370426e-09, 
    1.448812e-09, 1.17881e-09, 5.958933e-09, 5.526882e-09, 5.564127e-09, 
    5.132749e-09, 4.828268e-09, 4.209587e-09, 3.329527e-09, 3.644759e-09, 
    3.080151e-09, 2.974144e-09, 3.837761e-09, 3.290564e-09, 5.249631e-09, 
    4.891992e-09, 5.102976e-09, 5.924029e-09, 3.570399e-09, 4.681077e-09, 
    2.777524e-09, 3.269988e-09, 1.972803e-09, 2.565056e-09, 1.493163e-09, 
    1.140588e-09, 8.646354e-10, 6.018309e-10, 5.300113e-09, 5.583479e-09, 
    5.082982e-09, 4.440368e-09, 3.894098e-09, 3.238436e-09, 3.175763e-09, 
    3.063001e-09, 2.783141e-09, 2.561102e-09, 3.027854e-09, 2.507308e-09, 
    4.811283e-09, 3.483112e-09, 5.693094e-09, 4.952237e-09, 4.476704e-09, 
    4.681494e-09, 3.681989e-09, 3.468781e-09, 2.685121e-09, 3.073991e-09, 
    1.223791e-09, 1.909329e-09, 4.413377e-10, 7.202956e-10, 5.684771e-09, 
    5.301103e-09, 4.098981e-09, 4.645735e-09, 3.197462e-09, 2.893338e-09, 
    2.660487e-09, 2.380931e-09, 2.351971e-09, 2.196949e-09, 2.454581e-09, 
    2.206791e-09, 3.237124e-09, 2.74509e-09, 4.226321e-09, 3.827139e-09, 
    4.007585e-09, 4.211766e-09, 3.602637e-09, 3.020098e-09, 3.008445e-09, 
    2.836003e-09, 2.384771e-09, 3.192298e-09, 1.146766e-09, 2.252675e-09, 
    4.90259e-09, 4.247535e-09, 4.159048e-09, 4.402152e-09, 2.92294e-09, 
    3.413723e-09, 2.200654e-09, 2.494936e-09, 2.025092e-09, 2.250642e-09, 
    2.285131e-09, 2.600868e-09, 2.810979e-09, 3.390114e-09, 3.914677e-09, 
    4.366344e-09, 4.258442e-09, 3.772209e-09, 2.986627e-09, 2.349331e-09, 
    2.480514e-09, 2.058595e-09, 3.290834e-09, 2.728502e-09, 2.937734e-09, 
    2.412858e-09, 3.653372e-09, 2.576077e-09, 3.968951e-09, 3.83095e-09, 
    3.423971e-09, 2.692764e-09, 2.546205e-09, 2.395418e-09, 2.487771e-09, 
    2.968229e-09, 3.05228e-09, 3.43353e-09, 3.543943e-09, 3.860731e-09, 
    4.136502e-09, 3.884031e-09, 3.629933e-09, 2.968044e-09, 2.443497e-09, 
    1.944519e-09, 1.833451e-09, 1.359344e-09, 1.738236e-09, 1.141908e-09, 
    1.638831e-09, 8.501922e-10, 2.52107e-09, 1.655239e-09, 3.406181e-09, 
    3.1775e-09, 2.789609e-09, 2.019184e-09, 2.415172e-09, 1.956579e-09, 
    3.055609e-09, 3.756074e-09, 3.952977e-09, 4.337942e-09, 3.944448e-09, 
    3.975547e-09, 3.619706e-09, 3.731692e-09, 2.947537e-09, 3.353797e-09, 
    2.285986e-09, 1.959973e-09, 1.205421e-09, 8.51399e-10, 5.700418e-10, 
    4.682473e-10, 4.398248e-10, 4.282862e-10,
  4.32761e-13, 4.280988e-13, 4.289675e-13, 4.254785e-13, 4.273767e-13, 
    4.251458e-13, 4.317767e-13, 4.279234e-13, 4.303444e-13, 4.323216e-13, 
    4.195388e-13, 4.253299e-13, 4.14551e-13, 4.174955e-13, 4.107719e-13, 
    4.149849e-13, 4.100349e-13, 4.108805e-13, 4.084764e-13, 4.091226e-13, 
    4.064874e-13, 4.081893e-13, 4.053598e-13, 4.068683e-13, 4.066147e-13, 
    4.082503e-13, 4.240825e-13, 4.20205e-13, 4.243268e-13, 4.237415e-13, 
    4.24003e-13, 4.273364e-13, 4.291286e-13, 4.331378e-13, 4.323839e-13, 
    4.294522e-13, 4.234815e-13, 4.254066e-13, 4.207484e-13, 4.208466e-13, 
    4.163674e-13, 4.182963e-13, 4.118184e-13, 4.134656e-13, 4.09095e-13, 
    4.10084e-13, 4.091398e-13, 4.094193e-13, 4.091362e-13, 4.106159e-13, 
    4.09963e-13, 4.113355e-13, 4.179238e-13, 4.15772e-13, 4.227617e-13, 
    4.278366e-13, 4.316005e-13, 4.344703e-13, 4.340543e-13, 4.332706e-13, 
    4.294356e-13, 4.261139e-13, 4.237596e-13, 4.222676e-13, 4.208608e-13, 
    4.169701e-13, 4.151264e-13, 4.11503e-13, 4.121074e-13, 4.110961e-13, 
    4.101863e-13, 4.087775e-13, 4.089994e-13, 4.084141e-13, 4.111222e-13, 
    4.092639e-13, 4.124612e-13, 4.115211e-13, 4.204877e-13, 4.248772e-13, 
    4.269196e-13, 4.287991e-13, 4.337367e-13, 4.302706e-13, 4.316066e-13, 
    4.284918e-13, 4.266244e-13, 4.275373e-13, 4.222277e-13, 4.242009e-13, 
    4.150216e-13, 4.186147e-13, 4.102897e-13, 4.119816e-13, 4.099103e-13, 
    4.109333e-13, 4.092224e-13, 4.10753e-13, 4.082034e-13, 4.077107e-13, 
    4.08045e-13, 4.068152e-13, 4.108427e-13, 4.091397e-13, 4.275631e-13, 
    4.274127e-13, 4.267194e-13, 4.298578e-13, 4.300575e-13, 4.331585e-13, 
    4.303893e-13, 4.292591e-13, 4.265188e-13, 4.249823e-13, 4.235787e-13, 
    4.20682e-13, 4.177427e-13, 4.141279e-13, 4.118665e-13, 4.104985e-13, 
    4.113237e-13, 4.10593e-13, 4.11412e-13, 4.118105e-13, 4.078927e-13, 
    4.09957e-13, 4.069832e-13, 4.071286e-13, 4.084005e-13, 4.071121e-13, 
    4.273075e-13, 4.281784e-13, 4.313476e-13, 4.288481e-13, 4.335088e-13, 
    4.308416e-13, 4.29375e-13, 4.241582e-13, 4.231031e-13, 4.221526e-13, 
    4.20354e-13, 4.18194e-13, 4.147899e-13, 4.12206e-13, 4.101351e-13, 
    4.102779e-13, 4.102274e-13, 4.097978e-13, 4.108856e-13, 4.096268e-13, 
    4.094259e-13, 4.099573e-13, 4.071483e-13, 4.078844e-13, 4.071318e-13, 
    4.076044e-13, 4.278933e-13, 4.264485e-13, 4.272227e-13, 4.257791e-13, 
    4.267905e-13, 4.224909e-13, 4.212992e-13, 4.162876e-13, 4.182349e-13, 
    4.152053e-13, 4.1791e-13, 4.174086e-13, 4.151123e-13, 4.177562e-13, 
    4.123395e-13, 4.158639e-13, 4.097814e-13, 4.128004e-13, 4.096105e-13, 
    4.101435e-13, 4.09272e-13, 4.085371e-13, 4.076723e-13, 4.062438e-13, 
    4.065558e-13, 4.054805e-13, 4.243899e-13, 4.22689e-13, 4.228357e-13, 
    4.211363e-13, 4.19936e-13, 4.174948e-13, 4.140165e-13, 4.152632e-13, 
    4.130297e-13, 4.126101e-13, 4.160261e-13, 4.138623e-13, 4.215969e-13, 
    4.201873e-13, 4.21019e-13, 4.242525e-13, 4.149692e-13, 4.193555e-13, 
    4.118313e-13, 4.137809e-13, 4.086392e-13, 4.109893e-13, 4.067323e-13, 
    4.053335e-13, 4.042316e-13, 4.031807e-13, 4.217958e-13, 4.229119e-13, 
    4.209402e-13, 4.184058e-13, 4.162487e-13, 4.136561e-13, 4.134081e-13, 
    4.129618e-13, 4.118536e-13, 4.109736e-13, 4.128227e-13, 4.107604e-13, 
    4.198691e-13, 4.14624e-13, 4.233435e-13, 4.204248e-13, 4.185492e-13, 
    4.193571e-13, 4.154104e-13, 4.145674e-13, 4.114652e-13, 4.130053e-13, 
    4.056597e-13, 4.083871e-13, 4.025382e-13, 4.036546e-13, 4.233107e-13, 
    4.217997e-13, 4.17058e-13, 4.192161e-13, 4.13494e-13, 4.1229e-13, 
    4.113676e-13, 4.102592e-13, 4.101443e-13, 4.095292e-13, 4.105513e-13, 
    4.095683e-13, 4.136509e-13, 4.117028e-13, 4.175609e-13, 4.159841e-13, 
    4.166971e-13, 4.175034e-13, 4.150967e-13, 4.12792e-13, 4.127458e-13, 
    4.12063e-13, 4.102744e-13, 4.134735e-13, 4.053582e-13, 4.097504e-13, 
    4.202291e-13, 4.176447e-13, 4.172952e-13, 4.18255e-13, 4.124073e-13, 
    4.143496e-13, 4.095439e-13, 4.107113e-13, 4.088469e-13, 4.097423e-13, 
    4.098791e-13, 4.111313e-13, 4.119638e-13, 4.142562e-13, 4.1633e-13, 
    4.181137e-13, 4.176877e-13, 4.15767e-13, 4.126595e-13, 4.101338e-13, 
    4.106541e-13, 4.0898e-13, 4.138634e-13, 4.116371e-13, 4.124659e-13, 
    4.103858e-13, 4.152973e-13, 4.11033e-13, 4.165444e-13, 4.159992e-13, 
    4.143901e-13, 4.114955e-13, 4.109146e-13, 4.103167e-13, 4.106829e-13, 
    4.125866e-13, 4.129194e-13, 4.144279e-13, 4.148646e-13, 4.161168e-13, 
    4.172062e-13, 4.162089e-13, 4.152046e-13, 4.125859e-13, 4.105073e-13, 
    4.085269e-13, 4.080856e-13, 4.061996e-13, 4.077071e-13, 4.053388e-13, 
    4.073118e-13, 4.041739e-13, 4.108149e-13, 4.073771e-13, 4.143197e-13, 
    4.13415e-13, 4.118792e-13, 4.088234e-13, 4.10395e-13, 4.085748e-13, 
    4.129325e-13, 4.157033e-13, 4.164813e-13, 4.180015e-13, 4.164476e-13, 
    4.165705e-13, 4.151642e-13, 4.156069e-13, 4.125047e-13, 4.141125e-13, 
    4.098825e-13, 4.085883e-13, 4.055865e-13, 4.041787e-13, 4.030535e-13, 
    4.02646e-13, 4.025321e-13, 4.024859e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949654e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.94965e-07, 8.949651e-07, 8.949648e-07, 8.94965e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.94965e-07, 8.949651e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.94965e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.00961e-16, 6.025902e-16, 6.022737e-16, 6.035866e-16, 6.028587e-16, 
    6.03718e-16, 6.012916e-16, 6.026546e-16, 6.017848e-16, 6.01108e-16, 
    6.061305e-16, 6.036452e-16, 6.087103e-16, 6.07128e-16, 6.111002e-16, 
    6.084638e-16, 6.116314e-16, 6.110248e-16, 6.128513e-16, 6.123283e-16, 
    6.146609e-16, 6.130927e-16, 6.158697e-16, 6.142869e-16, 6.145344e-16, 
    6.130408e-16, 6.041462e-16, 6.058212e-16, 6.040468e-16, 6.042857e-16, 
    6.041786e-16, 6.028735e-16, 6.02215e-16, 6.008367e-16, 6.010871e-16, 
    6.020996e-16, 6.043933e-16, 6.036154e-16, 6.055761e-16, 6.055319e-16, 
    6.077115e-16, 6.067292e-16, 6.103881e-16, 6.093494e-16, 6.123502e-16, 
    6.115959e-16, 6.123147e-16, 6.120968e-16, 6.123175e-16, 6.112111e-16, 
    6.116852e-16, 6.107115e-16, 6.069131e-16, 6.080303e-16, 6.046955e-16, 
    6.02686e-16, 6.013514e-16, 6.004032e-16, 6.005373e-16, 6.007927e-16, 
    6.021055e-16, 6.033393e-16, 6.042788e-16, 6.049069e-16, 6.055255e-16, 
    6.073952e-16, 6.08385e-16, 6.105979e-16, 6.101992e-16, 6.108749e-16, 
    6.115209e-16, 6.126041e-16, 6.124259e-16, 6.129029e-16, 6.108575e-16, 
    6.12217e-16, 6.099722e-16, 6.105862e-16, 6.056918e-16, 6.038254e-16, 
    6.030298e-16, 6.023345e-16, 6.006403e-16, 6.018103e-16, 6.013492e-16, 
    6.024466e-16, 6.031432e-16, 6.027988e-16, 6.04924e-16, 6.040981e-16, 
    6.084437e-16, 6.065734e-16, 6.114456e-16, 6.10281e-16, 6.117246e-16, 
    6.109883e-16, 6.122495e-16, 6.111145e-16, 6.130805e-16, 6.13508e-16, 
    6.132159e-16, 6.143387e-16, 6.110514e-16, 6.123145e-16, 6.02789e-16, 
    6.028452e-16, 6.031071e-16, 6.019556e-16, 6.018852e-16, 6.008298e-16, 
    6.017691e-16, 6.021688e-16, 6.031837e-16, 6.037834e-16, 6.043533e-16, 
    6.056059e-16, 6.070032e-16, 6.089555e-16, 6.103565e-16, 6.112952e-16, 
    6.107198e-16, 6.112277e-16, 6.106598e-16, 6.103937e-16, 6.133477e-16, 
    6.116895e-16, 6.141772e-16, 6.140397e-16, 6.129142e-16, 6.140552e-16, 
    6.028846e-16, 6.025613e-16, 6.014378e-16, 6.023171e-16, 6.007149e-16, 
    6.016117e-16, 6.02127e-16, 6.041149e-16, 6.045518e-16, 6.049562e-16, 
    6.057551e-16, 6.067795e-16, 6.085746e-16, 6.10135e-16, 6.115585e-16, 
    6.114543e-16, 6.11491e-16, 6.118086e-16, 6.110214e-16, 6.119378e-16, 
    6.120914e-16, 6.116896e-16, 6.140213e-16, 6.133555e-16, 6.140368e-16, 
    6.136034e-16, 6.026665e-16, 6.032105e-16, 6.029166e-16, 6.034692e-16, 
    6.030797e-16, 6.048103e-16, 6.053288e-16, 6.077532e-16, 6.067592e-16, 
    6.083414e-16, 6.069201e-16, 6.07172e-16, 6.083922e-16, 6.069971e-16, 
    6.100489e-16, 6.079798e-16, 6.11821e-16, 6.097567e-16, 6.119502e-16, 
    6.115524e-16, 6.122112e-16, 6.128008e-16, 6.135427e-16, 6.149099e-16, 
    6.145934e-16, 6.157364e-16, 6.040214e-16, 6.047262e-16, 6.046645e-16, 
    6.054021e-16, 6.059473e-16, 6.071286e-16, 6.090211e-16, 6.083098e-16, 
    6.096157e-16, 6.098776e-16, 6.078937e-16, 6.091118e-16, 6.05198e-16, 
    6.058306e-16, 6.054543e-16, 6.040768e-16, 6.084733e-16, 6.062183e-16, 
    6.103796e-16, 6.091604e-16, 6.127167e-16, 6.109486e-16, 6.144192e-16, 
    6.158994e-16, 6.172929e-16, 6.189177e-16, 6.051111e-16, 6.046323e-16, 
    6.054899e-16, 6.066749e-16, 6.077745e-16, 6.092347e-16, 6.093842e-16, 
    6.096575e-16, 6.103653e-16, 6.109602e-16, 6.097435e-16, 6.111093e-16, 
    6.059766e-16, 6.08669e-16, 6.044509e-16, 6.057218e-16, 6.066052e-16, 
    6.062181e-16, 6.082286e-16, 6.087019e-16, 6.106235e-16, 6.096308e-16, 
    6.155339e-16, 6.129248e-16, 6.201549e-16, 6.181377e-16, 6.044649e-16, 
    6.051096e-16, 6.073509e-16, 6.06285e-16, 6.093324e-16, 6.100814e-16, 
    6.1069e-16, 6.114675e-16, 6.115516e-16, 6.120121e-16, 6.112574e-16, 
    6.119825e-16, 6.092379e-16, 6.104649e-16, 6.070954e-16, 6.07916e-16, 
    6.075387e-16, 6.071244e-16, 6.084026e-16, 6.097627e-16, 6.097923e-16, 
    6.102277e-16, 6.114539e-16, 6.093447e-16, 6.158692e-16, 6.118419e-16, 
    6.058124e-16, 6.070521e-16, 6.072298e-16, 6.067496e-16, 6.100063e-16, 
    6.08827e-16, 6.12001e-16, 6.111439e-16, 6.125482e-16, 6.118504e-16, 
    6.117477e-16, 6.108513e-16, 6.102926e-16, 6.08881e-16, 6.077313e-16, 
    6.068193e-16, 6.070315e-16, 6.080331e-16, 6.098459e-16, 6.11559e-16, 
    6.111838e-16, 6.124415e-16, 6.091116e-16, 6.105083e-16, 6.099686e-16, 
    6.11376e-16, 6.082908e-16, 6.109166e-16, 6.076186e-16, 6.079082e-16, 
    6.088036e-16, 6.106026e-16, 6.110012e-16, 6.114258e-16, 6.11164e-16, 
    6.09892e-16, 6.096838e-16, 6.08782e-16, 6.085326e-16, 6.078452e-16, 
    6.072756e-16, 6.077958e-16, 6.08342e-16, 6.098928e-16, 6.112884e-16, 
    6.128091e-16, 6.131813e-16, 6.149542e-16, 6.135103e-16, 6.158915e-16, 
    6.138661e-16, 6.17371e-16, 6.110695e-16, 6.138077e-16, 6.088445e-16, 
    6.093802e-16, 6.103475e-16, 6.125661e-16, 6.113694e-16, 6.127691e-16, 
    6.096757e-16, 6.080674e-16, 6.076517e-16, 6.068747e-16, 6.076695e-16, 
    6.076048e-16, 6.08365e-16, 6.081208e-16, 6.099443e-16, 6.089651e-16, 
    6.11745e-16, 6.127582e-16, 6.156165e-16, 6.173656e-16, 6.191449e-16, 
    6.199294e-16, 6.201682e-16, 6.20268e-16 ;

 CWDC_TO_LITR2C =
  4.567303e-16, 4.579685e-16, 4.57728e-16, 4.587258e-16, 4.581726e-16, 
    4.588256e-16, 4.569816e-16, 4.580175e-16, 4.573564e-16, 4.568421e-16, 
    4.606592e-16, 4.587703e-16, 4.626199e-16, 4.614172e-16, 4.644362e-16, 
    4.624325e-16, 4.648399e-16, 4.643788e-16, 4.65767e-16, 4.653695e-16, 
    4.671423e-16, 4.659504e-16, 4.680609e-16, 4.66858e-16, 4.670461e-16, 
    4.65911e-16, 4.591511e-16, 4.604241e-16, 4.590756e-16, 4.592572e-16, 
    4.591758e-16, 4.581838e-16, 4.576834e-16, 4.566359e-16, 4.568263e-16, 
    4.575957e-16, 4.593389e-16, 4.587477e-16, 4.602378e-16, 4.602042e-16, 
    4.618608e-16, 4.611141e-16, 4.63895e-16, 4.631056e-16, 4.653862e-16, 
    4.648129e-16, 4.653591e-16, 4.651936e-16, 4.653613e-16, 4.645205e-16, 
    4.648808e-16, 4.641408e-16, 4.61254e-16, 4.621031e-16, 4.595686e-16, 
    4.580414e-16, 4.570271e-16, 4.563064e-16, 4.564083e-16, 4.566025e-16, 
    4.576002e-16, 4.585379e-16, 4.592519e-16, 4.597292e-16, 4.601994e-16, 
    4.616203e-16, 4.623726e-16, 4.640544e-16, 4.637514e-16, 4.64265e-16, 
    4.647559e-16, 4.655791e-16, 4.654437e-16, 4.658062e-16, 4.642517e-16, 
    4.652849e-16, 4.635789e-16, 4.640455e-16, 4.603257e-16, 4.589073e-16, 
    4.583026e-16, 4.577742e-16, 4.564866e-16, 4.573759e-16, 4.570254e-16, 
    4.578594e-16, 4.583888e-16, 4.581271e-16, 4.597423e-16, 4.591145e-16, 
    4.624172e-16, 4.609958e-16, 4.646986e-16, 4.638136e-16, 4.649107e-16, 
    4.643511e-16, 4.653097e-16, 4.64447e-16, 4.659412e-16, 4.662661e-16, 
    4.66044e-16, 4.668974e-16, 4.643991e-16, 4.65359e-16, 4.581197e-16, 
    4.581623e-16, 4.583614e-16, 4.574863e-16, 4.574328e-16, 4.566306e-16, 
    4.573445e-16, 4.576483e-16, 4.584196e-16, 4.588754e-16, 4.593085e-16, 
    4.602604e-16, 4.613224e-16, 4.628062e-16, 4.63871e-16, 4.645843e-16, 
    4.641471e-16, 4.645331e-16, 4.641015e-16, 4.638992e-16, 4.661443e-16, 
    4.64884e-16, 4.667747e-16, 4.666702e-16, 4.658148e-16, 4.66682e-16, 
    4.581924e-16, 4.579466e-16, 4.570927e-16, 4.57761e-16, 4.565433e-16, 
    4.572249e-16, 4.576165e-16, 4.591273e-16, 4.594594e-16, 4.597667e-16, 
    4.603738e-16, 4.611524e-16, 4.625167e-16, 4.637026e-16, 4.647845e-16, 
    4.647053e-16, 4.647331e-16, 4.649746e-16, 4.643763e-16, 4.650728e-16, 
    4.651895e-16, 4.648841e-16, 4.666562e-16, 4.661502e-16, 4.66668e-16, 
    4.663386e-16, 4.580266e-16, 4.5844e-16, 4.582166e-16, 4.586366e-16, 
    4.583406e-16, 4.596559e-16, 4.600499e-16, 4.618924e-16, 4.61137e-16, 
    4.623395e-16, 4.612593e-16, 4.614507e-16, 4.623781e-16, 4.613178e-16, 
    4.636372e-16, 4.620646e-16, 4.649839e-16, 4.634151e-16, 4.650822e-16, 
    4.647798e-16, 4.652805e-16, 4.657286e-16, 4.662924e-16, 4.673315e-16, 
    4.67091e-16, 4.679597e-16, 4.590562e-16, 4.595919e-16, 4.59545e-16, 
    4.601056e-16, 4.605199e-16, 4.614178e-16, 4.62856e-16, 4.623155e-16, 
    4.63308e-16, 4.63507e-16, 4.619992e-16, 4.629249e-16, 4.599505e-16, 
    4.604313e-16, 4.601452e-16, 4.590984e-16, 4.624396e-16, 4.607259e-16, 
    4.638885e-16, 4.629619e-16, 4.656647e-16, 4.643209e-16, 4.669586e-16, 
    4.680835e-16, 4.691426e-16, 4.703775e-16, 4.598845e-16, 4.595206e-16, 
    4.601723e-16, 4.610729e-16, 4.619087e-16, 4.630184e-16, 4.63132e-16, 
    4.633397e-16, 4.638776e-16, 4.643297e-16, 4.634051e-16, 4.64443e-16, 
    4.605422e-16, 4.625884e-16, 4.593827e-16, 4.603486e-16, 4.6102e-16, 
    4.607258e-16, 4.622537e-16, 4.626134e-16, 4.640738e-16, 4.633194e-16, 
    4.678058e-16, 4.658229e-16, 4.713177e-16, 4.697846e-16, 4.593933e-16, 
    4.598834e-16, 4.615867e-16, 4.607766e-16, 4.630926e-16, 4.636619e-16, 
    4.641244e-16, 4.647153e-16, 4.647793e-16, 4.651292e-16, 4.645556e-16, 
    4.651067e-16, 4.630208e-16, 4.639533e-16, 4.613925e-16, 4.620162e-16, 
    4.617294e-16, 4.614145e-16, 4.62386e-16, 4.634196e-16, 4.634421e-16, 
    4.63773e-16, 4.647049e-16, 4.63102e-16, 4.680606e-16, 4.649999e-16, 
    4.604174e-16, 4.613596e-16, 4.614947e-16, 4.611297e-16, 4.636048e-16, 
    4.627085e-16, 4.651208e-16, 4.644694e-16, 4.655366e-16, 4.650063e-16, 
    4.649283e-16, 4.64247e-16, 4.638224e-16, 4.627496e-16, 4.618758e-16, 
    4.611827e-16, 4.61344e-16, 4.621052e-16, 4.634829e-16, 4.647849e-16, 
    4.644996e-16, 4.654556e-16, 4.629248e-16, 4.639863e-16, 4.635762e-16, 
    4.646457e-16, 4.62301e-16, 4.642966e-16, 4.617901e-16, 4.620102e-16, 
    4.626907e-16, 4.64058e-16, 4.643609e-16, 4.646836e-16, 4.644846e-16, 
    4.63518e-16, 4.633597e-16, 4.626743e-16, 4.624848e-16, 4.619623e-16, 
    4.615294e-16, 4.619249e-16, 4.623399e-16, 4.635186e-16, 4.645792e-16, 
    4.657349e-16, 4.660178e-16, 4.673652e-16, 4.662678e-16, 4.680775e-16, 
    4.665382e-16, 4.69202e-16, 4.644128e-16, 4.664938e-16, 4.627218e-16, 
    4.631289e-16, 4.638641e-16, 4.655502e-16, 4.646407e-16, 4.657045e-16, 
    4.633535e-16, 4.621312e-16, 4.618153e-16, 4.612248e-16, 4.618288e-16, 
    4.617797e-16, 4.623574e-16, 4.621718e-16, 4.635577e-16, 4.628135e-16, 
    4.649262e-16, 4.656962e-16, 4.678685e-16, 4.691979e-16, 4.705501e-16, 
    4.711464e-16, 4.713278e-16, 4.714036e-16 ;

 CWDC_TO_LITR3C =
  1.442306e-16, 1.446217e-16, 1.445457e-16, 1.448608e-16, 1.446861e-16, 
    1.448923e-16, 1.4431e-16, 1.446371e-16, 1.444284e-16, 1.442659e-16, 
    1.454713e-16, 1.448748e-16, 1.460905e-16, 1.457107e-16, 1.466641e-16, 
    1.460313e-16, 1.467916e-16, 1.46646e-16, 1.470843e-16, 1.469588e-16, 
    1.475186e-16, 1.471422e-16, 1.478087e-16, 1.474289e-16, 1.474882e-16, 
    1.471298e-16, 1.449951e-16, 1.453971e-16, 1.449712e-16, 1.450286e-16, 
    1.450029e-16, 1.446896e-16, 1.445316e-16, 1.442008e-16, 1.442609e-16, 
    1.445039e-16, 1.450544e-16, 1.448677e-16, 1.453383e-16, 1.453277e-16, 
    1.458508e-16, 1.45615e-16, 1.464932e-16, 1.462439e-16, 1.46964e-16, 
    1.46783e-16, 1.469555e-16, 1.469032e-16, 1.469562e-16, 1.466907e-16, 
    1.468045e-16, 1.465708e-16, 1.456591e-16, 1.459273e-16, 1.451269e-16, 
    1.446447e-16, 1.443243e-16, 1.440968e-16, 1.441289e-16, 1.441902e-16, 
    1.445053e-16, 1.448014e-16, 1.450269e-16, 1.451776e-16, 1.453261e-16, 
    1.457748e-16, 1.460124e-16, 1.465435e-16, 1.464478e-16, 1.4661e-16, 
    1.46765e-16, 1.47025e-16, 1.469822e-16, 1.470967e-16, 1.466058e-16, 
    1.469321e-16, 1.463933e-16, 1.465407e-16, 1.45366e-16, 1.449181e-16, 
    1.447271e-16, 1.445603e-16, 1.441537e-16, 1.444345e-16, 1.443238e-16, 
    1.445872e-16, 1.447544e-16, 1.446717e-16, 1.451818e-16, 1.449835e-16, 
    1.460265e-16, 1.455776e-16, 1.467469e-16, 1.464675e-16, 1.468139e-16, 
    1.466372e-16, 1.469399e-16, 1.466675e-16, 1.471393e-16, 1.472419e-16, 
    1.471718e-16, 1.474413e-16, 1.466523e-16, 1.469555e-16, 1.446694e-16, 
    1.446828e-16, 1.447457e-16, 1.444693e-16, 1.444525e-16, 1.441992e-16, 
    1.444246e-16, 1.445205e-16, 1.447641e-16, 1.44908e-16, 1.450448e-16, 
    1.453454e-16, 1.456808e-16, 1.461493e-16, 1.464856e-16, 1.467108e-16, 
    1.465728e-16, 1.466947e-16, 1.465584e-16, 1.464945e-16, 1.472035e-16, 
    1.468055e-16, 1.474025e-16, 1.473695e-16, 1.470994e-16, 1.473733e-16, 
    1.446923e-16, 1.446147e-16, 1.443451e-16, 1.445561e-16, 1.441716e-16, 
    1.443868e-16, 1.445105e-16, 1.449876e-16, 1.450924e-16, 1.451895e-16, 
    1.453812e-16, 1.456271e-16, 1.460579e-16, 1.464324e-16, 1.46774e-16, 
    1.46749e-16, 1.467578e-16, 1.468341e-16, 1.466451e-16, 1.468651e-16, 
    1.469019e-16, 1.468055e-16, 1.473651e-16, 1.472053e-16, 1.473688e-16, 
    1.472648e-16, 1.4464e-16, 1.447705e-16, 1.447e-16, 1.448326e-16, 
    1.447391e-16, 1.451545e-16, 1.452789e-16, 1.458608e-16, 1.456222e-16, 
    1.460019e-16, 1.456608e-16, 1.457213e-16, 1.460141e-16, 1.456793e-16, 
    1.464117e-16, 1.459151e-16, 1.46837e-16, 1.463416e-16, 1.46868e-16, 
    1.467726e-16, 1.469307e-16, 1.470722e-16, 1.472502e-16, 1.475784e-16, 
    1.475024e-16, 1.477767e-16, 1.449651e-16, 1.451343e-16, 1.451195e-16, 
    1.452965e-16, 1.454273e-16, 1.457109e-16, 1.461651e-16, 1.459943e-16, 
    1.463078e-16, 1.463706e-16, 1.458945e-16, 1.461868e-16, 1.452475e-16, 
    1.453994e-16, 1.45309e-16, 1.449784e-16, 1.460336e-16, 1.454924e-16, 
    1.464911e-16, 1.461985e-16, 1.47052e-16, 1.466277e-16, 1.474606e-16, 
    1.478159e-16, 1.481503e-16, 1.485403e-16, 1.452267e-16, 1.451118e-16, 
    1.453176e-16, 1.45602e-16, 1.458659e-16, 1.462163e-16, 1.462522e-16, 
    1.463178e-16, 1.464877e-16, 1.466304e-16, 1.463385e-16, 1.466662e-16, 
    1.454344e-16, 1.460806e-16, 1.450682e-16, 1.453732e-16, 1.455852e-16, 
    1.454923e-16, 1.459749e-16, 1.460885e-16, 1.465496e-16, 1.463114e-16, 
    1.477281e-16, 1.47102e-16, 1.488372e-16, 1.483531e-16, 1.450716e-16, 
    1.452263e-16, 1.457642e-16, 1.455084e-16, 1.462398e-16, 1.464195e-16, 
    1.465656e-16, 1.467522e-16, 1.467724e-16, 1.468829e-16, 1.467018e-16, 
    1.468758e-16, 1.462171e-16, 1.465116e-16, 1.457029e-16, 1.458998e-16, 
    1.458093e-16, 1.457099e-16, 1.460166e-16, 1.46343e-16, 1.463502e-16, 
    1.464546e-16, 1.467489e-16, 1.462427e-16, 1.478086e-16, 1.468421e-16, 
    1.45395e-16, 1.456925e-16, 1.457352e-16, 1.456199e-16, 1.464015e-16, 
    1.461185e-16, 1.468802e-16, 1.466745e-16, 1.470116e-16, 1.468441e-16, 
    1.468195e-16, 1.466043e-16, 1.464702e-16, 1.461314e-16, 1.458555e-16, 
    1.456366e-16, 1.456876e-16, 1.459279e-16, 1.46363e-16, 1.467742e-16, 
    1.466841e-16, 1.46986e-16, 1.461868e-16, 1.46522e-16, 1.463925e-16, 
    1.467302e-16, 1.459898e-16, 1.4662e-16, 1.458285e-16, 1.45898e-16, 
    1.461129e-16, 1.465446e-16, 1.466403e-16, 1.467422e-16, 1.466793e-16, 
    1.463741e-16, 1.463241e-16, 1.461077e-16, 1.460478e-16, 1.458828e-16, 
    1.457461e-16, 1.45871e-16, 1.460021e-16, 1.463743e-16, 1.467092e-16, 
    1.470742e-16, 1.471635e-16, 1.47589e-16, 1.472425e-16, 1.478139e-16, 
    1.473279e-16, 1.48169e-16, 1.466567e-16, 1.473138e-16, 1.461227e-16, 
    1.462512e-16, 1.464834e-16, 1.470159e-16, 1.467286e-16, 1.470646e-16, 
    1.463222e-16, 1.459362e-16, 1.458364e-16, 1.456499e-16, 1.458407e-16, 
    1.458252e-16, 1.460076e-16, 1.45949e-16, 1.463866e-16, 1.461516e-16, 
    1.468188e-16, 1.47062e-16, 1.47748e-16, 1.481677e-16, 1.485948e-16, 
    1.487831e-16, 1.488404e-16, 1.488643e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  9.134606e-19, 9.159371e-19, 9.154561e-19, 9.174516e-19, 9.163451e-19, 
    9.176513e-19, 9.139633e-19, 9.16035e-19, 9.147129e-19, 9.136843e-19, 
    9.213184e-19, 9.175407e-19, 9.252397e-19, 9.228345e-19, 9.288723e-19, 
    9.248651e-19, 9.296798e-19, 9.287577e-19, 9.31534e-19, 9.307391e-19, 
    9.342847e-19, 9.319009e-19, 9.361219e-19, 9.337161e-19, 9.340923e-19, 
    9.318221e-19, 9.183022e-19, 9.208482e-19, 9.18151e-19, 9.185144e-19, 
    9.183515e-19, 9.163677e-19, 9.153669e-19, 9.132718e-19, 9.136525e-19, 
    9.151914e-19, 9.186777e-19, 9.174954e-19, 9.204757e-19, 9.204085e-19, 
    9.237215e-19, 9.222283e-19, 9.2779e-19, 9.262112e-19, 9.307723e-19, 
    9.296258e-19, 9.307183e-19, 9.303871e-19, 9.307225e-19, 9.29041e-19, 
    9.297616e-19, 9.282815e-19, 9.225079e-19, 9.242061e-19, 9.191371e-19, 
    9.160828e-19, 9.14054e-19, 9.126129e-19, 9.128167e-19, 9.132049e-19, 
    9.152004e-19, 9.170758e-19, 9.185038e-19, 9.194584e-19, 9.203988e-19, 
    9.232406e-19, 9.247452e-19, 9.281087e-19, 9.275027e-19, 9.285299e-19, 
    9.295117e-19, 9.311582e-19, 9.308875e-19, 9.316124e-19, 9.285033e-19, 
    9.305698e-19, 9.271578e-19, 9.280911e-19, 9.206515e-19, 9.178146e-19, 
    9.166052e-19, 9.155484e-19, 9.129732e-19, 9.147517e-19, 9.140507e-19, 
    9.157188e-19, 9.167777e-19, 9.162541e-19, 9.194846e-19, 9.18229e-19, 
    9.248344e-19, 9.219915e-19, 9.293972e-19, 9.276272e-19, 9.298214e-19, 
    9.287021e-19, 9.306193e-19, 9.288939e-19, 9.318823e-19, 9.325322e-19, 
    9.320881e-19, 9.337948e-19, 9.287982e-19, 9.30718e-19, 9.162393e-19, 
    9.163247e-19, 9.167227e-19, 9.149725e-19, 9.148656e-19, 9.132613e-19, 
    9.146891e-19, 9.152965e-19, 9.168392e-19, 9.177508e-19, 9.186172e-19, 
    9.205209e-19, 9.226448e-19, 9.256123e-19, 9.27742e-19, 9.291686e-19, 
    9.282941e-19, 9.290662e-19, 9.282029e-19, 9.277983e-19, 9.322886e-19, 
    9.297681e-19, 9.335493e-19, 9.333404e-19, 9.316295e-19, 9.333639e-19, 
    9.163847e-19, 9.158933e-19, 9.141853e-19, 9.155221e-19, 9.130865e-19, 
    9.144498e-19, 9.152331e-19, 9.182546e-19, 9.189188e-19, 9.195335e-19, 
    9.207477e-19, 9.223047e-19, 9.250335e-19, 9.274051e-19, 9.295689e-19, 
    9.294105e-19, 9.294663e-19, 9.299491e-19, 9.287525e-19, 9.301456e-19, 
    9.303789e-19, 9.297682e-19, 9.333123e-19, 9.323004e-19, 9.333359e-19, 
    9.326772e-19, 9.160531e-19, 9.1688e-19, 9.164332e-19, 9.172732e-19, 
    9.166811e-19, 9.193117e-19, 9.200998e-19, 9.237849e-19, 9.222739e-19, 
    9.246789e-19, 9.225186e-19, 9.229013e-19, 9.247561e-19, 9.226356e-19, 
    9.272743e-19, 9.241293e-19, 9.299679e-19, 9.268301e-19, 9.301643e-19, 
    9.295596e-19, 9.30561e-19, 9.314573e-19, 9.325848e-19, 9.34663e-19, 
    9.34182e-19, 9.359194e-19, 9.181125e-19, 9.191839e-19, 9.190901e-19, 
    9.202111e-19, 9.210398e-19, 9.228355e-19, 9.25712e-19, 9.246309e-19, 
    9.266159e-19, 9.27014e-19, 9.239985e-19, 9.258499e-19, 9.199009e-19, 
    9.208625e-19, 9.202905e-19, 9.181967e-19, 9.248793e-19, 9.214518e-19, 
    9.27777e-19, 9.259239e-19, 9.313294e-19, 9.286419e-19, 9.339171e-19, 
    9.36167e-19, 9.382852e-19, 9.407549e-19, 9.197689e-19, 9.190412e-19, 
    9.203446e-19, 9.221458e-19, 9.238173e-19, 9.260369e-19, 9.262641e-19, 
    9.266795e-19, 9.277552e-19, 9.286594e-19, 9.268103e-19, 9.288861e-19, 
    9.210844e-19, 9.251769e-19, 9.187654e-19, 9.206972e-19, 9.220399e-19, 
    9.214516e-19, 9.245074e-19, 9.25227e-19, 9.281476e-19, 9.266388e-19, 
    9.356115e-19, 9.316458e-19, 9.426354e-19, 9.395693e-19, 9.187866e-19, 
    9.197666e-19, 9.231735e-19, 9.215532e-19, 9.261852e-19, 9.273238e-19, 
    9.282487e-19, 9.294306e-19, 9.295585e-19, 9.302585e-19, 9.291113e-19, 
    9.302134e-19, 9.260415e-19, 9.279066e-19, 9.227849e-19, 9.240323e-19, 
    9.234587e-19, 9.228291e-19, 9.247719e-19, 9.268392e-19, 9.268843e-19, 
    9.275461e-19, 9.294099e-19, 9.26204e-19, 9.361211e-19, 9.299997e-19, 
    9.208348e-19, 9.227192e-19, 9.229893e-19, 9.222594e-19, 9.272096e-19, 
    9.25417e-19, 9.302415e-19, 9.289386e-19, 9.310733e-19, 9.300127e-19, 
    9.298566e-19, 9.284939e-19, 9.276448e-19, 9.254991e-19, 9.237516e-19, 
    9.223654e-19, 9.226879e-19, 9.242103e-19, 9.269658e-19, 9.295698e-19, 
    9.289993e-19, 9.309111e-19, 9.258496e-19, 9.279726e-19, 9.271523e-19, 
    9.292915e-19, 9.246019e-19, 9.285932e-19, 9.235802e-19, 9.240204e-19, 
    9.253814e-19, 9.281159e-19, 9.287219e-19, 9.293672e-19, 9.289692e-19, 
    9.270359e-19, 9.267193e-19, 9.253485e-19, 9.249696e-19, 9.239247e-19, 
    9.230588e-19, 9.238497e-19, 9.246798e-19, 9.270371e-19, 9.291584e-19, 
    9.314699e-19, 9.320356e-19, 9.347304e-19, 9.325357e-19, 9.36155e-19, 
    9.330764e-19, 9.384039e-19, 9.288256e-19, 9.329877e-19, 9.254437e-19, 
    9.262578e-19, 9.277282e-19, 9.311005e-19, 9.292815e-19, 9.31409e-19, 
    9.26707e-19, 9.242624e-19, 9.236306e-19, 9.224496e-19, 9.236576e-19, 
    9.235594e-19, 9.247148e-19, 9.243436e-19, 9.271153e-19, 9.256269e-19, 
    9.298524e-19, 9.313924e-19, 9.35737e-19, 9.383957e-19, 9.411003e-19, 
    9.422927e-19, 9.426556e-19, 9.428073e-19 ;

 CWDN_TO_LITR3N =
  2.884613e-19, 2.892433e-19, 2.890914e-19, 2.897216e-19, 2.893722e-19, 
    2.897846e-19, 2.8862e-19, 2.892742e-19, 2.888567e-19, 2.885319e-19, 
    2.909427e-19, 2.897497e-19, 2.921809e-19, 2.914214e-19, 2.933281e-19, 
    2.920626e-19, 2.935831e-19, 2.932919e-19, 2.941686e-19, 2.939176e-19, 
    2.950373e-19, 2.942845e-19, 2.956174e-19, 2.948577e-19, 2.949765e-19, 
    2.942596e-19, 2.899902e-19, 2.907942e-19, 2.899424e-19, 2.900572e-19, 
    2.900057e-19, 2.893793e-19, 2.890632e-19, 2.884016e-19, 2.885218e-19, 
    2.890078e-19, 2.901088e-19, 2.897354e-19, 2.906765e-19, 2.906553e-19, 
    2.917015e-19, 2.9123e-19, 2.929863e-19, 2.924877e-19, 2.939281e-19, 
    2.93566e-19, 2.93911e-19, 2.938065e-19, 2.939124e-19, 2.933813e-19, 
    2.936089e-19, 2.931415e-19, 2.913183e-19, 2.918545e-19, 2.902538e-19, 
    2.892893e-19, 2.886487e-19, 2.881935e-19, 2.882579e-19, 2.883805e-19, 
    2.890107e-19, 2.896029e-19, 2.900538e-19, 2.903553e-19, 2.906522e-19, 
    2.915497e-19, 2.920248e-19, 2.93087e-19, 2.928956e-19, 2.9322e-19, 
    2.9353e-19, 2.9405e-19, 2.939645e-19, 2.941934e-19, 2.932116e-19, 
    2.938642e-19, 2.927867e-19, 2.930814e-19, 2.90732e-19, 2.898362e-19, 
    2.894543e-19, 2.891206e-19, 2.883073e-19, 2.88869e-19, 2.886476e-19, 
    2.891744e-19, 2.895087e-19, 2.893434e-19, 2.903635e-19, 2.899671e-19, 
    2.92053e-19, 2.911552e-19, 2.934939e-19, 2.929349e-19, 2.936278e-19, 
    2.932744e-19, 2.938798e-19, 2.933349e-19, 2.942787e-19, 2.944839e-19, 
    2.943436e-19, 2.948825e-19, 2.933047e-19, 2.939109e-19, 2.893387e-19, 
    2.893657e-19, 2.894914e-19, 2.889387e-19, 2.889049e-19, 2.883983e-19, 
    2.888492e-19, 2.89041e-19, 2.895282e-19, 2.89816e-19, 2.900896e-19, 
    2.906908e-19, 2.913615e-19, 2.922986e-19, 2.929711e-19, 2.934217e-19, 
    2.931455e-19, 2.933893e-19, 2.931167e-19, 2.92989e-19, 2.944069e-19, 
    2.93611e-19, 2.948051e-19, 2.947391e-19, 2.941988e-19, 2.947465e-19, 
    2.893846e-19, 2.892294e-19, 2.886901e-19, 2.891122e-19, 2.883431e-19, 
    2.887736e-19, 2.89021e-19, 2.899752e-19, 2.901849e-19, 2.90379e-19, 
    2.907624e-19, 2.912541e-19, 2.921158e-19, 2.928648e-19, 2.935481e-19, 
    2.934981e-19, 2.935157e-19, 2.936681e-19, 2.932903e-19, 2.937302e-19, 
    2.938039e-19, 2.93611e-19, 2.947302e-19, 2.944107e-19, 2.947377e-19, 
    2.945296e-19, 2.892799e-19, 2.895411e-19, 2.893999e-19, 2.896652e-19, 
    2.894783e-19, 2.90309e-19, 2.905578e-19, 2.917215e-19, 2.912444e-19, 
    2.920039e-19, 2.913217e-19, 2.914425e-19, 2.920283e-19, 2.913586e-19, 
    2.928235e-19, 2.918303e-19, 2.936741e-19, 2.926832e-19, 2.937361e-19, 
    2.935451e-19, 2.938614e-19, 2.941444e-19, 2.945005e-19, 2.951567e-19, 
    2.950048e-19, 2.955535e-19, 2.899303e-19, 2.902686e-19, 2.90239e-19, 
    2.90593e-19, 2.908547e-19, 2.914217e-19, 2.923301e-19, 2.919887e-19, 
    2.926156e-19, 2.927413e-19, 2.91789e-19, 2.923737e-19, 2.904951e-19, 
    2.907987e-19, 2.90618e-19, 2.899569e-19, 2.920672e-19, 2.909848e-19, 
    2.929822e-19, 2.92397e-19, 2.94104e-19, 2.932553e-19, 2.949212e-19, 
    2.956317e-19, 2.963006e-19, 2.970805e-19, 2.904534e-19, 2.902235e-19, 
    2.906351e-19, 2.912039e-19, 2.917318e-19, 2.924327e-19, 2.925045e-19, 
    2.926356e-19, 2.929753e-19, 2.932609e-19, 2.926769e-19, 2.933325e-19, 
    2.908688e-19, 2.921611e-19, 2.901364e-19, 2.907465e-19, 2.911705e-19, 
    2.909847e-19, 2.919497e-19, 2.921769e-19, 2.930992e-19, 2.926228e-19, 
    2.954562e-19, 2.942039e-19, 2.976743e-19, 2.967061e-19, 2.901432e-19, 
    2.904526e-19, 2.915285e-19, 2.910168e-19, 2.924795e-19, 2.928391e-19, 
    2.931312e-19, 2.935044e-19, 2.935448e-19, 2.937658e-19, 2.934036e-19, 
    2.937516e-19, 2.924342e-19, 2.930231e-19, 2.914058e-19, 2.917997e-19, 
    2.916185e-19, 2.914197e-19, 2.920332e-19, 2.926861e-19, 2.927003e-19, 
    2.929093e-19, 2.934978e-19, 2.924855e-19, 2.956172e-19, 2.936841e-19, 
    2.907899e-19, 2.91385e-19, 2.914703e-19, 2.912398e-19, 2.92803e-19, 
    2.92237e-19, 2.937605e-19, 2.933491e-19, 2.940231e-19, 2.936882e-19, 
    2.936389e-19, 2.932086e-19, 2.929405e-19, 2.922629e-19, 2.91711e-19, 
    2.912733e-19, 2.913751e-19, 2.918559e-19, 2.927261e-19, 2.935483e-19, 
    2.933682e-19, 2.939719e-19, 2.923736e-19, 2.93044e-19, 2.927849e-19, 
    2.934605e-19, 2.919796e-19, 2.932399e-19, 2.916569e-19, 2.917959e-19, 
    2.922257e-19, 2.930892e-19, 2.932806e-19, 2.934844e-19, 2.933587e-19, 
    2.927482e-19, 2.926482e-19, 2.922154e-19, 2.920956e-19, 2.917657e-19, 
    2.914923e-19, 2.91742e-19, 2.920041e-19, 2.927486e-19, 2.934184e-19, 
    2.941484e-19, 2.94327e-19, 2.95178e-19, 2.94485e-19, 2.956279e-19, 
    2.946557e-19, 2.963381e-19, 2.933133e-19, 2.946277e-19, 2.922454e-19, 
    2.925025e-19, 2.929668e-19, 2.940317e-19, 2.934573e-19, 2.941292e-19, 
    2.926443e-19, 2.918723e-19, 2.916728e-19, 2.912998e-19, 2.916813e-19, 
    2.916503e-19, 2.920152e-19, 2.91898e-19, 2.927733e-19, 2.923032e-19, 
    2.936376e-19, 2.941239e-19, 2.954959e-19, 2.963355e-19, 2.971896e-19, 
    2.975661e-19, 2.976807e-19, 2.977286e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.809097e-14, 2.821622e-14, 2.819179e-14, 2.829291e-14, 2.823676e-14, 
    2.830296e-14, 2.81162e-14, 2.822105e-14, 2.815406e-14, 2.810199e-14, 
    2.848918e-14, 2.829722e-14, 2.868855e-14, 2.856595e-14, 2.887388e-14, 
    2.866944e-14, 2.89151e-14, 2.886786e-14, 2.90098e-14, 2.896908e-14, 
    2.915086e-14, 2.902851e-14, 2.924503e-14, 2.912156e-14, 2.914086e-14, 
    2.902437e-14, 2.833595e-14, 2.846547e-14, 2.832824e-14, 2.834671e-14, 
    2.833838e-14, 2.823783e-14, 2.818724e-14, 2.808113e-14, 2.810034e-14, 
    2.817823e-14, 2.835483e-14, 2.829477e-14, 2.844593e-14, 2.844252e-14, 
    2.861098e-14, 2.853498e-14, 2.88184e-14, 2.873774e-14, 2.897075e-14, 
    2.891209e-14, 2.896796e-14, 2.895097e-14, 2.896811e-14, 2.888214e-14, 
    2.891892e-14, 2.884328e-14, 2.854952e-14, 2.863594e-14, 2.837823e-14, 
    2.822353e-14, 2.812071e-14, 2.804786e-14, 2.80581e-14, 2.807775e-14, 
    2.817864e-14, 2.827349e-14, 2.834585e-14, 2.839425e-14, 2.844195e-14, 
    2.858668e-14, 2.866317e-14, 2.883468e-14, 2.880365e-14, 2.885613e-14, 
    2.890623e-14, 2.899042e-14, 2.897654e-14, 2.901363e-14, 2.885457e-14, 
    2.896027e-14, 2.878577e-14, 2.883348e-14, 2.845539e-14, 2.831106e-14, 
    2.824994e-14, 2.819627e-14, 2.806601e-14, 2.815595e-14, 2.812046e-14, 
    2.820474e-14, 2.825836e-14, 2.823179e-14, 2.839555e-14, 2.833183e-14, 
    2.866767e-14, 2.852292e-14, 2.890042e-14, 2.880996e-14, 2.892201e-14, 
    2.886481e-14, 2.896281e-14, 2.887456e-14, 2.902739e-14, 2.906072e-14, 
    2.90379e-14, 2.912532e-14, 2.886952e-14, 2.896773e-14, 2.82312e-14, 
    2.823553e-14, 2.825565e-14, 2.816708e-14, 2.816164e-14, 2.808047e-14, 
    2.815261e-14, 2.818338e-14, 2.826139e-14, 2.830757e-14, 2.835147e-14, 
    2.844812e-14, 2.855611e-14, 2.870719e-14, 2.881579e-14, 2.88886e-14, 
    2.88439e-14, 2.888332e-14, 2.883921e-14, 2.88185e-14, 2.904817e-14, 
    2.891918e-14, 2.911267e-14, 2.910196e-14, 2.901433e-14, 2.910309e-14, 
    2.823852e-14, 2.821358e-14, 2.812721e-14, 2.819475e-14, 2.807158e-14, 
    2.814053e-14, 2.818016e-14, 2.833317e-14, 2.836674e-14, 2.839796e-14, 
    2.845957e-14, 2.853869e-14, 2.867764e-14, 2.879857e-14, 2.890903e-14, 
    2.89009e-14, 2.890374e-14, 2.892841e-14, 2.886723e-14, 2.89384e-14, 
    2.895034e-14, 2.891907e-14, 2.910045e-14, 2.90486e-14, 2.910163e-14, 
    2.906782e-14, 2.822164e-14, 2.82635e-14, 2.824083e-14, 2.828342e-14, 
    2.825338e-14, 2.838682e-14, 2.842682e-14, 2.861415e-14, 2.853714e-14, 
    2.865961e-14, 2.854951e-14, 2.856902e-14, 2.866361e-14, 2.855537e-14, 
    2.879187e-14, 2.863153e-14, 2.892934e-14, 2.876919e-14, 2.893933e-14, 
    2.890835e-14, 2.895953e-14, 2.900544e-14, 2.906311e-14, 2.916972e-14, 
    2.914496e-14, 2.923413e-14, 2.832594e-14, 2.83803e-14, 2.837546e-14, 
    2.843234e-14, 2.847443e-14, 2.856571e-14, 2.871221e-14, 2.865704e-14, 
    2.875819e-14, 2.877853e-14, 2.862474e-14, 2.871916e-14, 2.841643e-14, 
    2.84653e-14, 2.843614e-14, 2.832987e-14, 2.866959e-14, 2.849514e-14, 
    2.881729e-14, 2.872266e-14, 2.899883e-14, 2.886146e-14, 2.913136e-14, 
    2.924698e-14, 2.935564e-14, 2.94829e-14, 2.840992e-14, 2.837292e-14, 
    2.843905e-14, 2.853071e-14, 2.861563e-14, 2.872874e-14, 2.874026e-14, 
    2.876143e-14, 2.881629e-14, 2.886249e-14, 2.876811e-14, 2.8874e-14, 
    2.84767e-14, 2.868471e-14, 2.835865e-14, 2.845682e-14, 2.852494e-14, 
    2.8495e-14, 2.865041e-14, 2.868704e-14, 2.883612e-14, 2.8759e-14, 
    2.92184e-14, 2.901501e-14, 2.957969e-14, 2.942175e-14, 2.835999e-14, 
    2.840967e-14, 2.858288e-14, 2.850043e-14, 2.87362e-14, 2.879431e-14, 
    2.884148e-14, 2.890193e-14, 2.890837e-14, 2.89442e-14, 2.888545e-14, 
    2.894181e-14, 2.872871e-14, 2.882388e-14, 2.856275e-14, 2.862625e-14, 
    2.859699e-14, 2.856491e-14, 2.86638e-14, 2.876933e-14, 2.877149e-14, 
    2.880531e-14, 2.890086e-14, 2.873669e-14, 2.92447e-14, 2.893087e-14, 
    2.846389e-14, 2.85598e-14, 2.85734e-14, 2.853624e-14, 2.878842e-14, 
    2.8697e-14, 2.894331e-14, 2.887665e-14, 2.898578e-14, 2.893154e-14, 
    2.892351e-14, 2.885385e-14, 2.881046e-14, 2.8701e-14, 2.861192e-14, 
    2.854133e-14, 2.855768e-14, 2.863524e-14, 2.87757e-14, 2.890868e-14, 
    2.887952e-14, 2.897716e-14, 2.871858e-14, 2.882699e-14, 2.878505e-14, 
    2.889428e-14, 2.865549e-14, 2.885945e-14, 2.860339e-14, 2.862577e-14, 
    2.869511e-14, 2.883476e-14, 2.886552e-14, 2.889856e-14, 2.887811e-14, 
    2.877944e-14, 2.876322e-14, 2.869324e-14, 2.867394e-14, 2.862066e-14, 
    2.857653e-14, 2.861682e-14, 2.865909e-14, 2.877926e-14, 2.888761e-14, 
    2.900579e-14, 2.90347e-14, 2.917306e-14, 2.906047e-14, 2.924633e-14, 
    2.908839e-14, 2.936175e-14, 2.887111e-14, 2.908413e-14, 2.869825e-14, 
    2.873973e-14, 2.88149e-14, 2.898726e-14, 2.889407e-14, 2.9003e-14, 
    2.876256e-14, 2.863799e-14, 2.860567e-14, 2.85456e-14, 2.8607e-14, 
    2.860201e-14, 2.866081e-14, 2.864186e-14, 2.878318e-14, 2.870724e-14, 
    2.892299e-14, 2.900183e-14, 2.922452e-14, 2.936117e-14, 2.950029e-14, 
    2.956173e-14, 2.958043e-14, 2.958823e-14 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  6.523794, 6.540125, 6.536952, 6.550135, 6.542829, 6.551457, 6.527113, 
    6.540763, 6.532053, 6.525279, 6.575651, 6.550726, 6.601721, 6.585755, 
    6.627564, 6.599216, 6.632985, 6.626819, 6.645467, 6.640121, 6.663968, 
    6.647936, 6.676415, 6.660152, 6.662682, 6.647403, 6.555763, 6.572534, 
    6.554764, 6.557154, 6.556088, 6.54297, 6.536342, 6.522566, 6.52507, 
    6.535199, 6.55823, 6.550441, 6.570138, 6.569693, 6.591645, 6.581743, 
    6.620341, 6.608221, 6.640345, 6.632642, 6.639977, 6.637756, 6.640007, 
    6.628716, 6.633549, 6.623633, 6.583592, 6.59486, 6.561271, 6.541056, 
    6.527707, 6.51823, 6.519569, 6.522116, 6.535258, 6.547664, 6.5571, 
    6.563406, 6.569628, 6.58841, 6.598429, 6.622461, 6.618424, 6.625282, 
    6.631878, 6.642933, 6.641116, 6.645985, 6.625119, 6.63897, 6.614541, 
    6.622359, 6.571227, 6.552548, 6.544515, 6.537559, 6.520597, 6.5323, 
    6.527681, 6.538696, 6.545691, 6.542234, 6.563578, 6.555283, 6.599024, 
    6.580162, 6.631109, 6.619255, 6.633957, 6.626454, 6.639307, 6.627739, 
    6.647806, 6.652172, 6.649186, 6.6607, 6.627095, 6.639968, 6.542132, 
    6.542696, 6.545331, 6.533754, 6.533053, 6.522493, 6.531897, 6.535898, 
    6.546104, 6.552127, 6.557842, 6.57043, 6.584489, 6.604214, 6.620022, 
    6.62958, 6.623724, 6.628893, 6.623111, 6.620407, 6.650529, 6.633588, 
    6.659042, 6.657634, 6.646096, 6.657794, 6.543093, 6.53985, 6.528574, 
    6.537397, 6.521346, 6.530313, 6.535468, 6.555437, 6.559839, 6.563895, 
    6.571935, 6.58225, 6.600362, 6.617761, 6.632266, 6.631204, 6.631577, 
    6.634811, 6.626788, 6.636131, 6.63769, 6.633598, 6.657445, 6.650624, 
    6.657604, 6.653165, 6.540906, 6.546369, 6.543415, 6.548965, 6.545046, 
    6.562413, 6.567619, 6.592047, 6.582041, 6.598, 6.583668, 6.586199, 
    6.59848, 6.584448, 6.615288, 6.594326, 6.634938, 6.612304, 6.636257, 
    6.632203, 6.638927, 6.644943, 6.652539, 6.666549, 6.663306, 6.675056, 
    6.554515, 6.561577, 6.560972, 6.568383, 6.573865, 6.585772, 6.604887, 
    6.597697, 6.610922, 6.613573, 6.593496, 6.605799, 6.566321, 6.572671, 
    6.568903, 6.555061, 6.599329, 6.576578, 6.620254, 6.606301, 6.644083, 
    6.626027, 6.661517, 6.676698, 6.691111, 6.707887, 6.565454, 6.560649, 
    6.56927, 6.581177, 6.592283, 6.607052, 6.608574, 6.61134, 6.620117, 
    6.626167, 6.612196, 6.627687, 6.574109, 6.601316, 6.558817, 6.571572, 
    6.580483, 6.576594, 6.596881, 6.601666, 6.622725, 6.611075, 6.67293, 
    6.646187, 6.720757, 6.699817, 6.558967, 6.565445, 6.587999, 6.57727, 
    6.608048, 6.615639, 6.623421, 6.631325, 6.632193, 6.636885, 6.629196, 
    6.636589, 6.607083, 6.621125, 6.585441, 6.593712, 6.589911, 6.585732, 
    6.598638, 6.612387, 6.61271, 6.618703, 6.631105, 6.608173, 6.676331, 
    6.635073, 6.572515, 6.584974, 6.586788, 6.581955, 6.614877, 6.602925, 
    6.636775, 6.628039, 6.642367, 6.635241, 6.634192, 6.625059, 6.619373, 
    6.603467, 6.591845, 6.58266, 6.584796, 6.594891, 6.613235, 6.632258, 
    6.628428, 6.641278, 6.60581, 6.621556, 6.614483, 6.6304, 6.5975, 
    6.625647, 6.590718, 6.593641, 6.602688, 6.622499, 6.626585, 6.6309, 
    6.628244, 6.613707, 6.611603, 6.602475, 6.599943, 6.593007, 6.587257, 
    6.592503, 6.598011, 6.613726, 6.629498, 6.645024, 6.648841, 6.666961, 
    6.652164, 6.676555, 6.655746, 6.691844, 6.627234, 6.6552, 6.60311, 
    6.608534, 6.61991, 6.642516, 6.630333, 6.644598, 6.611523, 6.595225, 
    6.591051, 6.583212, 6.59123, 6.590579, 6.59826, 6.595792, 6.614248, 
    6.60433, 6.634156, 6.644493, 6.673812, 6.691833, 6.710282, 6.718425, 
    6.720909, 6.721945 ;

 EFLX_LH_TOT_R =
  6.523794, 6.540125, 6.536952, 6.550135, 6.542829, 6.551457, 6.527113, 
    6.540763, 6.532053, 6.525279, 6.575651, 6.550726, 6.601721, 6.585755, 
    6.627564, 6.599216, 6.632985, 6.626819, 6.645467, 6.640121, 6.663968, 
    6.647936, 6.676415, 6.660152, 6.662682, 6.647403, 6.555763, 6.572534, 
    6.554764, 6.557154, 6.556088, 6.54297, 6.536342, 6.522566, 6.52507, 
    6.535199, 6.55823, 6.550441, 6.570138, 6.569693, 6.591645, 6.581743, 
    6.620341, 6.608221, 6.640345, 6.632642, 6.639977, 6.637756, 6.640007, 
    6.628716, 6.633549, 6.623633, 6.583592, 6.59486, 6.561271, 6.541056, 
    6.527707, 6.51823, 6.519569, 6.522116, 6.535258, 6.547664, 6.5571, 
    6.563406, 6.569628, 6.58841, 6.598429, 6.622461, 6.618424, 6.625282, 
    6.631878, 6.642933, 6.641116, 6.645985, 6.625119, 6.63897, 6.614541, 
    6.622359, 6.571227, 6.552548, 6.544515, 6.537559, 6.520597, 6.5323, 
    6.527681, 6.538696, 6.545691, 6.542234, 6.563578, 6.555283, 6.599024, 
    6.580162, 6.631109, 6.619255, 6.633957, 6.626454, 6.639307, 6.627739, 
    6.647806, 6.652172, 6.649186, 6.6607, 6.627095, 6.639968, 6.542132, 
    6.542696, 6.545331, 6.533754, 6.533053, 6.522493, 6.531897, 6.535898, 
    6.546104, 6.552127, 6.557842, 6.57043, 6.584489, 6.604214, 6.620022, 
    6.62958, 6.623724, 6.628893, 6.623111, 6.620407, 6.650529, 6.633588, 
    6.659042, 6.657634, 6.646096, 6.657794, 6.543093, 6.53985, 6.528574, 
    6.537397, 6.521346, 6.530313, 6.535468, 6.555437, 6.559839, 6.563895, 
    6.571935, 6.58225, 6.600362, 6.617761, 6.632266, 6.631204, 6.631577, 
    6.634811, 6.626788, 6.636131, 6.63769, 6.633598, 6.657445, 6.650624, 
    6.657604, 6.653165, 6.540906, 6.546369, 6.543415, 6.548965, 6.545046, 
    6.562413, 6.567619, 6.592047, 6.582041, 6.598, 6.583668, 6.586199, 
    6.59848, 6.584448, 6.615288, 6.594326, 6.634938, 6.612304, 6.636257, 
    6.632203, 6.638927, 6.644943, 6.652539, 6.666549, 6.663306, 6.675056, 
    6.554515, 6.561577, 6.560972, 6.568383, 6.573865, 6.585772, 6.604887, 
    6.597697, 6.610922, 6.613573, 6.593496, 6.605799, 6.566321, 6.572671, 
    6.568903, 6.555061, 6.599329, 6.576578, 6.620254, 6.606301, 6.644083, 
    6.626027, 6.661517, 6.676698, 6.691111, 6.707887, 6.565454, 6.560649, 
    6.56927, 6.581177, 6.592283, 6.607052, 6.608574, 6.61134, 6.620117, 
    6.626167, 6.612196, 6.627687, 6.574109, 6.601316, 6.558817, 6.571572, 
    6.580483, 6.576594, 6.596881, 6.601666, 6.622725, 6.611075, 6.67293, 
    6.646187, 6.720757, 6.699817, 6.558967, 6.565445, 6.587999, 6.57727, 
    6.608048, 6.615639, 6.623421, 6.631325, 6.632193, 6.636885, 6.629196, 
    6.636589, 6.607083, 6.621125, 6.585441, 6.593712, 6.589911, 6.585732, 
    6.598638, 6.612387, 6.61271, 6.618703, 6.631105, 6.608173, 6.676331, 
    6.635073, 6.572515, 6.584974, 6.586788, 6.581955, 6.614877, 6.602925, 
    6.636775, 6.628039, 6.642367, 6.635241, 6.634192, 6.625059, 6.619373, 
    6.603467, 6.591845, 6.58266, 6.584796, 6.594891, 6.613235, 6.632258, 
    6.628428, 6.641278, 6.60581, 6.621556, 6.614483, 6.6304, 6.5975, 
    6.625647, 6.590718, 6.593641, 6.602688, 6.622499, 6.626585, 6.6309, 
    6.628244, 6.613707, 6.611603, 6.602475, 6.599943, 6.593007, 6.587257, 
    6.592503, 6.598011, 6.613726, 6.629498, 6.645024, 6.648841, 6.666961, 
    6.652164, 6.676555, 6.655746, 6.691844, 6.627234, 6.6552, 6.60311, 
    6.608534, 6.61991, 6.642516, 6.630333, 6.644598, 6.611523, 6.595225, 
    6.591051, 6.583212, 6.59123, 6.590579, 6.59826, 6.595792, 6.614248, 
    6.60433, 6.634156, 6.644493, 6.673812, 6.691833, 6.710282, 6.718425, 
    6.720909, 6.721945 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.356978e-08, 6.384934e-08, 6.379499e-08, 6.402048e-08, 6.389539e-08, 
    6.404304e-08, 6.362645e-08, 6.386044e-08, 6.371106e-08, 6.359494e-08, 
    6.445807e-08, 6.403054e-08, 6.490213e-08, 6.462948e-08, 6.531439e-08, 
    6.485971e-08, 6.540607e-08, 6.530126e-08, 6.561668e-08, 6.552632e-08, 
    6.592977e-08, 6.565838e-08, 6.61389e-08, 6.586495e-08, 6.590781e-08, 
    6.564943e-08, 6.411657e-08, 6.440485e-08, 6.409949e-08, 6.41406e-08, 
    6.412215e-08, 6.389798e-08, 6.378502e-08, 6.354841e-08, 6.359136e-08, 
    6.376514e-08, 6.415908e-08, 6.402535e-08, 6.436237e-08, 6.435476e-08, 
    6.472996e-08, 6.456079e-08, 6.51914e-08, 6.501217e-08, 6.553009e-08, 
    6.539984e-08, 6.552398e-08, 6.548633e-08, 6.552447e-08, 6.533344e-08, 
    6.541529e-08, 6.524719e-08, 6.459248e-08, 6.478489e-08, 6.421101e-08, 
    6.386593e-08, 6.363672e-08, 6.347406e-08, 6.349706e-08, 6.35409e-08, 
    6.376616e-08, 6.397794e-08, 6.413933e-08, 6.42473e-08, 6.435366e-08, 
    6.467567e-08, 6.484608e-08, 6.522765e-08, 6.515878e-08, 6.527544e-08, 
    6.538689e-08, 6.557399e-08, 6.55432e-08, 6.562563e-08, 6.527236e-08, 
    6.550714e-08, 6.511956e-08, 6.522556e-08, 6.438261e-08, 6.406143e-08, 
    6.392494e-08, 6.380544e-08, 6.351474e-08, 6.371549e-08, 6.363636e-08, 
    6.382462e-08, 6.394425e-08, 6.388508e-08, 6.425024e-08, 6.410828e-08, 
    6.485618e-08, 6.453404e-08, 6.537388e-08, 6.517291e-08, 6.542206e-08, 
    6.529492e-08, 6.551276e-08, 6.53167e-08, 6.565631e-08, 6.573026e-08, 
    6.567973e-08, 6.587384e-08, 6.530584e-08, 6.552398e-08, 6.388343e-08, 
    6.389308e-08, 6.393803e-08, 6.374042e-08, 6.372833e-08, 6.354723e-08, 
    6.370837e-08, 6.377699e-08, 6.395118e-08, 6.405422e-08, 6.415217e-08, 
    6.436752e-08, 6.460803e-08, 6.494434e-08, 6.518594e-08, 6.53479e-08, 
    6.524859e-08, 6.533626e-08, 6.523825e-08, 6.519231e-08, 6.570255e-08, 
    6.541605e-08, 6.584592e-08, 6.582213e-08, 6.562759e-08, 6.582481e-08, 
    6.389985e-08, 6.384432e-08, 6.365153e-08, 6.38024e-08, 6.352751e-08, 
    6.368138e-08, 6.376987e-08, 6.411125e-08, 6.418625e-08, 6.425581e-08, 
    6.439316e-08, 6.456945e-08, 6.487869e-08, 6.514775e-08, 6.539337e-08, 
    6.537537e-08, 6.538171e-08, 6.543657e-08, 6.530066e-08, 6.545889e-08, 
    6.548544e-08, 6.541601e-08, 6.581894e-08, 6.570383e-08, 6.582162e-08, 
    6.574668e-08, 6.386237e-08, 6.395581e-08, 6.390532e-08, 6.400027e-08, 
    6.393338e-08, 6.42308e-08, 6.431998e-08, 6.473723e-08, 6.456598e-08, 
    6.483852e-08, 6.459366e-08, 6.463705e-08, 6.484741e-08, 6.460689e-08, 
    6.513292e-08, 6.47763e-08, 6.543871e-08, 6.50826e-08, 6.546102e-08, 
    6.53923e-08, 6.550608e-08, 6.560798e-08, 6.573618e-08, 6.597273e-08, 
    6.591795e-08, 6.611577e-08, 6.40951e-08, 6.42163e-08, 6.420562e-08, 
    6.433245e-08, 6.442625e-08, 6.462955e-08, 6.49556e-08, 6.483299e-08, 
    6.505808e-08, 6.510327e-08, 6.476129e-08, 6.497127e-08, 6.42974e-08, 
    6.440629e-08, 6.434146e-08, 6.410467e-08, 6.486125e-08, 6.447298e-08, 
    6.518994e-08, 6.49796e-08, 6.559345e-08, 6.528818e-08, 6.58878e-08, 
    6.614415e-08, 6.638538e-08, 6.666732e-08, 6.428244e-08, 6.420009e-08, 
    6.434753e-08, 6.455154e-08, 6.47408e-08, 6.499243e-08, 6.501818e-08, 
    6.506531e-08, 6.518741e-08, 6.529008e-08, 6.508023e-08, 6.531582e-08, 
    6.443155e-08, 6.489495e-08, 6.416896e-08, 6.438758e-08, 6.453951e-08, 
    6.447286e-08, 6.481897e-08, 6.490055e-08, 6.523204e-08, 6.506068e-08, 
    6.608088e-08, 6.562952e-08, 6.688197e-08, 6.653197e-08, 6.417132e-08, 
    6.428215e-08, 6.466789e-08, 6.448436e-08, 6.500922e-08, 6.513842e-08, 
    6.524344e-08, 6.53777e-08, 6.539219e-08, 6.547174e-08, 6.534139e-08, 
    6.546659e-08, 6.499297e-08, 6.520462e-08, 6.46238e-08, 6.476517e-08, 
    6.470013e-08, 6.46288e-08, 6.484896e-08, 6.508353e-08, 6.508854e-08, 
    6.516375e-08, 6.537572e-08, 6.501136e-08, 6.613915e-08, 6.544267e-08, 
    6.440301e-08, 6.461651e-08, 6.464699e-08, 6.456429e-08, 6.512547e-08, 
    6.492213e-08, 6.54698e-08, 6.532179e-08, 6.55643e-08, 6.544379e-08, 
    6.542606e-08, 6.527128e-08, 6.517492e-08, 6.493146e-08, 6.473337e-08, 
    6.457628e-08, 6.461281e-08, 6.478536e-08, 6.509788e-08, 6.539351e-08, 
    6.532875e-08, 6.554587e-08, 6.497117e-08, 6.521216e-08, 6.511902e-08, 
    6.536187e-08, 6.482973e-08, 6.52829e-08, 6.471389e-08, 6.476378e-08, 
    6.49181e-08, 6.522851e-08, 6.529717e-08, 6.53705e-08, 6.532525e-08, 
    6.510581e-08, 6.506986e-08, 6.491435e-08, 6.487141e-08, 6.475292e-08, 
    6.465483e-08, 6.474446e-08, 6.483858e-08, 6.51059e-08, 6.53468e-08, 
    6.560944e-08, 6.567371e-08, 6.59806e-08, 6.573079e-08, 6.614304e-08, 
    6.579257e-08, 6.639924e-08, 6.530915e-08, 6.578225e-08, 6.492512e-08, 
    6.501746e-08, 6.518448e-08, 6.556754e-08, 6.536073e-08, 6.560259e-08, 
    6.506844e-08, 6.479132e-08, 6.471961e-08, 6.458583e-08, 6.472267e-08, 
    6.471154e-08, 6.484247e-08, 6.48004e-08, 6.511478e-08, 6.494591e-08, 
    6.542562e-08, 6.560068e-08, 6.609504e-08, 6.63981e-08, 6.670659e-08, 
    6.684278e-08, 6.688423e-08, 6.690156e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRSEB =
  -4.643258e-15, -9.367801e-15, -1.306504e-14, -5.39862e-16, -6.8848e-15, 
    -9.790279e-15, -7.297412e-15, -3.607906e-15, 1.209054e-15, -8.643101e-15, 
    -1.05012e-14, -1.580187e-14, -1.564697e-14, -9.126037e-15, -1.571044e-14, 
    -5.931534e-16, 1.596547e-15, -9.39685e-15, -2.014121e-14, -1.575292e-14, 
    -5.938803e-15, -5.264326e-15, -9.975355e-15, -5.478088e-15, 
    -1.684662e-14, -9.708356e-15, -9.615011e-15, -9.928033e-15, 
    -2.321841e-15, -6.850571e-15, -1.181895e-14, -9.430252e-15, 
    -1.049139e-14, -1.181165e-14, -4.14518e-15, -6.828756e-15, -4.768786e-15, 
    -6.413302e-15, -5.967873e-15, -6.544592e-15, -1.060856e-14, 
    -1.810425e-14, -1.004962e-14, -5.589013e-15, -8.338262e-15, -1.62676e-14, 
    -1.108147e-14, -1.060988e-14, -1.479528e-14, -8.931064e-15, 
    -1.333297e-14, -1.183362e-14, -1.133727e-14, -6.29335e-15, -1.82562e-14, 
    -1.205435e-14, -8.906852e-15, -7.638388e-15, -1.148976e-14, 
    -1.050009e-14, -4.893368e-15, -7.996775e-15, -3.809233e-15, 
    -7.451539e-15, -6.941775e-15, -4.109995e-15, -7.125787e-15, 
    -6.834199e-15, -8.169619e-15, -9.882036e-15, -1.657789e-14, 
    -5.026977e-15, -9.987054e-15, -1.07897e-14, -4.898056e-15, -1.435007e-14, 
    -1.251607e-15, -6.086202e-15, -1.879846e-15, -8.088449e-15, 
    -1.632774e-15, -2.584241e-15, -1.423219e-14, -1.112068e-14, 
    -8.494693e-15, -9.951566e-15, -4.854741e-15, -8.897402e-15, 6.011158e-16, 
    -7.336836e-15, -9.470081e-15, -1.328596e-14, -7.610667e-15, 
    -9.653956e-15, -2.441186e-14, -1.830398e-14, -1.050772e-14, 
    -1.237934e-14, -5.181783e-15, -1.007766e-14, -1.327154e-14, 
    -8.110437e-15, -7.226944e-15, -3.37185e-15, -1.128555e-14, -1.909283e-14, 
    -1.32679e-14, -1.422976e-14, -1.476654e-14, -1.644741e-14, -1.246719e-15, 
    -6.16099e-15, -1.826129e-15, -1.355221e-14, -1.068991e-14, -1.53046e-14, 
    -1.610203e-14, -1.433807e-14, -1.743637e-14, -1.136958e-14, 
    -3.381332e-15, -7.49435e-15, -6.942547e-15, -7.214324e-15, -1.422976e-14, 
    -4.301135e-15, -1.009108e-14, -6.362039e-15, -7.447435e-15, 3.068852e-15, 
    -1.331214e-14, -3.462345e-16, 5.574679e-15, -8.416589e-15, -2.307093e-14, 
    -1.275866e-15, -9.413001e-15, -7.17159e-15, -1.758063e-14, -1.322994e-14, 
    -4.993161e-15, -7.148476e-15, -1.277723e-14, -9.905775e-15, 
    -1.480422e-15, -7.682233e-15, -1.28246e-14, -1.403744e-14, 1.445524e-15, 
    -3.690917e-16, -9.07752e-15, -6.410959e-15, -1.019148e-14, 3.721751e-15, 
    -1.019523e-14, -1.032541e-14, -1.972116e-14, -3.54234e-16, -9.301947e-15, 
    -1.317802e-14, -1.182062e-14, -3.412248e-15, -1.064577e-14, 
    -3.289948e-15, -5.042475e-15, -9.880948e-15, -7.068398e-15, 
    -8.134152e-16, -2.765744e-15, -1.0733e-14, -1.097789e-14, -2.830213e-15, 
    -6.220889e-16, -5.416704e-15, -7.444385e-15, 7.82965e-16, -5.077498e-15, 
    -1.045739e-14, -8.643295e-15, -1.605808e-14, -1.210299e-14, 2.097406e-15, 
    -3.223969e-15, -1.109892e-14, -1.00434e-14, -1.669492e-14, 4.392409e-16, 
    -1.019399e-14, -1.168215e-14, 1.718506e-15, -1.577669e-14, -1.120727e-14, 
    -1.657573e-14, -3.157908e-15, -4.61886e-15, -9.403496e-15, -8.677892e-15, 
    -1.822277e-14, 2.598638e-15, -4.496613e-15, -1.218079e-14, -1.099392e-15, 
    -5.173263e-15, -1.617004e-14, -1.539868e-14, -1.206732e-14, 
    -1.260039e-14, -1.503798e-15, -3.150272e-15, -9.09167e-15, -6.190776e-15, 
    -1.267334e-15, -1.346029e-14, -1.027098e-14, -5.877122e-15, 
    -1.287222e-14, -1.001498e-14, -7.115044e-15, -6.619287e-15, 
    -1.123545e-14, -8.217566e-15, -1.50527e-14, -1.014829e-14, -6.885886e-17, 
    6.010935e-15, -4.14069e-15, -1.253889e-14, -1.147066e-14, -1.50038e-14, 
    -7.019027e-15, -7.143009e-15, -7.755201e-15, -1.094641e-14, 
    -7.583227e-15, -1.716818e-14, -9.792056e-15, -4.992074e-15, -1.28976e-14, 
    1.787789e-15, -8.36789e-15, 1.397624e-16, -8.341423e-15, -1.836751e-15, 
    -1.053711e-14, -8.337542e-15, -1.064758e-14, -8.492661e-15, 
    -6.308425e-15, -1.43104e-14, -9.730194e-15, -1.478474e-14, -9.163422e-15, 
    -8.458404e-15, -1.372751e-14, -7.300026e-15, -1.017004e-14, -4.55858e-15, 
    -5.444349e-15, -4.235462e-15, -8.563946e-15, -1.517483e-14, 
    -1.268553e-14, -4.947947e-15, -1.477747e-14, -5.99418e-15, -1.398433e-14, 
    -9.005255e-15, -1.329016e-14, 4.992677e-16, -8.098809e-15, 3.573859e-16, 
    -6.291194e-15, -1.573147e-14, -1.535686e-14, -8.193902e-15, -1.13033e-14, 
    -1.166382e-14, -7.463769e-15, -4.607307e-15, -5.396685e-15, 
    -1.082556e-14, -1.00714e-14, -8.57942e-15, -1.414407e-14, -1.429508e-14, 
    -8.147845e-15, -5.149469e-15, -9.931403e-15, -1.169968e-14, 
    -5.455674e-15, -6.557662e-15, -5.82905e-15, -1.177913e-14, -1.275052e-14, 
    4.455899e-16, -1.373441e-14, -6.141258e-15, -5.117297e-15, -1.662262e-14, 
    -7.847162e-15, -1.129397e-14, -5.364809e-15, -4.209966e-15, 
    -1.877304e-14, -1.198109e-14, -6.481075e-15, -5.119728e-15, 
    -8.121426e-15, -1.568192e-14, -4.452002e-15, -7.409073e-15, 
    -6.154919e-15, -6.580334e-15, -5.001218e-15, -9.647013e-15, 
    -1.039469e-14, -2.745359e-15, -9.111106e-15, -1.568762e-14, 
    -9.217701e-15, -1.032317e-14, -9.180882e-15, -1.417649e-14, 
    -7.255539e-15, -5.971398e-15, -4.903922e-15, -8.717683e-15, 
    -1.344532e-14, -1.307574e-14, -9.69786e-15, -8.620786e-15, -8.333576e-15, 
    -9.160559e-15, -5.796393e-15, -1.223654e-14, -5.413009e-15, 
    -2.168326e-15, -1.187231e-14 ;

 ERRSOI =
  -71.26398, -71.35706, -71.33938, -71.41357, -71.37308, -71.42117, 
    -71.28365, -71.36004, -71.31173, -71.27346, -71.5556, -71.41708, 
    -71.7077, -71.61771, -71.84664, -71.69258, -71.87809, -71.84405, 
    -71.95113, -71.92053, -72.05389, -71.96526, -72.12624, -72.0337, 
    -72.04746, -71.96204, -71.44669, -71.53773, -71.44088, -71.45395, 
    -71.4485, -71.37328, -71.33424, -71.25813, -71.27227, -71.32886, 
    -71.45987, -71.41656, -71.52937, -71.52687, -71.6516, -71.59527, 
    -71.80697, -71.74704, -71.92185, -71.87756, -71.91944, -71.90697, 
    -71.91961, -71.85477, -71.88244, -71.82603, -71.60547, -71.66956, 
    -71.47775, -71.36008, -71.28667, -71.23326, -71.2408, -71.25481, 
    -71.32915, -71.40075, -71.45483, -71.49078, -71.52647, -71.62996, 
    -71.68887, -71.81818, -71.79639, -71.83452, -71.87323, -71.93616, 
    -71.92603, -71.95341, -71.83466, -71.91297, -71.78352, -71.81876, 
    -71.52995, -71.42852, -71.38014, -71.34254, -71.24648, -71.31246, 
    -71.28629, -71.34989, -71.38945, -71.37013, -71.49178, -71.4442, 
    -71.69238, -71.58533, -71.86873, -71.80099, -71.8852, -71.84251, 
    -71.91516, -71.84979, -71.9641, -71.98832, -71.97163, -72.0379, -71.846, 
    -71.91885, -71.3693, -71.37241, -71.38764, -71.32062, -71.31688, 
    -71.25742, -71.31089, -71.33316, -71.39224, -71.42605, -71.45864, 
    -71.53048, -71.6098, -71.72284, -71.80531, -71.86036, -71.82701, 
    -71.8564, -71.8233, -71.80807, -71.97884, -71.88232, -72.02835, 
    -72.02047, -71.95381, -72.02138, -71.3747, -71.3566, -71.2918, -71.34252, 
    -71.25105, -71.30144, -71.32997, -71.44383, -71.47038, -71.49307, 
    -71.53938, -71.59812, -71.70099, -71.79183, -71.87575, -71.86972, 
    -71.87178, -71.8899, -71.84415, -71.89748, -71.90582, -71.88305, 
    -72.01938, -71.98046, -72.0203, -71.9951, -71.36264, -71.3934, -71.37667, 
    -71.40778, -71.38537, -71.48335, -71.51274, -71.65245, -71.5966, 
    -71.68723, -71.6063, -71.62027, -71.68755, -71.61108, -71.78551, 
    -71.6648, -71.89062, -71.76713, -71.89822, -71.87537, -71.91382, 
    -71.9476, -71.99129, -72.07024, -72.0522, -72.11933, -71.43987, 
    -71.47929, -71.47697, -71.5191, -71.55, -71.61855, -71.72737, -71.68678, 
    -71.76261, -71.77744, -71.66296, -71.73209, -71.50658, -71.54169, 
    -71.52165, -71.44229, -71.69452, -71.56414, -71.80646, -71.73573, 
    -71.94262, -71.83841, -72.04199, -72.12628, -72.2113, -72.30445, 
    -71.50209, -71.47516, -71.52444, -71.59056, -71.65535, -71.73981, 
    -71.74911, -71.7646, -71.80634, -71.84079, -71.76836, -71.84956, 
    -71.54749, -71.7064, -71.46389, -71.53518, -71.58718, -71.56554, 
    -71.68245, -71.70963, -71.81999, -71.76353, -72.10442, -71.95307, 
    -72.37952, -72.25906, -71.46546, -71.50255, -71.63016, -71.56957, 
    -71.74608, -71.78912, -71.82528, -71.86949, -71.87514, -71.90152, 
    -71.85816, -71.90026, -71.73998, -71.81176, -71.61695, -71.66356, 
    -71.64252, -71.61858, -71.69236, -71.7692, -71.77275, -71.7972, 
    -71.86252, -71.74683, -72.1205, -71.88602, -71.5429, -71.6119, -71.62407, 
    -71.59691, -71.78474, -71.71633, -71.90115, -71.85153, -71.93335, 
    -71.8925, -71.88641, -71.83447, -71.80166, -71.7191, -71.6527, -71.60108, 
    -71.61322, -71.66999, -71.77435, -71.8748, -71.85252, -71.92715, 
    -71.73318, -71.81346, -71.78172, -71.86472, -71.68528, -71.83231, 
    -71.64716, -71.66374, -71.71499, -71.81763, -71.84319, -71.86707, 
    -71.85273, -71.77735, -71.76589, -71.7142, -71.69901, -71.66028, 
    -71.62734, -71.65696, -71.68768, -71.77818, -71.85895, -71.9478, 
    -71.9703, -72.06968, -71.98614, -72.12142, -72.00241, -72.21064, 
    -71.84362, -72.00279, -71.71796, -71.74899, -71.80323, -71.93185, 
    -71.86435, -71.94421, -71.76559, -71.671, -71.64893, -71.60387, 
    -71.64996, -71.64629, -71.69031, -71.67627, -71.78121, -71.72488, 
    -71.88574, -71.94405, -72.1116, -72.21349, -72.32056, -72.36691, 
    -72.3812, -72.38706 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.621211, -1.620114, -1.620322, -1.619446, -1.619924, -1.619356, 
    -1.620979, -1.620079, -1.620648, -1.621099, -1.617766, -1.619404, 
    -1.615975, -1.617031, -1.614345, -1.616153, -1.613973, -1.614374, 
    -1.613107, -1.61347, -1.611889, -1.61294, -1.611027, -1.612128, 
    -1.611965, -1.612978, -1.619054, -1.617978, -1.619122, -1.618968, 
    -1.619032, -1.619922, -1.620384, -1.62128, -1.621113, -1.620447, 
    -1.618898, -1.61941, -1.618073, -1.618103, -1.616633, -1.617294, 
    -1.614812, -1.615511, -1.613454, -1.613978, -1.613483, -1.61363, 
    -1.613481, -1.614248, -1.613921, -1.614587, -1.617175, -1.616423, 
    -1.618686, -1.62008, -1.620944, -1.621572, -1.621484, -1.621319, 
    -1.620443, -1.619597, -1.618957, -1.618531, -1.618108, -1.61689, 
    -1.616196, -1.61468, -1.614936, -1.614487, -1.614029, -1.613285, 
    -1.613405, -1.613081, -1.614485, -1.61356, -1.615081, -1.614673, 
    -1.61807, -1.619268, -1.619842, -1.620285, -1.621417, -1.62064, 
    -1.620948, -1.620198, -1.619731, -1.619959, -1.618519, -1.619083, 
    -1.616155, -1.617412, -1.614083, -1.614882, -1.613888, -1.614392, 
    -1.613534, -1.614306, -1.612954, -1.612667, -1.612865, -1.612078, 
    -1.614351, -1.61349, -1.619969, -1.619932, -1.619752, -1.620544, 
    -1.620588, -1.621288, -1.620658, -1.620396, -1.619697, -1.619298, 
    -1.618912, -1.618061, -1.617124, -1.615796, -1.614831, -1.614181, 
    -1.614575, -1.614228, -1.614619, -1.614798, -1.61278, -1.613922, 
    -1.612191, -1.612285, -1.613076, -1.612274, -1.619905, -1.620118, 
    -1.620883, -1.620285, -1.621363, -1.62077, -1.620434, -1.619088, 
    -1.618773, -1.618504, -1.617955, -1.617261, -1.616053, -1.61499, 
    -1.613999, -1.614071, -1.614046, -1.613832, -1.614373, -1.613743, 
    -1.613644, -1.613913, -1.612298, -1.612759, -1.612287, -1.612586, 
    -1.620047, -1.619684, -1.619881, -1.619514, -1.619779, -1.61862, 
    -1.618272, -1.616624, -1.617279, -1.616215, -1.617165, -1.617001, 
    -1.616213, -1.617108, -1.615059, -1.61648, -1.613824, -1.615277, 
    -1.613734, -1.614004, -1.613549, -1.61315, -1.612631, -1.611694, 
    -1.611908, -1.611109, -1.619134, -1.618668, -1.618695, -1.618195, 
    -1.617829, -1.617021, -1.615742, -1.616219, -1.615327, -1.615153, 
    -1.616499, -1.615687, -1.618344, -1.617929, -1.618165, -1.619106, 
    -1.61613, -1.617662, -1.614818, -1.615644, -1.613209, -1.614442, 
    -1.612029, -1.611027, -1.61001, -1.608896, -1.618397, -1.618716, 
    -1.618132, -1.617351, -1.616589, -1.615596, -1.615486, -1.615304, 
    -1.614819, -1.614412, -1.615261, -1.614309, -1.617861, -1.615989, 
    -1.61885, -1.618006, -1.61739, -1.617644, -1.61627, -1.61595, -1.614659, 
    -1.615317, -1.611288, -1.613086, -1.607993, -1.60944, -1.618831, 
    -1.618392, -1.616885, -1.617597, -1.615522, -1.615016, -1.614595, 
    -1.614074, -1.614007, -1.613695, -1.614207, -1.61371, -1.615594, 
    -1.614755, -1.617039, -1.616493, -1.616739, -1.61702, -1.616154, 
    -1.615251, -1.615208, -1.614927, -1.61416, -1.615513, -1.611099, 
    -1.613882, -1.617913, -1.6171, -1.616956, -1.617275, -1.615067, 
    -1.615872, -1.613699, -1.614285, -1.613318, -1.613801, -1.613874, 
    -1.614487, -1.614874, -1.615839, -1.61662, -1.617226, -1.617083, 
    -1.616417, -1.61519, -1.614011, -1.614275, -1.613391, -1.615674, 
    -1.614735, -1.615103, -1.61413, -1.616237, -1.614516, -1.616685, 
    -1.61649, -1.615888, -1.614687, -1.614384, -1.614103, -1.614271, 
    -1.615155, -1.615289, -1.615897, -1.616076, -1.616531, -1.616917, 
    -1.61657, -1.616209, -1.615144, -1.614199, -1.613147, -1.61288, 
    -1.611702, -1.612694, -1.611088, -1.612504, -1.610021, -1.614381, 
    -1.612497, -1.615852, -1.615488, -1.614857, -1.613337, -1.614134, 
    -1.613191, -1.615293, -1.616406, -1.616664, -1.617193, -1.616652, 
    -1.616695, -1.616178, -1.616343, -1.615109, -1.615771, -1.613882, 
    -1.613192, -1.611201, -1.609985, -1.608701, -1.608145, -1.607973, 
    -1.607902 ;

 FCH4 =
  1.821471e-13, 1.820607e-13, 1.820786e-13, 1.82001e-13, 1.820453e-13, 
    1.819928e-13, 1.821307e-13, 1.820569e-13, 1.821052e-13, 1.8214e-13, 
    1.818218e-13, 1.819974e-13, 1.806104e-13, 1.805992e-13, 1.805664e-13, 
    1.806105e-13, 1.805461e-13, 1.805693e-13, 1.80484e-13, 1.805134e-13, 
    1.803494e-13, 1.80469e-13, 1.802309e-13, 1.803816e-13, 1.803606e-13, 
    1.804723e-13, 1.819653e-13, 1.818457e-13, 1.819718e-13, 1.819559e-13, 
    1.819631e-13, 1.820443e-13, 1.820815e-13, 1.821534e-13, 1.82141e-13, 
    1.820881e-13, 1.819487e-13, 1.819994e-13, 1.818651e-13, 1.818684e-13, 
    1.80607e-13, 1.805916e-13, 1.805878e-13, 1.806064e-13, 1.805123e-13, 
    1.805478e-13, 1.805141e-13, 1.805251e-13, 1.805139e-13, 1.805627e-13, 
    1.80544e-13, 1.805791e-13, 1.805953e-13, 1.806094e-13, 1.819282e-13, 
    1.820548e-13, 1.821276e-13, 1.82174e-13, 1.821676e-13, 1.821554e-13, 
    1.820877e-13, 1.820165e-13, 1.819566e-13, 1.819136e-13, 1.818689e-13, 
    1.806028e-13, 1.806106e-13, 1.805822e-13, 1.805923e-13, 1.80574e-13, 
    1.805509e-13, 1.804983e-13, 1.805082e-13, 1.804808e-13, 1.805747e-13, 
    1.80519e-13, 1.805971e-13, 1.805827e-13, 1.818555e-13, 1.819861e-13, 
    1.820347e-13, 1.820752e-13, 1.821627e-13, 1.821037e-13, 1.821277e-13, 
    1.82069e-13, 1.820284e-13, 1.820488e-13, 1.819124e-13, 1.819685e-13, 
    1.806106e-13, 1.80588e-13, 1.805539e-13, 1.805904e-13, 1.805423e-13, 
    1.805706e-13, 1.805174e-13, 1.805663e-13, 1.804697e-13, 1.80441e-13, 
    1.804609e-13, 1.803775e-13, 1.805684e-13, 1.80514e-13, 1.820494e-13, 
    1.820461e-13, 1.820306e-13, 1.820959e-13, 1.820997e-13, 1.821536e-13, 
    1.82106e-13, 1.820843e-13, 1.82026e-13, 1.819888e-13, 1.819515e-13, 
    1.818628e-13, 1.805969e-13, 1.806095e-13, 1.805886e-13, 1.805597e-13, 
    1.80579e-13, 1.805622e-13, 1.805807e-13, 1.805878e-13, 1.804521e-13, 
    1.805437e-13, 1.803907e-13, 1.804017e-13, 1.8048e-13, 1.804004e-13, 
    1.820438e-13, 1.820625e-13, 1.821233e-13, 1.820763e-13, 1.821592e-13, 
    1.821142e-13, 1.820865e-13, 1.819672e-13, 1.819382e-13, 1.8191e-13, 
    1.818516e-13, 1.805926e-13, 1.806107e-13, 1.805936e-13, 1.805494e-13, 
    1.805536e-13, 1.805521e-13, 1.805386e-13, 1.805694e-13, 1.805327e-13, 
    1.805253e-13, 1.805438e-13, 1.804031e-13, 1.804517e-13, 1.804019e-13, 
    1.804344e-13, 1.820565e-13, 1.820244e-13, 1.820419e-13, 1.820085e-13, 
    1.820321e-13, 1.819201e-13, 1.81883e-13, 1.806072e-13, 1.805922e-13, 
    1.806106e-13, 1.805955e-13, 1.805999e-13, 1.806103e-13, 1.80597e-13, 
    1.805952e-13, 1.806089e-13, 1.80538e-13, 1.806004e-13, 1.805321e-13, 
    1.805497e-13, 1.805195e-13, 1.804869e-13, 1.804387e-13, 1.803272e-13, 
    1.803557e-13, 1.802453e-13, 1.819735e-13, 1.81926e-13, 1.819305e-13, 
    1.81878e-13, 1.818369e-13, 1.805993e-13, 1.806091e-13, 1.806107e-13, 
    1.80603e-13, 1.805987e-13, 1.806086e-13, 1.806084e-13, 1.818927e-13, 
    1.818455e-13, 1.81874e-13, 1.819698e-13, 1.806107e-13, 1.818155e-13, 
    1.80588e-13, 1.806081e-13, 1.804919e-13, 1.805716e-13, 1.803706e-13, 
    1.802274e-13, 1.800597e-13, 1.798201e-13, 1.81899e-13, 1.819327e-13, 
    1.818715e-13, 1.805902e-13, 1.806076e-13, 1.806074e-13, 1.80606e-13, 
    1.806023e-13, 1.805885e-13, 1.805715e-13, 1.806008e-13, 1.805664e-13, 
    1.818339e-13, 1.806106e-13, 1.819449e-13, 1.818538e-13, 1.805887e-13, 
    1.818158e-13, 1.806105e-13, 1.806107e-13, 1.805815e-13, 1.806028e-13, 
    1.802659e-13, 1.804792e-13, 1.796059e-13, 1.79941e-13, 1.819441e-13, 
    1.818992e-13, 1.806026e-13, 1.818105e-13, 1.806065e-13, 1.805948e-13, 
    1.805798e-13, 1.80553e-13, 1.805497e-13, 1.805291e-13, 1.805611e-13, 
    1.805306e-13, 1.806074e-13, 1.805859e-13, 1.805987e-13, 1.806087e-13, 
    1.806052e-13, 1.805992e-13, 1.806109e-13, 1.806005e-13, 1.806003e-13, 
    1.805916e-13, 1.805526e-13, 1.806064e-13, 1.8023e-13, 1.805363e-13, 
    1.818473e-13, 1.805977e-13, 1.806009e-13, 1.805921e-13, 1.805963e-13, 
    1.806102e-13, 1.805297e-13, 1.805652e-13, 1.805015e-13, 1.805367e-13, 
    1.805413e-13, 1.805749e-13, 1.805902e-13, 1.806099e-13, 1.806071e-13, 
    1.805936e-13, 1.805976e-13, 1.806094e-13, 1.805991e-13, 1.805492e-13, 
    1.805636e-13, 1.805074e-13, 1.806086e-13, 1.805847e-13, 1.805969e-13, 
    1.805566e-13, 1.806106e-13, 1.805721e-13, 1.806061e-13, 1.806087e-13, 
    1.806103e-13, 1.805819e-13, 1.805701e-13, 1.805546e-13, 1.805645e-13, 
    1.805984e-13, 1.806019e-13, 1.806105e-13, 1.806108e-13, 1.806083e-13, 
    1.806017e-13, 1.806078e-13, 1.806107e-13, 1.805985e-13, 1.805598e-13, 
    1.804864e-13, 1.804633e-13, 1.803226e-13, 1.804405e-13, 1.802276e-13, 
    1.804139e-13, 1.800485e-13, 1.805673e-13, 1.804189e-13, 1.806102e-13, 
    1.80606e-13, 1.805886e-13, 1.805002e-13, 1.805569e-13, 1.804886e-13, 
    1.806021e-13, 1.806095e-13, 1.806065e-13, 1.805946e-13, 1.806066e-13, 
    1.80606e-13, 1.806109e-13, 1.806101e-13, 1.805975e-13, 1.806096e-13, 
    1.805413e-13, 1.804893e-13, 1.802578e-13, 1.800497e-13, 1.797833e-13, 
    1.796472e-13, 1.796036e-13, 1.79585e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  8.145005, 8.160238, 8.157275, 8.16958, 8.162753, 8.170814, 8.148092, 
    8.160842, 8.152701, 8.146379, 8.193417, 8.170131, 8.217695, 8.202786, 
    8.241909, 8.215369, 8.246958, 8.241193, 8.258574, 8.253591, 8.275857, 
    8.260876, 8.287442, 8.27228, 8.274648, 8.260381, 8.174816, 8.190512, 
    8.173886, 8.176123, 8.17512, 8.162892, 8.156726, 8.143846, 8.146183, 
    8.155646, 8.177128, 8.169851, 8.18821, 8.187796, 8.208279, 8.199038, 
    8.235152, 8.223732, 8.253799, 8.24662, 8.25346, 8.251387, 8.253488, 
    8.242963, 8.24747, 8.23822, 8.200767, 8.211283, 8.179957, 8.161136, 
    8.14865, 8.139802, 8.141052, 8.143435, 8.155701, 8.167261, 8.176057, 
    8.181937, 8.187736, 8.2053, 8.214625, 8.237142, 8.23336, 8.23977, 
    8.245907, 8.256218, 8.25452, 8.259066, 8.239604, 8.25253, 8.229622, 
    8.237031, 8.189297, 8.171817, 8.164357, 8.157844, 8.142014, 8.152941, 
    8.14863, 8.158894, 8.165421, 8.162192, 8.182097, 8.174366, 8.215179, 
    8.197574, 8.245192, 8.234138, 8.247845, 8.240847, 8.25284, 8.242044, 
    8.260759, 8.264839, 8.262051, 8.272778, 8.241446, 8.253458, 8.162101, 
    8.162627, 8.165083, 8.154298, 8.153641, 8.143781, 8.152555, 8.156293, 
    8.165801, 8.171425, 8.176754, 8.18849, 8.201613, 8.220011, 8.234853, 
    8.243762, 8.238298, 8.243121, 8.23773, 8.235206, 8.263309, 8.24751, 
    8.271233, 8.269918, 8.259172, 8.270067, 8.162997, 8.159968, 8.149457, 
    8.157681, 8.142709, 8.151083, 8.155902, 8.174524, 8.178612, 8.182399, 
    8.18989, 8.199511, 8.216415, 8.232752, 8.246265, 8.245275, 8.245624, 
    8.248644, 8.24116, 8.249873, 8.251334, 8.247511, 8.269743, 8.263384, 
    8.269891, 8.26575, 8.160954, 8.166053, 8.163296, 8.168479, 8.164825, 
    8.181033, 8.185891, 8.208672, 8.19932, 8.214215, 8.200832, 8.2032, 
    8.214693, 8.201556, 8.230347, 8.210805, 8.248762, 8.22758, 8.249991, 
    8.246207, 8.252476, 8.258093, 8.26517, 8.278242, 8.275213, 8.286165, 
    8.173649, 8.180245, 8.179667, 8.186579, 8.191694, 8.202793, 8.22063, 
    8.213917, 8.226249, 8.228726, 8.209995, 8.221486, 8.184665, 8.190599, 
    8.187068, 8.174168, 8.215459, 8.19424, 8.235072, 8.221946, 8.257291, 
    8.240468, 8.273546, 8.287724, 8.301121, 8.316783, 8.183851, 8.179365, 
    8.187402, 8.198528, 8.208872, 8.222648, 8.224061, 8.226645, 8.234936, 
    8.24058, 8.227457, 8.241997, 8.19197, 8.217306, 8.177668, 8.189579, 
    8.197873, 8.194238, 8.213151, 8.217616, 8.237384, 8.226392, 8.284219, 
    8.259273, 8.328751, 8.309258, 8.177798, 8.183837, 8.204885, 8.194866, 
    8.223571, 8.230655, 8.238016, 8.245399, 8.2462, 8.25058, 8.243403, 
    8.250299, 8.222677, 8.23588, 8.20248, 8.210205, 8.206651, 8.202753, 
    8.214792, 8.227638, 8.227919, 8.233631, 8.245265, 8.223686, 8.28743, 
    8.248955, 8.190428, 8.202074, 8.203745, 8.19923, 8.229944, 8.218797, 
    8.250475, 8.242324, 8.255685, 8.249042, 8.248065, 8.239546, 8.234247, 
    8.219306, 8.208465, 8.199885, 8.20188, 8.211308, 8.228426, 8.24627, 
    8.242702, 8.254669, 8.221484, 8.236291, 8.229587, 8.24453, 8.213737, 
    8.240163, 8.207403, 8.210131, 8.218575, 8.237185, 8.24097, 8.245003, 
    8.242516, 8.228862, 8.226892, 8.218372, 8.216019, 8.209538, 8.204175, 
    8.209073, 8.21422, 8.22887, 8.243697, 8.258172, 8.261721, 8.278664, 
    8.264857, 8.287642, 8.26825, 8.301865, 8.241614, 8.267697, 8.218963, 
    8.224022, 8.234766, 8.255854, 8.244467, 8.257789, 8.226816, 8.211631, 
    8.207715, 8.200405, 8.207883, 8.207274, 8.214437, 8.212135, 8.229357, 
    8.2201, 8.248038, 8.257685, 8.285013, 8.301818, 8.318983, 8.32657, 
    8.328881, 8.329847 ;

 FGR =
  -324.1767, -324.9395, -324.7916, -325.4059, -325.0658, -325.4676, 
    -324.3321, -324.969, -324.5629, -324.2465, -326.5954, -325.4335, 
    -327.8078, -327.067, -328.9406, -327.6914, -329.1908, -328.9067, 
    -329.7664, -329.5202, -330.6161, -329.88, -331.1873, -330.4413, 
    -330.5573, -329.8555, -325.6691, -326.4501, -325.6224, -325.7339, 
    -325.6842, -325.0722, -324.7625, -324.1197, -324.2367, -324.7095, 
    -325.784, -325.4206, -326.3401, -326.3194, -327.3407, -326.8805, 
    -328.6074, -328.1097, -329.5305, -329.1754, -329.5135, -329.4112, 
    -329.5148, -328.9942, -329.2172, -328.7596, -326.9664, -327.4898, 
    -325.9262, -324.9822, -324.3597, -323.9167, -323.9793, -324.0984, 
    -324.7123, -325.2912, -325.7317, -326.0261, -326.3163, -327.1895, 
    -327.6552, -328.7052, -328.519, -328.8355, -329.1402, -329.6496, 
    -329.5659, -329.79, -328.8283, -329.4669, -328.4024, -328.7007, 
    -326.3891, -325.5189, -325.1436, -324.8198, -324.0273, -324.5742, 
    -324.3585, -324.8731, -325.1992, -325.0381, -326.0341, -325.6467, 
    -327.6828, -326.8066, -329.1046, -328.5573, -329.2361, -328.89, 
    -329.4825, -328.9493, -329.8739, -330.0746, -329.9373, -330.4667, 
    -328.9196, -329.5129, -325.0334, -325.0596, -325.1825, -324.6421, 
    -324.6094, -324.1161, -324.5556, -324.7422, -325.2186, -325.4992, 
    -325.7662, -326.3535, -327.0079, -327.9237, -328.5927, -329.0343, 
    -328.7639, -329.0025, -328.7356, -328.6107, -329.999, -329.2189, 
    -330.3905, -330.3259, -329.7951, -330.3332, -325.0781, -324.927, 
    -324.4003, -324.8125, -324.0625, -324.4815, -324.722, -325.6535, 
    -325.8596, -326.0487, -326.4238, -326.904, -327.7451, -328.4881, 
    -329.1582, -329.1092, -329.1264, -329.2754, -328.9053, -329.3362, 
    -329.408, -329.2195, -330.3172, -330.0037, -330.3245, -330.1205, 
    -324.9763, -325.2308, -325.0932, -325.3517, -325.1691, -325.9792, 
    -326.222, -327.3589, -326.8942, -327.6355, -326.97, -327.0876, -327.6571, 
    -327.0064, -328.4363, -327.4646, -329.2812, -328.2979, -329.3421, 
    -329.1552, -329.4652, -329.7421, -330.0917, -330.735, -330.5862, 
    -331.1252, -325.6109, -325.9404, -325.9125, -326.2582, -326.5136, 
    -327.0679, -327.9551, -327.6218, -328.2348, -328.3575, -327.4268, 
    -327.9972, -326.1618, -326.4575, -326.2823, -325.6362, -327.6971, 
    -326.6396, -328.6034, -328.0207, -329.7025, -328.8698, -330.5041, 
    -331.1999, -331.8602, -332.6257, -326.1215, -325.8975, -326.2997, 
    -326.8537, -327.3703, -328.0554, -328.1261, -328.2541, -328.5973, 
    -328.8767, -328.2934, -328.9469, -326.5237, -327.7894, -325.8117, 
    -326.4062, -326.8216, -326.6407, -327.584, -327.8059, -328.7174, 
    -328.2419, -331.0272, -329.799, -333.2124, -332.2576, -325.8189, 
    -326.1213, -327.1711, -326.6722, -328.1017, -328.453, -328.7499, 
    -329.1145, -329.1548, -329.3709, -329.0165, -329.3574, -328.0568, 
    -328.6438, -327.0526, -327.4367, -327.2604, -327.0662, -327.6655, 
    -328.3022, -328.3176, -328.5317, -329.1029, -328.1075, -331.1823, 
    -329.2862, -326.4509, -327.0302, -327.1151, -326.8905, -328.4177, 
    -327.8642, -329.3659, -328.9631, -329.6236, -329.2952, -329.2469, 
    -328.8255, -328.5628, -327.8892, -327.3499, -326.9233, -327.0227, 
    -327.4914, -328.3415, -329.1576, -328.9808, -329.5735, -327.998, 
    -328.6635, -328.3993, -329.072, -327.6125, -328.8512, -327.2979, 
    -327.4336, -327.8532, -328.7067, -328.896, -329.0949, -328.9726, 
    -328.3634, -328.2662, -327.8434, -327.7258, -327.4042, -327.1371, 
    -327.3807, -327.6361, -328.3645, -329.0302, -329.7458, -329.9216, 
    -330.7532, -330.0737, -331.1924, -330.2374, -331.8927, -328.9251, 
    -330.2131, -327.8729, -328.1243, -328.5872, -329.6299, -329.0689, 
    -329.7259, -328.2625, -327.5066, -327.3133, -326.9489, -327.3217, 
    -327.2914, -327.648, -327.5335, -328.3887, -327.9294, -329.2451, 
    -329.7212, -331.0681, -331.8928, -332.7354, -333.1064, -333.2195, 
    -333.2667 ;

 FGR12 =
  -224.4644, -224.4258, -224.4332, -224.4026, -224.4193, -224.3996, 
    -224.4563, -224.4246, -224.4446, -224.4605, -224.3451, -224.4013, 
    -224.2853, -224.3206, -224.2326, -224.2912, -224.2207, -224.2337, 
    -224.1933, -224.2047, -224.1552, -224.188, -224.1288, -224.1627, 
    -224.1576, -224.1892, -224.3893, -224.3523, -224.3916, -224.3863, 
    -224.3885, -224.4192, -224.4352, -224.4669, -224.461, -224.4375, 
    -224.3839, -224.4015, -224.3557, -224.3568, -224.3072, -224.3295, 
    -224.2478, -224.2701, -224.2042, -224.221, -224.2052, -224.2099, 
    -224.2051, -224.2296, -224.2191, -224.2405, -224.3254, -224.3001, 
    -224.3766, -224.4246, -224.455, -224.4773, -224.4741, -224.4683, 
    -224.4373, -224.4079, -224.3859, -224.3713, -224.3569, -224.3157, 
    -224.2926, -224.2435, -224.2519, -224.2373, -224.2226, -224.1989, 
    -224.2027, -224.1924, -224.2373, -224.2076, -224.256, -224.2433, 
    -224.3554, -224.3966, -224.4163, -224.4318, -224.4718, -224.4442, 
    -224.4551, -224.4288, -224.4126, -224.4205, -224.3709, -224.3903, 
    -224.2912, -224.3334, -224.2243, -224.2501, -224.218, -224.2343, 
    -224.2068, -224.2315, -224.1884, -224.1794, -224.1857, -224.1611, 
    -224.2329, -224.2054, -224.4208, -224.4195, -224.4133, -224.4409, 
    -224.4424, -224.4672, -224.4449, -224.4357, -224.4114, -224.3976, 
    -224.3844, -224.3553, -224.3237, -224.2794, -224.2484, -224.2274, 
    -224.2402, -224.229, -224.2416, -224.2474, -224.183, -224.2192, 
    -224.1646, -224.1675, -224.1923, -224.1672, -224.4186, -224.4261, 
    -224.4529, -224.4318, -224.4699, -224.4488, -224.437, -224.3904, 
    -224.3797, -224.3703, -224.3517, -224.3283, -224.2879, -224.2536, 
    -224.2216, -224.2239, -224.2231, -224.2163, -224.2336, -224.2134, 
    -224.2103, -224.2189, -224.1679, -224.1824, -224.1676, -224.1769, 
    -224.4236, -224.4109, -224.4178, -224.4051, -224.4142, -224.3743, 
    -224.3624, -224.3069, -224.3289, -224.2933, -224.3251, -224.3195, 
    -224.2931, -224.3232, -224.2552, -224.3021, -224.216, -224.2623, 
    -224.2132, -224.2218, -224.2073, -224.1946, -224.1783, -224.1492, 
    -224.1559, -224.1313, -224.392, -224.376, -224.377, -224.3598, -224.3475, 
    -224.3202, -224.2776, -224.2935, -224.264, -224.2583, -224.3028, 
    -224.2758, -224.3649, -224.3508, -224.3588, -224.3911, -224.2904, 
    -224.3418, -224.248, -224.2744, -224.1965, -224.2358, -224.1596, 
    -224.1288, -224.0981, -224.0651, -224.3667, -224.3777, -224.3577, 
    -224.3313, -224.3058, -224.2728, -224.2693, -224.2633, -224.248, 
    -224.2349, -224.2618, -224.2315, -224.3485, -224.2858, -224.3823, 
    -224.3533, -224.3327, -224.3412, -224.2952, -224.2845, -224.2428, 
    -224.2637, -224.1368, -224.1926, -224.0387, -224.0811, -224.3817, 
    -224.3665, -224.3156, -224.3397, -224.2704, -224.2538, -224.2408, 
    -224.224, -224.2219, -224.2119, -224.2283, -224.2124, -224.2728, 
    -224.246, -224.3209, -224.3025, -224.3108, -224.3202, -224.2913, 
    -224.2615, -224.2601, -224.2515, -224.2267, -224.2702, -224.131, 
    -224.2179, -224.3503, -224.3228, -224.3181, -224.3288, -224.2555, 
    -224.282, -224.212, -224.2308, -224.1999, -224.2153, -224.2176, 
    -224.2373, -224.2498, -224.2809, -224.3068, -224.3272, -224.3224, -224.3, 
    -224.2595, -224.222, -224.2305, -224.2022, -224.2755, -224.2453, 
    -224.2567, -224.2258, -224.2941, -224.2381, -224.309, -224.3025, 
    -224.2825, -224.2437, -224.234, -224.2249, -224.2303, -224.2584, 
    -224.2628, -224.2828, -224.2887, -224.3038, -224.3168, -224.3051, 
    -224.2931, -224.258, -224.228, -224.1945, -224.1862, -224.1495, 
    -224.1803, -224.1307, -224.1744, -224.0984, -224.2339, -224.1741, 
    -224.2813, -224.2693, -224.2493, -224.2005, -224.226, -224.1959, 
    -224.2629, -224.2996, -224.3083, -224.3261, -224.3079, -224.3093, 
    -224.2921, -224.2976, -224.2569, -224.2786, -224.2179, -224.196, 
    -224.1341, -224.0974, -224.0593, -224.0431, -224.0381, -224.0361 ;

 FGR_R =
  -324.1767, -324.9395, -324.7916, -325.4059, -325.0658, -325.4676, 
    -324.3321, -324.969, -324.5629, -324.2465, -326.5954, -325.4335, 
    -327.8078, -327.067, -328.9406, -327.6914, -329.1908, -328.9067, 
    -329.7664, -329.5202, -330.6161, -329.88, -331.1873, -330.4413, 
    -330.5573, -329.8555, -325.6691, -326.4501, -325.6224, -325.7339, 
    -325.6842, -325.0722, -324.7625, -324.1197, -324.2367, -324.7095, 
    -325.784, -325.4206, -326.3401, -326.3194, -327.3407, -326.8805, 
    -328.6074, -328.1097, -329.5305, -329.1754, -329.5135, -329.4112, 
    -329.5148, -328.9942, -329.2172, -328.7596, -326.9664, -327.4898, 
    -325.9262, -324.9822, -324.3597, -323.9167, -323.9793, -324.0984, 
    -324.7123, -325.2912, -325.7317, -326.0261, -326.3163, -327.1895, 
    -327.6552, -328.7052, -328.519, -328.8355, -329.1402, -329.6496, 
    -329.5659, -329.79, -328.8283, -329.4669, -328.4024, -328.7007, 
    -326.3891, -325.5189, -325.1436, -324.8198, -324.0273, -324.5742, 
    -324.3585, -324.8731, -325.1992, -325.0381, -326.0341, -325.6467, 
    -327.6828, -326.8066, -329.1046, -328.5573, -329.2361, -328.89, 
    -329.4825, -328.9493, -329.8739, -330.0746, -329.9373, -330.4667, 
    -328.9196, -329.5129, -325.0334, -325.0596, -325.1825, -324.6421, 
    -324.6094, -324.1161, -324.5556, -324.7422, -325.2186, -325.4992, 
    -325.7662, -326.3535, -327.0079, -327.9237, -328.5927, -329.0343, 
    -328.7639, -329.0025, -328.7356, -328.6107, -329.999, -329.2189, 
    -330.3905, -330.3259, -329.7951, -330.3332, -325.0781, -324.927, 
    -324.4003, -324.8125, -324.0625, -324.4815, -324.722, -325.6535, 
    -325.8596, -326.0487, -326.4238, -326.904, -327.7451, -328.4881, 
    -329.1582, -329.1092, -329.1264, -329.2754, -328.9053, -329.3362, 
    -329.408, -329.2195, -330.3172, -330.0037, -330.3245, -330.1205, 
    -324.9763, -325.2308, -325.0932, -325.3517, -325.1691, -325.9792, 
    -326.222, -327.3589, -326.8942, -327.6355, -326.97, -327.0876, -327.6571, 
    -327.0064, -328.4363, -327.4646, -329.2812, -328.2979, -329.3421, 
    -329.1552, -329.4652, -329.7421, -330.0917, -330.735, -330.5862, 
    -331.1252, -325.6109, -325.9404, -325.9125, -326.2582, -326.5136, 
    -327.0679, -327.9551, -327.6218, -328.2348, -328.3575, -327.4268, 
    -327.9972, -326.1618, -326.4575, -326.2823, -325.6362, -327.6971, 
    -326.6396, -328.6034, -328.0207, -329.7025, -328.8698, -330.5041, 
    -331.1999, -331.8602, -332.6257, -326.1215, -325.8975, -326.2997, 
    -326.8537, -327.3703, -328.0554, -328.1261, -328.2541, -328.5973, 
    -328.8767, -328.2934, -328.9469, -326.5237, -327.7894, -325.8117, 
    -326.4062, -326.8216, -326.6407, -327.584, -327.8059, -328.7174, 
    -328.2419, -331.0272, -329.799, -333.2124, -332.2576, -325.8189, 
    -326.1213, -327.1711, -326.6722, -328.1017, -328.453, -328.7499, 
    -329.1145, -329.1548, -329.3709, -329.0165, -329.3574, -328.0568, 
    -328.6438, -327.0526, -327.4367, -327.2604, -327.0662, -327.6655, 
    -328.3022, -328.3176, -328.5317, -329.1029, -328.1075, -331.1823, 
    -329.2862, -326.4509, -327.0302, -327.1151, -326.8905, -328.4177, 
    -327.8642, -329.3659, -328.9631, -329.6236, -329.2952, -329.2469, 
    -328.8255, -328.5628, -327.8892, -327.3499, -326.9233, -327.0227, 
    -327.4914, -328.3415, -329.1576, -328.9808, -329.5735, -327.998, 
    -328.6635, -328.3993, -329.072, -327.6125, -328.8512, -327.2979, 
    -327.4336, -327.8532, -328.7067, -328.896, -329.0949, -328.9726, 
    -328.3634, -328.2662, -327.8434, -327.7258, -327.4042, -327.1371, 
    -327.3807, -327.6361, -328.3645, -329.0302, -329.7458, -329.9216, 
    -330.7532, -330.0737, -331.1924, -330.2374, -331.8927, -328.9251, 
    -330.2131, -327.8729, -328.1243, -328.5872, -329.6299, -329.0689, 
    -329.7259, -328.2625, -327.5066, -327.3133, -326.9489, -327.3217, 
    -327.2914, -327.648, -327.5335, -328.3887, -327.9294, -329.2451, 
    -329.7212, -331.0681, -331.8928, -332.7354, -333.1064, -333.2195, 
    -333.2667 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  74.74778, 74.80091, 74.79061, 74.83339, 74.80971, 74.83768, 74.75861, 
    74.80296, 74.77468, 74.75264, 74.9163, 74.83531, 75.00118, 74.9493, 
    75.07941, 74.99303, 75.09693, 75.07703, 75.13724, 75.12, 75.19672, 
    75.1452, 75.2367, 75.18449, 75.1926, 75.14348, 74.85173, 74.90617, 
    74.84848, 74.85625, 74.85279, 74.81015, 74.78858, 74.7438, 74.75196, 
    74.7849, 74.85974, 74.83441, 74.89851, 74.89707, 74.96848, 74.93624, 
    75.05608, 75.02235, 75.12072, 75.09586, 75.11953, 75.11237, 75.11962, 
    75.08316, 75.09878, 75.06673, 74.94225, 74.97892, 74.86966, 74.80388, 
    74.76054, 74.72967, 74.73403, 74.74232, 74.78509, 74.8254, 74.8561, 
    74.87663, 74.89686, 74.95787, 74.99049, 75.06291, 75.04988, 75.07205, 
    75.09338, 75.12906, 75.12321, 75.13889, 75.07155, 75.11626, 75.04286, 
    75.06261, 74.90192, 74.84126, 74.81512, 74.79257, 74.73738, 74.77547, 
    74.76044, 74.79629, 74.81899, 74.80779, 74.87718, 74.85017, 74.99243, 
    74.93108, 75.0909, 75.05257, 75.10011, 75.07587, 75.11736, 75.08002, 
    75.14477, 75.15881, 75.14921, 75.18626, 75.07793, 75.11949, 74.80745, 
    74.80927, 74.81783, 74.7802, 74.77792, 74.74356, 74.77418, 74.78718, 
    74.82035, 74.83989, 74.85851, 74.89945, 74.94515, 75.0093, 75.05505, 
    75.08597, 75.06704, 75.08375, 75.06505, 75.0563, 75.15352, 75.09889, 
    75.18093, 75.17641, 75.13924, 75.17693, 74.81056, 74.80004, 74.76336, 
    74.79207, 74.73983, 74.76901, 74.78576, 74.85065, 74.86501, 74.8782, 
    74.90435, 74.93789, 74.9968, 75.04771, 75.09465, 75.09122, 75.09242, 
    75.10286, 75.07694, 75.10712, 75.11214, 75.09895, 75.1758, 75.15385, 
    75.17632, 75.16203, 74.80347, 74.8212, 74.81161, 74.82961, 74.81689, 
    74.87335, 74.89027, 74.96974, 74.9372, 74.98912, 74.94251, 74.95074, 
    74.99062, 74.94506, 75.04523, 74.97714, 75.10326, 75.03552, 75.10753, 
    75.09444, 75.11615, 75.13554, 75.16001, 75.20504, 75.19463, 75.23236, 
    74.84767, 74.87065, 74.86871, 74.89281, 74.91061, 74.94937, 75.01151, 
    74.98817, 75.03111, 75.03971, 74.97451, 75.01446, 74.88609, 74.90669, 
    74.89449, 74.84944, 74.99343, 74.91939, 75.05579, 75.01611, 75.13276, 
    75.07445, 75.18888, 75.23758, 75.2838, 75.33734, 74.88328, 74.86766, 
    74.8957, 74.93436, 74.97055, 75.01854, 75.0235, 75.03246, 75.05537, 
    75.07494, 75.03522, 75.07986, 74.91131, 74.99989, 74.86167, 74.90312, 
    74.93212, 74.91946, 74.98552, 75.00106, 75.06377, 75.03162, 75.22549, 
    75.13951, 75.3784, 75.31159, 74.86218, 74.88326, 74.9566, 74.92167, 
    75.02179, 75.0464, 75.06606, 75.09159, 75.09441, 75.10955, 75.08473, 
    75.1086, 75.01864, 75.05862, 74.9483, 74.9752, 74.96285, 74.94925, 
    74.99123, 75.03583, 75.03692, 75.05077, 75.09075, 75.02219, 75.23633, 
    75.10359, 74.90623, 74.94672, 74.95267, 74.93694, 75.04393, 75.00513, 
    75.1092, 75.08099, 75.12724, 75.10425, 75.10086, 75.07135, 75.05295, 
    75.00689, 74.96912, 74.93924, 74.9462, 74.97903, 75.03859, 75.0946, 
    75.08222, 75.12373, 75.01452, 75.06, 75.04264, 75.08862, 74.98752, 
    75.07313, 74.96548, 74.97498, 75.00437, 75.06302, 75.07629, 75.09022, 
    75.08165, 75.04012, 75.03331, 75.00368, 74.99545, 74.97292, 74.95422, 
    74.97128, 74.98917, 75.0402, 75.08569, 75.1358, 75.14811, 75.20631, 
    75.15874, 75.23704, 75.17019, 75.28605, 75.07832, 75.1685, 75.00575, 
    75.02337, 75.05465, 75.12767, 75.08839, 75.1344, 75.03306, 74.98009, 
    74.96656, 74.94103, 74.96714, 74.96503, 74.99, 74.98198, 75.04189, 
    75.00971, 75.10074, 75.13406, 75.22836, 75.28607, 75.34502, 75.37098, 
    75.37889, 75.38219 ;

 FIRA_R =
  74.74778, 74.80091, 74.79061, 74.83339, 74.80971, 74.83768, 74.75861, 
    74.80296, 74.77468, 74.75264, 74.9163, 74.83531, 75.00118, 74.9493, 
    75.07941, 74.99303, 75.09693, 75.07703, 75.13724, 75.12, 75.19672, 
    75.1452, 75.2367, 75.18449, 75.1926, 75.14348, 74.85173, 74.90617, 
    74.84848, 74.85625, 74.85279, 74.81015, 74.78858, 74.7438, 74.75196, 
    74.7849, 74.85974, 74.83441, 74.89851, 74.89707, 74.96848, 74.93624, 
    75.05608, 75.02235, 75.12072, 75.09586, 75.11953, 75.11237, 75.11962, 
    75.08316, 75.09878, 75.06673, 74.94225, 74.97892, 74.86966, 74.80388, 
    74.76054, 74.72967, 74.73403, 74.74232, 74.78509, 74.8254, 74.8561, 
    74.87663, 74.89686, 74.95787, 74.99049, 75.06291, 75.04988, 75.07205, 
    75.09338, 75.12906, 75.12321, 75.13889, 75.07155, 75.11626, 75.04286, 
    75.06261, 74.90192, 74.84126, 74.81512, 74.79257, 74.73738, 74.77547, 
    74.76044, 74.79629, 74.81899, 74.80779, 74.87718, 74.85017, 74.99243, 
    74.93108, 75.0909, 75.05257, 75.10011, 75.07587, 75.11736, 75.08002, 
    75.14477, 75.15881, 75.14921, 75.18626, 75.07793, 75.11949, 74.80745, 
    74.80927, 74.81783, 74.7802, 74.77792, 74.74356, 74.77418, 74.78718, 
    74.82035, 74.83989, 74.85851, 74.89945, 74.94515, 75.0093, 75.05505, 
    75.08597, 75.06704, 75.08375, 75.06505, 75.0563, 75.15352, 75.09889, 
    75.18093, 75.17641, 75.13924, 75.17693, 74.81056, 74.80004, 74.76336, 
    74.79207, 74.73983, 74.76901, 74.78576, 74.85065, 74.86501, 74.8782, 
    74.90435, 74.93789, 74.9968, 75.04771, 75.09465, 75.09122, 75.09242, 
    75.10286, 75.07694, 75.10712, 75.11214, 75.09895, 75.1758, 75.15385, 
    75.17632, 75.16203, 74.80347, 74.8212, 74.81161, 74.82961, 74.81689, 
    74.87335, 74.89027, 74.96974, 74.9372, 74.98912, 74.94251, 74.95074, 
    74.99062, 74.94506, 75.04523, 74.97714, 75.10326, 75.03552, 75.10753, 
    75.09444, 75.11615, 75.13554, 75.16001, 75.20504, 75.19463, 75.23236, 
    74.84767, 74.87065, 74.86871, 74.89281, 74.91061, 74.94937, 75.01151, 
    74.98817, 75.03111, 75.03971, 74.97451, 75.01446, 74.88609, 74.90669, 
    74.89449, 74.84944, 74.99343, 74.91939, 75.05579, 75.01611, 75.13276, 
    75.07445, 75.18888, 75.23758, 75.2838, 75.33734, 74.88328, 74.86766, 
    74.8957, 74.93436, 74.97055, 75.01854, 75.0235, 75.03246, 75.05537, 
    75.07494, 75.03522, 75.07986, 74.91131, 74.99989, 74.86167, 74.90312, 
    74.93212, 74.91946, 74.98552, 75.00106, 75.06377, 75.03162, 75.22549, 
    75.13951, 75.3784, 75.31159, 74.86218, 74.88326, 74.9566, 74.92167, 
    75.02179, 75.0464, 75.06606, 75.09159, 75.09441, 75.10955, 75.08473, 
    75.1086, 75.01864, 75.05862, 74.9483, 74.9752, 74.96285, 74.94925, 
    74.99123, 75.03583, 75.03692, 75.05077, 75.09075, 75.02219, 75.23633, 
    75.10359, 74.90623, 74.94672, 74.95267, 74.93694, 75.04393, 75.00513, 
    75.1092, 75.08099, 75.12724, 75.10425, 75.10086, 75.07135, 75.05295, 
    75.00689, 74.96912, 74.93924, 74.9462, 74.97903, 75.03859, 75.0946, 
    75.08222, 75.12373, 75.01452, 75.06, 75.04264, 75.08862, 74.98752, 
    75.07313, 74.96548, 74.97498, 75.00437, 75.06302, 75.07629, 75.09022, 
    75.08165, 75.04012, 75.03331, 75.00368, 74.99545, 74.97292, 74.95422, 
    74.97128, 74.98917, 75.0402, 75.08569, 75.1358, 75.14811, 75.20631, 
    75.15874, 75.23704, 75.17019, 75.28605, 75.07832, 75.1685, 75.00575, 
    75.02337, 75.05465, 75.12767, 75.08839, 75.1344, 75.03306, 74.98009, 
    74.96656, 74.94103, 74.96714, 74.96503, 74.99, 74.98198, 75.04189, 
    75.00971, 75.10074, 75.13406, 75.22836, 75.28607, 75.34502, 75.37098, 
    75.37889, 75.38219 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.7087, 263.7618, 263.7516, 263.7943, 263.7706, 263.7986, 263.7195, 
    263.7639, 263.7356, 263.7136, 263.8772, 263.7962, 263.9621, 263.9102, 
    264.0403, 263.954, 264.0579, 264.038, 264.0982, 264.0809, 264.1577, 
    264.1061, 264.1976, 264.1454, 264.1535, 264.1044, 263.8127, 263.8671, 
    263.8094, 263.8172, 263.8137, 263.7711, 263.7495, 263.7047, 263.7129, 
    263.7458, 263.8207, 263.7953, 263.8595, 263.858, 263.9294, 263.8972, 
    264.017, 263.9833, 264.0817, 264.0568, 264.0805, 264.0733, 264.0806, 
    264.0441, 264.0597, 264.0277, 263.9032, 263.9398, 263.8306, 263.7648, 
    263.7215, 263.6906, 263.695, 263.7033, 263.746, 263.7863, 263.817, 
    263.8376, 263.8578, 263.9188, 263.9514, 264.0239, 264.0108, 264.033, 
    264.0543, 264.09, 264.0841, 264.0998, 264.0325, 264.0772, 264.0038, 
    264.0236, 263.8629, 263.8022, 263.7761, 263.7535, 263.6983, 263.7364, 
    263.7214, 263.7572, 263.7799, 263.7687, 263.8381, 263.8111, 263.9534, 
    263.892, 264.0518, 264.0135, 264.061, 264.0368, 264.0783, 264.041, 
    264.1057, 264.1198, 264.1101, 264.1472, 264.0389, 264.0804, 263.7684, 
    263.7702, 263.7788, 263.7411, 263.7389, 263.7045, 263.7351, 263.7481, 
    263.7813, 263.8008, 263.8195, 263.8604, 263.9061, 263.9702, 264.016, 
    264.0469, 264.028, 264.0447, 264.026, 264.0172, 264.1145, 264.0598, 
    264.1419, 264.1374, 264.1002, 264.1378, 263.7715, 263.761, 263.7243, 
    263.753, 263.7008, 263.7299, 263.7467, 263.8116, 263.826, 263.8391, 
    263.8653, 263.8988, 263.9577, 264.0087, 264.0556, 264.0522, 264.0533, 
    264.0638, 264.0379, 264.0681, 264.0731, 264.0599, 264.1367, 264.1148, 
    264.1373, 264.123, 263.7644, 263.7821, 263.7726, 263.7906, 263.7778, 
    263.8343, 263.8512, 263.9307, 263.8981, 263.95, 263.9034, 263.9117, 
    263.9516, 263.906, 264.0062, 263.9381, 264.0642, 263.9965, 264.0685, 
    264.0554, 264.0771, 264.0965, 264.1209, 264.166, 264.1556, 264.1933, 
    263.8086, 263.8316, 263.8297, 263.8538, 263.8716, 263.9103, 263.9724, 
    263.9491, 263.9921, 264.0006, 263.9355, 263.9754, 263.847, 263.8676, 
    263.8554, 263.8104, 263.9544, 263.8803, 264.0167, 263.9771, 264.0937, 
    264.0354, 264.1498, 264.1985, 264.2447, 264.2983, 263.8442, 263.8286, 
    263.8566, 263.8953, 263.9315, 263.9795, 263.9844, 263.9934, 264.0163, 
    264.0359, 263.9962, 264.0408, 263.8723, 263.9608, 263.8226, 263.8641, 
    263.8931, 263.8804, 263.9465, 263.962, 264.0247, 263.9926, 264.1864, 
    264.1005, 264.3393, 264.2725, 263.8231, 263.8442, 263.9175, 263.8826, 
    263.9827, 264.0074, 264.027, 264.0525, 264.0554, 264.0705, 264.0457, 
    264.0695, 263.9796, 264.0196, 263.9092, 263.9361, 263.9238, 263.9102, 
    263.9522, 263.9968, 263.9979, 264.0117, 264.0517, 263.9831, 264.1973, 
    264.0645, 263.8672, 263.9077, 263.9136, 263.8979, 264.0049, 263.9661, 
    264.0701, 264.0419, 264.0882, 264.0652, 264.0618, 264.0323, 264.0139, 
    263.9678, 263.9301, 263.9002, 263.9071, 263.94, 263.9995, 264.0555, 
    264.0432, 264.0847, 263.9755, 264.0209, 264.0036, 264.0496, 263.9485, 
    264.0341, 263.9264, 263.9359, 263.9653, 264.024, 264.0372, 264.0511, 
    264.0426, 264.0011, 263.9943, 263.9646, 263.9564, 263.9339, 263.9152, 
    263.9322, 263.9501, 264.0011, 264.0466, 264.0967, 264.109, 264.1672, 
    264.1197, 264.198, 264.1311, 264.247, 264.0392, 264.1295, 263.9667, 
    263.9843, 264.0156, 264.0886, 264.0493, 264.0953, 263.994, 263.941, 
    263.9275, 263.902, 263.9281, 263.926, 263.9509, 263.9429, 264.0028, 
    263.9706, 264.0617, 264.095, 264.1893, 264.247, 264.306, 264.3319, 
    264.3398, 264.3431 ;

 FIRE_R =
  263.7087, 263.7618, 263.7516, 263.7943, 263.7706, 263.7986, 263.7195, 
    263.7639, 263.7356, 263.7136, 263.8772, 263.7962, 263.9621, 263.9102, 
    264.0403, 263.954, 264.0579, 264.038, 264.0982, 264.0809, 264.1577, 
    264.1061, 264.1976, 264.1454, 264.1535, 264.1044, 263.8127, 263.8671, 
    263.8094, 263.8172, 263.8137, 263.7711, 263.7495, 263.7047, 263.7129, 
    263.7458, 263.8207, 263.7953, 263.8595, 263.858, 263.9294, 263.8972, 
    264.017, 263.9833, 264.0817, 264.0568, 264.0805, 264.0733, 264.0806, 
    264.0441, 264.0597, 264.0277, 263.9032, 263.9398, 263.8306, 263.7648, 
    263.7215, 263.6906, 263.695, 263.7033, 263.746, 263.7863, 263.817, 
    263.8376, 263.8578, 263.9188, 263.9514, 264.0239, 264.0108, 264.033, 
    264.0543, 264.09, 264.0841, 264.0998, 264.0325, 264.0772, 264.0038, 
    264.0236, 263.8629, 263.8022, 263.7761, 263.7535, 263.6983, 263.7364, 
    263.7214, 263.7572, 263.7799, 263.7687, 263.8381, 263.8111, 263.9534, 
    263.892, 264.0518, 264.0135, 264.061, 264.0368, 264.0783, 264.041, 
    264.1057, 264.1198, 264.1101, 264.1472, 264.0389, 264.0804, 263.7684, 
    263.7702, 263.7788, 263.7411, 263.7389, 263.7045, 263.7351, 263.7481, 
    263.7813, 263.8008, 263.8195, 263.8604, 263.9061, 263.9702, 264.016, 
    264.0469, 264.028, 264.0447, 264.026, 264.0172, 264.1145, 264.0598, 
    264.1419, 264.1374, 264.1002, 264.1378, 263.7715, 263.761, 263.7243, 
    263.753, 263.7008, 263.7299, 263.7467, 263.8116, 263.826, 263.8391, 
    263.8653, 263.8988, 263.9577, 264.0087, 264.0556, 264.0522, 264.0533, 
    264.0638, 264.0379, 264.0681, 264.0731, 264.0599, 264.1367, 264.1148, 
    264.1373, 264.123, 263.7644, 263.7821, 263.7726, 263.7906, 263.7778, 
    263.8343, 263.8512, 263.9307, 263.8981, 263.95, 263.9034, 263.9117, 
    263.9516, 263.906, 264.0062, 263.9381, 264.0642, 263.9965, 264.0685, 
    264.0554, 264.0771, 264.0965, 264.1209, 264.166, 264.1556, 264.1933, 
    263.8086, 263.8316, 263.8297, 263.8538, 263.8716, 263.9103, 263.9724, 
    263.9491, 263.9921, 264.0006, 263.9355, 263.9754, 263.847, 263.8676, 
    263.8554, 263.8104, 263.9544, 263.8803, 264.0167, 263.9771, 264.0937, 
    264.0354, 264.1498, 264.1985, 264.2447, 264.2983, 263.8442, 263.8286, 
    263.8566, 263.8953, 263.9315, 263.9795, 263.9844, 263.9934, 264.0163, 
    264.0359, 263.9962, 264.0408, 263.8723, 263.9608, 263.8226, 263.8641, 
    263.8931, 263.8804, 263.9465, 263.962, 264.0247, 263.9926, 264.1864, 
    264.1005, 264.3393, 264.2725, 263.8231, 263.8442, 263.9175, 263.8826, 
    263.9827, 264.0074, 264.027, 264.0525, 264.0554, 264.0705, 264.0457, 
    264.0695, 263.9796, 264.0196, 263.9092, 263.9361, 263.9238, 263.9102, 
    263.9522, 263.9968, 263.9979, 264.0117, 264.0517, 263.9831, 264.1973, 
    264.0645, 263.8672, 263.9077, 263.9136, 263.8979, 264.0049, 263.9661, 
    264.0701, 264.0419, 264.0882, 264.0652, 264.0618, 264.0323, 264.0139, 
    263.9678, 263.9301, 263.9002, 263.9071, 263.94, 263.9995, 264.0555, 
    264.0432, 264.0847, 263.9755, 264.0209, 264.0036, 264.0496, 263.9485, 
    264.0341, 263.9264, 263.9359, 263.9653, 264.024, 264.0372, 264.0511, 
    264.0426, 264.0011, 263.9943, 263.9646, 263.9564, 263.9339, 263.9152, 
    263.9322, 263.9501, 264.0011, 264.0466, 264.0967, 264.109, 264.1672, 
    264.1197, 264.198, 264.1311, 264.247, 264.0392, 264.1295, 263.9667, 
    263.9843, 264.0156, 264.0886, 264.0493, 264.0953, 263.994, 263.941, 
    263.9275, 263.902, 263.9281, 263.926, 263.9509, 263.9429, 264.0028, 
    263.9706, 264.0617, 264.095, 264.1893, 264.247, 264.306, 264.3319, 
    264.3398, 264.3431 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  242.9372, 243.6305, 243.4961, 244.0545, 243.7454, 244.1105, 243.0785, 
    243.6574, 243.2883, 243.0007, 245.1355, 244.0796, 246.237, 245.564, 
    247.2658, 246.1313, 247.493, 247.235, 248.0158, 247.7922, 248.7876, 
    248.119, 249.3063, 248.6288, 248.7342, 248.0967, 244.2937, 245.0035, 
    244.2513, 244.3526, 244.3075, 243.7512, 243.4697, 242.8854, 242.9918, 
    243.4216, 244.3982, 244.0679, 244.9036, 244.8847, 245.8127, 245.3946, 
    246.9632, 246.5113, 247.8016, 247.479, 247.7861, 247.6932, 247.7873, 
    247.3144, 247.517, 247.1014, 245.4727, 245.9482, 244.5274, 243.6694, 
    243.1036, 242.7009, 242.7579, 242.866, 243.4241, 243.9503, 244.3506, 
    244.6181, 244.882, 245.6754, 246.0984, 247.0519, 246.8828, 247.1703, 
    247.447, 247.9097, 247.8338, 248.0373, 247.1638, 247.7438, 246.7771, 
    247.0479, 244.9481, 244.1572, 243.8161, 243.5218, 242.8015, 243.2986, 
    243.1025, 243.5702, 243.8666, 243.7203, 244.6255, 244.2734, 246.1235, 
    245.3275, 247.4148, 246.9176, 247.5341, 247.2198, 247.7579, 247.2737, 
    248.1135, 248.2957, 248.1711, 248.6519, 247.2466, 247.7856, 243.7159, 
    243.7397, 243.8515, 243.3603, 243.3306, 242.8822, 243.2816, 243.4513, 
    243.8843, 244.1393, 244.382, 244.9158, 245.5103, 246.3423, 246.9498, 
    247.3508, 247.1053, 247.322, 247.0795, 246.9661, 248.2271, 247.5185, 
    248.5827, 248.524, 248.0419, 248.5306, 243.7566, 243.6192, 243.1405, 
    243.5152, 242.8335, 243.2143, 243.4329, 244.2795, 244.4668, 244.6387, 
    244.9796, 245.416, 246.1801, 246.8548, 247.4634, 247.4189, 247.4345, 
    247.5699, 247.2337, 247.6251, 247.6903, 247.5191, 248.5161, 248.2313, 
    248.5227, 248.3374, 243.664, 243.8954, 243.7703, 244.0052, 243.8392, 
    244.5755, 244.7962, 245.8293, 245.4071, 246.0805, 245.476, 245.5828, 
    246.1001, 245.509, 246.8079, 245.9252, 247.5752, 246.6822, 247.6304, 
    247.4607, 247.7422, 247.9938, 248.3112, 248.8955, 248.7604, 249.2499, 
    244.2408, 244.5403, 244.515, 244.8291, 245.0613, 245.5649, 246.3708, 
    246.0681, 246.6249, 246.7363, 245.891, 246.409, 244.7415, 245.0103, 
    244.851, 244.2638, 246.1364, 245.1758, 246.9595, 246.4304, 247.9578, 
    247.2015, 248.6858, 249.3177, 249.9174, 250.6126, 244.7049, 244.5013, 
    244.8668, 245.3703, 245.8396, 246.4619, 246.5261, 246.6424, 246.9539, 
    247.2077, 246.6781, 247.2715, 245.0705, 246.2203, 244.4233, 244.9637, 
    245.3411, 245.1768, 246.0338, 246.2353, 247.0631, 246.6313, 249.1609, 
    248.0454, 251.1454, 250.2783, 244.4299, 244.7047, 245.6587, 245.2054, 
    246.504, 246.8231, 247.0926, 247.4237, 247.4603, 247.6566, 247.3347, 
    247.6443, 246.4632, 246.9961, 245.551, 245.8999, 245.7398, 245.5633, 
    246.1078, 246.6861, 246.7001, 246.8943, 247.4132, 246.5093, 249.3017, 
    247.5796, 245.0043, 245.5306, 245.6078, 245.4037, 246.791, 246.2882, 
    247.6521, 247.2862, 247.8862, 247.5879, 247.5439, 247.1613, 246.9226, 
    246.311, 245.8211, 245.4335, 245.5238, 245.9496, 246.7218, 247.4628, 
    247.3022, 247.8406, 246.4098, 247.014, 246.7743, 247.3851, 246.0597, 
    247.1846, 245.7738, 245.8971, 246.2783, 247.0533, 247.2253, 247.4059, 
    247.2948, 246.7417, 246.6534, 246.2694, 246.1625, 245.8704, 245.6277, 
    245.849, 246.0811, 246.7427, 247.3472, 247.9971, 248.1568, 248.9121, 
    248.2949, 249.311, 248.4436, 249.9469, 247.2517, 248.4215, 246.2962, 
    246.5245, 246.9448, 247.8918, 247.3823, 247.979, 246.6501, 245.9634, 
    245.7878, 245.4568, 245.7954, 245.7679, 246.0919, 245.9879, 246.7647, 
    246.3475, 247.5424, 247.9747, 249.198, 249.947, 250.7122, 251.0491, 
    251.1518, 251.1947 ;

 FSH_G =
  256.0403, 256.7346, 256.5999, 257.1591, 256.8495, 257.2152, 256.1817, 
    256.7614, 256.3918, 256.1038, 258.2417, 257.1843, 259.3448, 258.6708, 
    260.3749, 259.2389, 260.6025, 260.3441, 261.1261, 260.9021, 261.8989, 
    261.2294, 262.4184, 261.7399, 261.8454, 261.2071, 257.3987, 258.1095, 
    257.3562, 257.4576, 257.4125, 256.8554, 256.5735, 255.9883, 256.0949, 
    256.5253, 257.5033, 257.1725, 258.0094, 257.9906, 258.9199, 258.5012, 
    260.0719, 259.6194, 260.9115, 260.5885, 260.8961, 260.803, 260.8973, 
    260.4237, 260.6265, 260.2103, 258.5793, 259.0555, 257.6327, 256.7734, 
    256.2069, 255.8036, 255.8606, 255.9689, 256.5278, 257.0547, 257.4557, 
    257.7236, 257.9878, 258.7823, 259.2059, 260.1608, 259.9915, 260.2794, 
    260.5565, 261.0198, 260.9438, 261.1476, 260.2728, 260.8536, 259.8856, 
    260.1568, 258.0539, 257.262, 256.9203, 256.6256, 255.9043, 256.4021, 
    256.2057, 256.6742, 256.971, 256.8244, 257.7309, 257.3784, 259.231, 
    258.434, 260.5242, 260.0263, 260.6437, 260.3289, 260.8678, 260.3828, 
    261.2239, 261.4064, 261.2815, 261.763, 260.3558, 260.8955, 256.82, 
    256.8439, 256.9558, 256.4639, 256.4341, 255.9851, 256.3852, 256.5551, 
    256.9886, 257.244, 257.4871, 258.0216, 258.6171, 259.4502, 260.0585, 
    260.4601, 260.2143, 260.4313, 260.1884, 260.0749, 261.3376, 260.6281, 
    261.6938, 261.635, 261.1522, 261.6416, 256.8607, 256.7232, 256.2438, 
    256.619, 255.9363, 256.3177, 256.5366, 257.3845, 257.5721, 257.7442, 
    258.0856, 258.5226, 259.2878, 259.9634, 260.5728, 260.5283, 260.5439, 
    260.6795, 260.3429, 260.7348, 260.8, 260.6286, 261.6271, 261.3419, 
    261.6337, 261.4482, 256.7681, 256.9998, 256.8745, 257.1098, 256.9435, 
    257.6809, 257.9019, 258.9364, 258.5137, 259.188, 258.5827, 258.6896, 
    259.2076, 258.6158, 259.9165, 259.0325, 260.6848, 259.7905, 260.7401, 
    260.5702, 260.8521, 261.104, 261.4219, 262.007, 261.8717, 262.362, 
    257.3457, 257.6456, 257.6203, 257.9349, 258.1673, 258.6717, 259.4787, 
    259.1756, 259.7332, 259.8448, 258.9982, 259.517, 257.8471, 258.1163, 
    257.9568, 257.3687, 259.244, 258.282, 260.0682, 259.5384, 261.0679, 
    260.3106, 261.797, 262.4298, 263.0304, 263.7265, 257.8105, 257.6065, 
    257.9726, 258.4768, 258.9468, 259.57, 259.6343, 259.7507, 260.0627, 
    260.3169, 259.7865, 260.3807, 258.1765, 259.328, 257.5285, 258.0696, 
    258.4476, 258.283, 259.1412, 259.3431, 260.172, 259.7397, 262.2727, 
    261.1557, 264.2602, 263.3918, 257.535, 257.8102, 258.7656, 258.3117, 
    259.6122, 259.9317, 260.2015, 260.5331, 260.5697, 260.7664, 260.444, 
    260.7541, 259.5713, 260.1049, 258.6578, 259.0072, 258.8468, 258.6701, 
    259.2154, 259.7944, 259.8085, 260.003, 260.5225, 259.6174, 262.4138, 
    260.6892, 258.1103, 258.6374, 258.7146, 258.5103, 259.8996, 259.3961, 
    260.7618, 260.3954, 260.9962, 260.6975, 260.6535, 260.2703, 260.0313, 
    259.4188, 258.9283, 258.5401, 258.6305, 259.0569, 259.8302, 260.5723, 
    260.4115, 260.9506, 259.5178, 260.1229, 259.8828, 260.4944, 259.1671, 
    260.2936, 258.881, 259.0044, 259.3861, 260.1621, 260.3344, 260.5153, 
    260.4041, 259.8502, 259.7617, 259.3772, 259.2702, 258.9776, 258.7346, 
    258.9562, 259.1886, 259.8511, 260.4565, 261.1073, 261.2673, 262.0236, 
    261.4055, 262.423, 261.5544, 263.0599, 260.3608, 261.5323, 259.404, 
    259.6327, 260.0535, 261.0019, 260.4916, 261.0892, 259.7584, 259.0708, 
    258.895, 258.5634, 258.9025, 258.875, 259.1994, 259.0953, 259.8732, 
    259.4554, 260.6519, 261.0849, 262.31, 263.06, 263.8263, 264.1638, 
    264.2666, 264.3095 ;

 FSH_NODYNLNDUSE =
  242.9372, 243.6305, 243.4961, 244.0545, 243.7454, 244.1105, 243.0785, 
    243.6574, 243.2883, 243.0007, 245.1355, 244.0796, 246.237, 245.564, 
    247.2658, 246.1313, 247.493, 247.235, 248.0158, 247.7922, 248.7876, 
    248.119, 249.3063, 248.6288, 248.7342, 248.0967, 244.2937, 245.0035, 
    244.2513, 244.3526, 244.3075, 243.7512, 243.4697, 242.8854, 242.9918, 
    243.4216, 244.3982, 244.0679, 244.9036, 244.8847, 245.8127, 245.3946, 
    246.9632, 246.5113, 247.8016, 247.479, 247.7861, 247.6932, 247.7873, 
    247.3144, 247.517, 247.1014, 245.4727, 245.9482, 244.5274, 243.6694, 
    243.1036, 242.7009, 242.7579, 242.866, 243.4241, 243.9503, 244.3506, 
    244.6181, 244.882, 245.6754, 246.0984, 247.0519, 246.8828, 247.1703, 
    247.447, 247.9097, 247.8338, 248.0373, 247.1638, 247.7438, 246.7771, 
    247.0479, 244.9481, 244.1572, 243.8161, 243.5218, 242.8015, 243.2986, 
    243.1025, 243.5702, 243.8666, 243.7203, 244.6255, 244.2734, 246.1235, 
    245.3275, 247.4148, 246.9176, 247.5341, 247.2198, 247.7579, 247.2737, 
    248.1135, 248.2957, 248.1711, 248.6519, 247.2466, 247.7856, 243.7159, 
    243.7397, 243.8515, 243.3603, 243.3306, 242.8822, 243.2816, 243.4513, 
    243.8843, 244.1393, 244.382, 244.9158, 245.5103, 246.3423, 246.9498, 
    247.3508, 247.1053, 247.322, 247.0795, 246.9661, 248.2271, 247.5185, 
    248.5827, 248.524, 248.0419, 248.5306, 243.7566, 243.6192, 243.1405, 
    243.5152, 242.8335, 243.2143, 243.4329, 244.2795, 244.4668, 244.6387, 
    244.9796, 245.416, 246.1801, 246.8548, 247.4634, 247.4189, 247.4345, 
    247.5699, 247.2337, 247.6251, 247.6903, 247.5191, 248.5161, 248.2313, 
    248.5227, 248.3374, 243.664, 243.8954, 243.7703, 244.0052, 243.8392, 
    244.5755, 244.7962, 245.8293, 245.4071, 246.0805, 245.476, 245.5828, 
    246.1001, 245.509, 246.8079, 245.9252, 247.5752, 246.6822, 247.6304, 
    247.4607, 247.7422, 247.9938, 248.3112, 248.8955, 248.7604, 249.2499, 
    244.2408, 244.5403, 244.515, 244.8291, 245.0613, 245.5649, 246.3708, 
    246.0681, 246.6249, 246.7363, 245.891, 246.409, 244.7415, 245.0103, 
    244.851, 244.2638, 246.1364, 245.1758, 246.9595, 246.4304, 247.9578, 
    247.2015, 248.6858, 249.3177, 249.9174, 250.6126, 244.7049, 244.5013, 
    244.8668, 245.3703, 245.8396, 246.4619, 246.5261, 246.6424, 246.9539, 
    247.2077, 246.6781, 247.2715, 245.0705, 246.2203, 244.4233, 244.9637, 
    245.3411, 245.1768, 246.0338, 246.2353, 247.0631, 246.6313, 249.1609, 
    248.0454, 251.1454, 250.2783, 244.4299, 244.7047, 245.6587, 245.2054, 
    246.504, 246.8231, 247.0926, 247.4237, 247.4603, 247.6566, 247.3347, 
    247.6443, 246.4632, 246.9961, 245.551, 245.8999, 245.7398, 245.5633, 
    246.1078, 246.6861, 246.7001, 246.8943, 247.4132, 246.5093, 249.3017, 
    247.5796, 245.0043, 245.5306, 245.6078, 245.4037, 246.791, 246.2882, 
    247.6521, 247.2862, 247.8862, 247.5879, 247.5439, 247.1613, 246.9226, 
    246.311, 245.8211, 245.4335, 245.5238, 245.9496, 246.7218, 247.4628, 
    247.3022, 247.8406, 246.4098, 247.014, 246.7743, 247.3851, 246.0597, 
    247.1846, 245.7738, 245.8971, 246.2783, 247.0533, 247.2253, 247.4059, 
    247.2948, 246.7417, 246.6534, 246.2694, 246.1625, 245.8704, 245.6277, 
    245.849, 246.0811, 246.7427, 247.3472, 247.9971, 248.1568, 248.9121, 
    248.2949, 249.311, 248.4436, 249.9469, 247.2517, 248.4215, 246.2962, 
    246.5245, 246.9448, 247.8918, 247.3823, 247.979, 246.6501, 245.9634, 
    245.7878, 245.4568, 245.7954, 245.7679, 246.0919, 245.9879, 246.7647, 
    246.3475, 247.5424, 247.9747, 249.198, 249.947, 250.7122, 251.0491, 
    251.1518, 251.1947 ;

 FSH_R =
  242.9372, 243.6305, 243.4961, 244.0545, 243.7454, 244.1105, 243.0785, 
    243.6574, 243.2883, 243.0007, 245.1355, 244.0796, 246.237, 245.564, 
    247.2658, 246.1313, 247.493, 247.235, 248.0158, 247.7922, 248.7876, 
    248.119, 249.3063, 248.6288, 248.7342, 248.0967, 244.2937, 245.0035, 
    244.2513, 244.3526, 244.3075, 243.7512, 243.4697, 242.8854, 242.9918, 
    243.4216, 244.3982, 244.0679, 244.9036, 244.8847, 245.8127, 245.3946, 
    246.9632, 246.5113, 247.8016, 247.479, 247.7861, 247.6932, 247.7873, 
    247.3144, 247.517, 247.1014, 245.4727, 245.9482, 244.5274, 243.6694, 
    243.1036, 242.7009, 242.7579, 242.866, 243.4241, 243.9503, 244.3506, 
    244.6181, 244.882, 245.6754, 246.0984, 247.0519, 246.8828, 247.1703, 
    247.447, 247.9097, 247.8338, 248.0373, 247.1638, 247.7438, 246.7771, 
    247.0479, 244.9481, 244.1572, 243.8161, 243.5218, 242.8015, 243.2986, 
    243.1025, 243.5702, 243.8666, 243.7203, 244.6255, 244.2734, 246.1235, 
    245.3275, 247.4148, 246.9176, 247.5341, 247.2198, 247.7579, 247.2737, 
    248.1135, 248.2957, 248.1711, 248.6519, 247.2466, 247.7856, 243.7159, 
    243.7397, 243.8515, 243.3603, 243.3306, 242.8822, 243.2816, 243.4513, 
    243.8843, 244.1393, 244.382, 244.9158, 245.5103, 246.3423, 246.9498, 
    247.3508, 247.1053, 247.322, 247.0795, 246.9661, 248.2271, 247.5185, 
    248.5827, 248.524, 248.0419, 248.5306, 243.7566, 243.6192, 243.1405, 
    243.5152, 242.8335, 243.2143, 243.4329, 244.2795, 244.4668, 244.6387, 
    244.9796, 245.416, 246.1801, 246.8548, 247.4634, 247.4189, 247.4345, 
    247.5699, 247.2337, 247.6251, 247.6903, 247.5191, 248.5161, 248.2313, 
    248.5227, 248.3374, 243.664, 243.8954, 243.7703, 244.0052, 243.8392, 
    244.5755, 244.7962, 245.8293, 245.4071, 246.0805, 245.476, 245.5828, 
    246.1001, 245.509, 246.8079, 245.9252, 247.5752, 246.6822, 247.6304, 
    247.4607, 247.7422, 247.9938, 248.3112, 248.8955, 248.7604, 249.2499, 
    244.2408, 244.5403, 244.515, 244.8291, 245.0613, 245.5649, 246.3708, 
    246.0681, 246.6249, 246.7363, 245.891, 246.409, 244.7415, 245.0103, 
    244.851, 244.2638, 246.1364, 245.1758, 246.9595, 246.4304, 247.9578, 
    247.2015, 248.6858, 249.3177, 249.9174, 250.6126, 244.7049, 244.5013, 
    244.8668, 245.3703, 245.8396, 246.4619, 246.5261, 246.6424, 246.9539, 
    247.2077, 246.6781, 247.2715, 245.0705, 246.2203, 244.4233, 244.9637, 
    245.3411, 245.1768, 246.0338, 246.2353, 247.0631, 246.6313, 249.1609, 
    248.0454, 251.1454, 250.2783, 244.4299, 244.7047, 245.6587, 245.2054, 
    246.504, 246.8231, 247.0926, 247.4237, 247.4603, 247.6566, 247.3347, 
    247.6443, 246.4632, 246.9961, 245.551, 245.8999, 245.7398, 245.5633, 
    246.1078, 246.6861, 246.7001, 246.8943, 247.4132, 246.5093, 249.3017, 
    247.5796, 245.0043, 245.5306, 245.6078, 245.4037, 246.791, 246.2882, 
    247.6521, 247.2862, 247.8862, 247.5879, 247.5439, 247.1613, 246.9226, 
    246.311, 245.8211, 245.4335, 245.5238, 245.9496, 246.7218, 247.4628, 
    247.3022, 247.8406, 246.4098, 247.014, 246.7743, 247.3851, 246.0597, 
    247.1846, 245.7738, 245.8971, 246.2783, 247.0533, 247.2253, 247.4059, 
    247.2948, 246.7417, 246.6534, 246.2694, 246.1625, 245.8704, 245.6277, 
    245.849, 246.0811, 246.7427, 247.3472, 247.9971, 248.1568, 248.9121, 
    248.2949, 249.311, 248.4436, 249.9469, 247.2517, 248.4215, 246.2962, 
    246.5245, 246.9448, 247.8918, 247.3823, 247.979, 246.6501, 245.9634, 
    245.7878, 245.4568, 245.7954, 245.7679, 246.0919, 245.9879, 246.7647, 
    246.3475, 247.5424, 247.9747, 249.198, 249.947, 250.7122, 251.0491, 
    251.1518, 251.1947 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.10301, -13.10401, -13.10382, -13.10462, -13.10418, -13.1047, -13.10322, 
    -13.10404, -13.10352, -13.10311, -13.10614, -13.10465, -13.10773, 
    -13.10679, -13.10917, -13.10757, -13.1095, -13.10914, -13.11026, 
    -13.10994, -13.11133, -13.11041, -13.11209, -13.11112, -13.11127, 
    -13.11037, -13.10497, -13.10595, -13.10491, -13.10505, -13.10499, 
    -13.10418, -13.10377, -13.10295, -13.1031, -13.10371, -13.10511, 
    -13.10465, -13.10586, -13.10583, -13.10715, -13.10656, -13.10875, 
    -13.10814, -13.10995, -13.10949, -13.10993, -13.1098, -13.10993, 
    -13.10925, -13.10954, -13.10895, -13.10666, -13.10733, -13.1053, 
    -13.10404, -13.10326, -13.10268, -13.10276, -13.10291, -13.10371, 
    -13.10448, -13.10506, -13.10544, -13.10583, -13.10692, -13.10753, 
    -13.10887, -13.10864, -13.10904, -13.10944, -13.1101, -13.11, -13.11028, 
    -13.10904, -13.10986, -13.10852, -13.10888, -13.10586, -13.10478, 
    -13.10426, -13.10385, -13.10282, -13.10353, -13.10325, -13.10393, 
    -13.10436, -13.10415, -13.10545, -13.10494, -13.10757, -13.10645, 
    -13.1094, -13.10869, -13.10957, -13.10912, -13.10988, -13.1092, 
    -13.11039, -13.11065, -13.11047, -13.11117, -13.10916, -13.10992, 
    -13.10414, -13.10417, -13.10434, -13.10362, -13.10358, -13.10294, 
    -13.10351, -13.10375, -13.10439, -13.10475, -13.1051, -13.10587, 
    -13.10671, -13.10789, -13.10874, -13.10931, -13.10896, -13.10927, 
    -13.10892, -13.10877, -13.11055, -13.10954, -13.11107, -13.11098, 
    -13.11029, -13.11099, -13.1042, -13.104, -13.10331, -13.10385, -13.10287, 
    -13.10341, -13.10372, -13.10494, -13.10523, -13.10547, -13.10597, 
    -13.10659, -13.10766, -13.1086, -13.10947, -13.10941, -13.10943, 
    -13.10962, -13.10914, -13.1097, -13.10979, -13.10955, -13.11097, 
    -13.11056, -13.11098, -13.11072, -13.10407, -13.1044, -13.10422, 
    -13.10455, -13.10431, -13.10536, -13.10568, -13.10715, -13.10657, 
    -13.10752, -13.10667, -13.10682, -13.10752, -13.10672, -13.10854, 
    -13.10728, -13.10963, -13.10835, -13.10971, -13.10947, -13.10987, 
    -13.11022, -13.11068, -13.1115, -13.11131, -13.11202, -13.1049, 
    -13.10532, -13.1053, -13.10575, -13.10608, -13.1068, -13.10794, 
    -13.10751, -13.1083, -13.10846, -13.10726, -13.10798, -13.10561, 
    -13.10599, -13.10577, -13.10492, -13.10759, -13.10623, -13.10875, 
    -13.10802, -13.11017, -13.10908, -13.11121, -13.11209, -13.11299, 
    -13.11397, -13.10557, -13.10528, -13.10581, -13.10651, -13.10718, 
    -13.10807, -13.10816, -13.10832, -13.10875, -13.10911, -13.10836, 
    -13.1092, -13.10605, -13.10772, -13.10515, -13.10592, -13.10647, 
    -13.10625, -13.10747, -13.10775, -13.10889, -13.10831, -13.11186, 
    -13.11028, -13.11476, -13.11349, -13.10517, -13.10557, -13.10692, 
    -13.10629, -13.10813, -13.10858, -13.10894, -13.10941, -13.10946, 
    -13.10974, -13.10929, -13.10973, -13.10807, -13.1088, -13.10678, 
    -13.10727, -13.10705, -13.1068, -13.10757, -13.10837, -13.10841, 
    -13.10865, -13.10933, -13.10814, -13.11203, -13.10958, -13.106, 
    -13.10673, -13.10686, -13.10658, -13.10853, -13.10782, -13.10974, 
    -13.10922, -13.11007, -13.10965, -13.10958, -13.10904, -13.1087, 
    -13.10785, -13.10716, -13.10662, -13.10675, -13.10734, -13.10842, 
    -13.10946, -13.10923, -13.11001, -13.108, -13.10882, -13.1085, -13.10936, 
    -13.1075, -13.10902, -13.1071, -13.10727, -13.10781, -13.10887, 
    -13.10913, -13.10938, -13.10923, -13.10845, -13.10834, -13.1078, 
    -13.10764, -13.10724, -13.10689, -13.1072, -13.10752, -13.10846, 
    -13.1093, -13.11022, -13.11046, -13.1115, -13.11062, -13.11204, 
    -13.11079, -13.11298, -13.10914, -13.1108, -13.10784, -13.10816, 
    -13.10872, -13.11006, -13.10935, -13.11019, -13.10833, -13.10735, 
    -13.10712, -13.10665, -13.10713, -13.10709, -13.10755, -13.1074, 
    -13.1085, -13.10791, -13.10958, -13.11018, -13.11194, -13.11301, 
    -13.11414, -13.11463, -13.11478, -13.11484 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531 ;

 FSRND =
  0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505 ;

 FSRVD =
  0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.809097e-14, 2.821622e-14, 2.819179e-14, 2.829291e-14, 2.823676e-14, 
    2.830296e-14, 2.81162e-14, 2.822105e-14, 2.815406e-14, 2.810199e-14, 
    2.848918e-14, 2.829722e-14, 2.868855e-14, 2.856595e-14, 2.887388e-14, 
    2.866944e-14, 2.89151e-14, 2.886786e-14, 2.90098e-14, 2.896908e-14, 
    2.915086e-14, 2.902851e-14, 2.924503e-14, 2.912156e-14, 2.914086e-14, 
    2.902437e-14, 2.833595e-14, 2.846547e-14, 2.832824e-14, 2.834671e-14, 
    2.833838e-14, 2.823783e-14, 2.818724e-14, 2.808113e-14, 2.810034e-14, 
    2.817823e-14, 2.835483e-14, 2.829477e-14, 2.844593e-14, 2.844252e-14, 
    2.861098e-14, 2.853498e-14, 2.88184e-14, 2.873774e-14, 2.897075e-14, 
    2.891209e-14, 2.896796e-14, 2.895097e-14, 2.896811e-14, 2.888214e-14, 
    2.891892e-14, 2.884328e-14, 2.854952e-14, 2.863594e-14, 2.837823e-14, 
    2.822353e-14, 2.812071e-14, 2.804786e-14, 2.80581e-14, 2.807775e-14, 
    2.817864e-14, 2.827349e-14, 2.834585e-14, 2.839425e-14, 2.844195e-14, 
    2.858668e-14, 2.866317e-14, 2.883468e-14, 2.880365e-14, 2.885613e-14, 
    2.890623e-14, 2.899042e-14, 2.897654e-14, 2.901363e-14, 2.885457e-14, 
    2.896027e-14, 2.878577e-14, 2.883348e-14, 2.845539e-14, 2.831106e-14, 
    2.824994e-14, 2.819627e-14, 2.806601e-14, 2.815595e-14, 2.812046e-14, 
    2.820474e-14, 2.825836e-14, 2.823179e-14, 2.839555e-14, 2.833183e-14, 
    2.866767e-14, 2.852292e-14, 2.890042e-14, 2.880996e-14, 2.892201e-14, 
    2.886481e-14, 2.896281e-14, 2.887456e-14, 2.902739e-14, 2.906072e-14, 
    2.90379e-14, 2.912532e-14, 2.886952e-14, 2.896773e-14, 2.82312e-14, 
    2.823553e-14, 2.825565e-14, 2.816708e-14, 2.816164e-14, 2.808047e-14, 
    2.815261e-14, 2.818338e-14, 2.826139e-14, 2.830757e-14, 2.835147e-14, 
    2.844812e-14, 2.855611e-14, 2.870719e-14, 2.881579e-14, 2.88886e-14, 
    2.88439e-14, 2.888332e-14, 2.883921e-14, 2.88185e-14, 2.904817e-14, 
    2.891918e-14, 2.911267e-14, 2.910196e-14, 2.901433e-14, 2.910309e-14, 
    2.823852e-14, 2.821358e-14, 2.812721e-14, 2.819475e-14, 2.807158e-14, 
    2.814053e-14, 2.818016e-14, 2.833317e-14, 2.836674e-14, 2.839796e-14, 
    2.845957e-14, 2.853869e-14, 2.867764e-14, 2.879857e-14, 2.890903e-14, 
    2.89009e-14, 2.890374e-14, 2.892841e-14, 2.886723e-14, 2.89384e-14, 
    2.895034e-14, 2.891907e-14, 2.910045e-14, 2.90486e-14, 2.910163e-14, 
    2.906782e-14, 2.822164e-14, 2.82635e-14, 2.824083e-14, 2.828342e-14, 
    2.825338e-14, 2.838682e-14, 2.842682e-14, 2.861415e-14, 2.853714e-14, 
    2.865961e-14, 2.854951e-14, 2.856902e-14, 2.866361e-14, 2.855537e-14, 
    2.879187e-14, 2.863153e-14, 2.892934e-14, 2.876919e-14, 2.893933e-14, 
    2.890835e-14, 2.895953e-14, 2.900544e-14, 2.906311e-14, 2.916972e-14, 
    2.914496e-14, 2.923413e-14, 2.832594e-14, 2.83803e-14, 2.837546e-14, 
    2.843234e-14, 2.847443e-14, 2.856571e-14, 2.871221e-14, 2.865704e-14, 
    2.875819e-14, 2.877853e-14, 2.862474e-14, 2.871916e-14, 2.841643e-14, 
    2.84653e-14, 2.843614e-14, 2.832987e-14, 2.866959e-14, 2.849514e-14, 
    2.881729e-14, 2.872266e-14, 2.899883e-14, 2.886146e-14, 2.913136e-14, 
    2.924698e-14, 2.935564e-14, 2.94829e-14, 2.840992e-14, 2.837292e-14, 
    2.843905e-14, 2.853071e-14, 2.861563e-14, 2.872874e-14, 2.874026e-14, 
    2.876143e-14, 2.881629e-14, 2.886249e-14, 2.876811e-14, 2.8874e-14, 
    2.84767e-14, 2.868471e-14, 2.835865e-14, 2.845682e-14, 2.852494e-14, 
    2.8495e-14, 2.865041e-14, 2.868704e-14, 2.883612e-14, 2.8759e-14, 
    2.92184e-14, 2.901501e-14, 2.957969e-14, 2.942175e-14, 2.835999e-14, 
    2.840967e-14, 2.858288e-14, 2.850043e-14, 2.87362e-14, 2.879431e-14, 
    2.884148e-14, 2.890193e-14, 2.890837e-14, 2.89442e-14, 2.888545e-14, 
    2.894181e-14, 2.872871e-14, 2.882388e-14, 2.856275e-14, 2.862625e-14, 
    2.859699e-14, 2.856491e-14, 2.86638e-14, 2.876933e-14, 2.877149e-14, 
    2.880531e-14, 2.890086e-14, 2.873669e-14, 2.92447e-14, 2.893087e-14, 
    2.846389e-14, 2.85598e-14, 2.85734e-14, 2.853624e-14, 2.878842e-14, 
    2.8697e-14, 2.894331e-14, 2.887665e-14, 2.898578e-14, 2.893154e-14, 
    2.892351e-14, 2.885385e-14, 2.881046e-14, 2.8701e-14, 2.861192e-14, 
    2.854133e-14, 2.855768e-14, 2.863524e-14, 2.87757e-14, 2.890868e-14, 
    2.887952e-14, 2.897716e-14, 2.871858e-14, 2.882699e-14, 2.878505e-14, 
    2.889428e-14, 2.865549e-14, 2.885945e-14, 2.860339e-14, 2.862577e-14, 
    2.869511e-14, 2.883476e-14, 2.886552e-14, 2.889856e-14, 2.887811e-14, 
    2.877944e-14, 2.876322e-14, 2.869324e-14, 2.867394e-14, 2.862066e-14, 
    2.857653e-14, 2.861682e-14, 2.865909e-14, 2.877926e-14, 2.888761e-14, 
    2.900579e-14, 2.90347e-14, 2.917306e-14, 2.906047e-14, 2.924633e-14, 
    2.908839e-14, 2.936175e-14, 2.887111e-14, 2.908413e-14, 2.869825e-14, 
    2.873973e-14, 2.88149e-14, 2.898726e-14, 2.889407e-14, 2.9003e-14, 
    2.876256e-14, 2.863799e-14, 2.860567e-14, 2.85456e-14, 2.8607e-14, 
    2.860201e-14, 2.866081e-14, 2.864186e-14, 2.878318e-14, 2.870724e-14, 
    2.892299e-14, 2.900183e-14, 2.922452e-14, 2.936117e-14, 2.950029e-14, 
    2.956173e-14, 2.958043e-14, 2.958823e-14 ;

 F_DENIT_vr =
  1.604023e-12, 1.611175e-12, 1.609781e-12, 1.615554e-12, 1.612348e-12, 
    1.616128e-12, 1.605464e-12, 1.611451e-12, 1.607626e-12, 1.604653e-12, 
    1.626762e-12, 1.6158e-12, 1.638146e-12, 1.631145e-12, 1.648729e-12, 
    1.637055e-12, 1.651082e-12, 1.648384e-12, 1.65649e-12, 1.654164e-12, 
    1.664544e-12, 1.657558e-12, 1.669921e-12, 1.662871e-12, 1.663973e-12, 
    1.657321e-12, 1.618012e-12, 1.625408e-12, 1.617572e-12, 1.618626e-12, 
    1.618151e-12, 1.61241e-12, 1.60952e-12, 1.603462e-12, 1.604558e-12, 
    1.609006e-12, 1.61909e-12, 1.615661e-12, 1.624292e-12, 1.624097e-12, 
    1.633717e-12, 1.629377e-12, 1.645561e-12, 1.640955e-12, 1.65426e-12, 
    1.65091e-12, 1.6541e-12, 1.65313e-12, 1.654109e-12, 1.6492e-12, 
    1.6513e-12, 1.646981e-12, 1.630207e-12, 1.635142e-12, 1.620426e-12, 
    1.611593e-12, 1.605721e-12, 1.601562e-12, 1.602147e-12, 1.603269e-12, 
    1.609029e-12, 1.614446e-12, 1.618578e-12, 1.621341e-12, 1.624065e-12, 
    1.632329e-12, 1.636697e-12, 1.64649e-12, 1.644718e-12, 1.647715e-12, 
    1.650576e-12, 1.655383e-12, 1.65459e-12, 1.656709e-12, 1.647626e-12, 
    1.653661e-12, 1.643697e-12, 1.646422e-12, 1.624832e-12, 1.616591e-12, 
    1.613101e-12, 1.610036e-12, 1.602598e-12, 1.607734e-12, 1.605707e-12, 
    1.61052e-12, 1.613582e-12, 1.612064e-12, 1.621415e-12, 1.617777e-12, 
    1.636953e-12, 1.628688e-12, 1.650244e-12, 1.645078e-12, 1.651477e-12, 
    1.64821e-12, 1.653807e-12, 1.648767e-12, 1.657494e-12, 1.659397e-12, 
    1.658094e-12, 1.663086e-12, 1.648479e-12, 1.654087e-12, 1.612031e-12, 
    1.612278e-12, 1.613427e-12, 1.608369e-12, 1.608059e-12, 1.603424e-12, 
    1.607543e-12, 1.6093e-12, 1.613755e-12, 1.616392e-12, 1.618898e-12, 
    1.624417e-12, 1.630583e-12, 1.63921e-12, 1.645411e-12, 1.649569e-12, 
    1.647017e-12, 1.649267e-12, 1.646749e-12, 1.645566e-12, 1.658681e-12, 
    1.651315e-12, 1.662364e-12, 1.661752e-12, 1.656748e-12, 1.661817e-12, 
    1.612449e-12, 1.611025e-12, 1.606093e-12, 1.609949e-12, 1.602916e-12, 
    1.606853e-12, 1.609116e-12, 1.617853e-12, 1.61977e-12, 1.621553e-12, 
    1.625071e-12, 1.629588e-12, 1.637523e-12, 1.644428e-12, 1.650736e-12, 
    1.650271e-12, 1.650433e-12, 1.651842e-12, 1.648349e-12, 1.652413e-12, 
    1.653094e-12, 1.651309e-12, 1.661666e-12, 1.658705e-12, 1.661733e-12, 
    1.659803e-12, 1.611485e-12, 1.613875e-12, 1.612581e-12, 1.615012e-12, 
    1.613297e-12, 1.620917e-12, 1.6232e-12, 1.633897e-12, 1.6295e-12, 
    1.636493e-12, 1.630206e-12, 1.631321e-12, 1.636722e-12, 1.630542e-12, 
    1.644045e-12, 1.63489e-12, 1.651895e-12, 1.64275e-12, 1.652466e-12, 
    1.650697e-12, 1.653619e-12, 1.65624e-12, 1.659533e-12, 1.665621e-12, 
    1.664208e-12, 1.669299e-12, 1.61744e-12, 1.620544e-12, 1.620268e-12, 
    1.623516e-12, 1.625919e-12, 1.631131e-12, 1.639497e-12, 1.636347e-12, 
    1.642123e-12, 1.643284e-12, 1.634502e-12, 1.639894e-12, 1.622608e-12, 
    1.625398e-12, 1.623733e-12, 1.617665e-12, 1.637063e-12, 1.627102e-12, 
    1.645497e-12, 1.640094e-12, 1.655863e-12, 1.648019e-12, 1.663431e-12, 
    1.670033e-12, 1.676237e-12, 1.683504e-12, 1.622236e-12, 1.620123e-12, 
    1.623899e-12, 1.629133e-12, 1.633982e-12, 1.64044e-12, 1.641098e-12, 
    1.642307e-12, 1.64544e-12, 1.648078e-12, 1.642689e-12, 1.648735e-12, 
    1.626049e-12, 1.637927e-12, 1.619309e-12, 1.624914e-12, 1.628804e-12, 
    1.627094e-12, 1.635968e-12, 1.63806e-12, 1.646572e-12, 1.642169e-12, 
    1.668401e-12, 1.656787e-12, 1.689031e-12, 1.680013e-12, 1.619384e-12, 
    1.622222e-12, 1.632112e-12, 1.627404e-12, 1.640866e-12, 1.644185e-12, 
    1.646878e-12, 1.65033e-12, 1.650698e-12, 1.652743e-12, 1.649389e-12, 
    1.652607e-12, 1.640439e-12, 1.645874e-12, 1.630963e-12, 1.634589e-12, 
    1.632918e-12, 1.631086e-12, 1.636733e-12, 1.642758e-12, 1.642882e-12, 
    1.644813e-12, 1.650269e-12, 1.640895e-12, 1.669902e-12, 1.651983e-12, 
    1.625318e-12, 1.630794e-12, 1.63157e-12, 1.629449e-12, 1.643848e-12, 
    1.638628e-12, 1.652693e-12, 1.648886e-12, 1.655118e-12, 1.652021e-12, 
    1.651562e-12, 1.647585e-12, 1.645107e-12, 1.638857e-12, 1.63377e-12, 
    1.629739e-12, 1.630673e-12, 1.635102e-12, 1.643122e-12, 1.650716e-12, 
    1.64905e-12, 1.654626e-12, 1.639861e-12, 1.646051e-12, 1.643656e-12, 
    1.649893e-12, 1.636258e-12, 1.647904e-12, 1.633283e-12, 1.634561e-12, 
    1.63852e-12, 1.646495e-12, 1.648251e-12, 1.650137e-12, 1.64897e-12, 
    1.643336e-12, 1.642409e-12, 1.638414e-12, 1.637311e-12, 1.634269e-12, 
    1.63175e-12, 1.63405e-12, 1.636464e-12, 1.643325e-12, 1.649513e-12, 
    1.656261e-12, 1.657911e-12, 1.665812e-12, 1.659383e-12, 1.669996e-12, 
    1.660977e-12, 1.676586e-12, 1.64857e-12, 1.660734e-12, 1.6387e-12, 
    1.641068e-12, 1.64536e-12, 1.655203e-12, 1.649881e-12, 1.656101e-12, 
    1.642372e-12, 1.635259e-12, 1.633414e-12, 1.629983e-12, 1.633489e-12, 
    1.633204e-12, 1.636562e-12, 1.63548e-12, 1.643549e-12, 1.639213e-12, 
    1.651533e-12, 1.656034e-12, 1.66875e-12, 1.676553e-12, 1.684497e-12, 
    1.688006e-12, 1.689073e-12, 1.689519e-12,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  7.54986e-16, 7.557574e-16, 7.556063e-16, 7.562241e-16, 7.558807e-16, 
    7.562836e-16, 7.551389e-16, 7.557841e-16, 7.553715e-16, 7.55049e-16, 
    7.574024e-16, 7.562462e-16, 7.585715e-16, 7.578514e-16, 7.596374e-16, 
    7.584596e-16, 7.598709e-16, 7.596001e-16, 7.60403e-16, 7.60173e-16, 
    7.611905e-16, 7.605066e-16, 7.617063e-16, 7.610258e-16, 7.611327e-16, 
    7.604811e-16, 7.564834e-16, 7.572652e-16, 7.564359e-16, 7.565481e-16, 
    7.564966e-16, 7.558856e-16, 7.55577e-16, 7.549192e-16, 7.550377e-16, 
    7.555193e-16, 7.565936e-16, 7.562285e-16, 7.571374e-16, 7.571171e-16, 
    7.581141e-16, 7.576662e-16, 7.593167e-16, 7.588507e-16, 7.601818e-16, 
    7.598493e-16, 7.601653e-16, 7.600683e-16, 7.601646e-16, 7.596777e-16, 
    7.598856e-16, 7.594546e-16, 7.577585e-16, 7.582661e-16, 7.567368e-16, 
    7.558001e-16, 7.551649e-16, 7.547125e-16, 7.547753e-16, 7.54898e-16, 
    7.555208e-16, 7.560988e-16, 7.565368e-16, 7.568274e-16, 7.571123e-16, 
    7.579741e-16, 7.584199e-16, 7.594097e-16, 7.592303e-16, 7.595311e-16, 
    7.598153e-16, 7.60291e-16, 7.602122e-16, 7.604205e-16, 7.595185e-16, 
    7.601198e-16, 7.591226e-16, 7.593971e-16, 7.572029e-16, 7.563296e-16, 
    7.559604e-16, 7.556296e-16, 7.548243e-16, 7.553814e-16, 7.551617e-16, 
    7.556787e-16, 7.560063e-16, 7.55843e-16, 7.568346e-16, 7.564502e-16, 
    7.584452e-16, 7.575939e-16, 7.59783e-16, 7.592655e-16, 7.599041e-16, 
    7.595785e-16, 7.601345e-16, 7.596332e-16, 7.604964e-16, 7.606838e-16, 
    7.605546e-16, 7.610415e-16, 7.596014e-16, 7.601594e-16, 7.558427e-16, 
    7.558693e-16, 7.559911e-16, 7.554493e-16, 7.554153e-16, 7.549122e-16, 
    7.553577e-16, 7.555475e-16, 7.560229e-16, 7.563031e-16, 7.565679e-16, 
    7.57148e-16, 7.577893e-16, 7.586727e-16, 7.592984e-16, 7.597134e-16, 
    7.594579e-16, 7.596823e-16, 7.594303e-16, 7.593106e-16, 7.606122e-16, 
    7.598854e-16, 7.609699e-16, 7.609103e-16, 7.604207e-16, 7.609151e-16, 
    7.558865e-16, 7.55733e-16, 7.552023e-16, 7.556167e-16, 7.548559e-16, 
    7.552834e-16, 7.555274e-16, 7.564587e-16, 7.566592e-16, 7.568475e-16, 
    7.572151e-16, 7.576843e-16, 7.585002e-16, 7.591989e-16, 7.598289e-16, 
    7.597818e-16, 7.597978e-16, 7.599374e-16, 7.595892e-16, 7.59993e-16, 
    7.600603e-16, 7.598828e-16, 7.609004e-16, 7.606113e-16, 7.609064e-16, 
    7.607171e-16, 7.557817e-16, 7.560366e-16, 7.558977e-16, 7.561575e-16, 
    7.559738e-16, 7.567824e-16, 7.570219e-16, 7.581309e-16, 7.576754e-16, 
    7.583956e-16, 7.577471e-16, 7.578628e-16, 7.584195e-16, 7.577801e-16, 
    7.591598e-16, 7.582293e-16, 7.599421e-16, 7.590286e-16, 7.599976e-16, 
    7.598208e-16, 7.6011e-16, 7.603694e-16, 7.60691e-16, 7.61284e-16, 
    7.611456e-16, 7.616367e-16, 7.564149e-16, 7.567428e-16, 7.567124e-16, 
    7.57053e-16, 7.573038e-16, 7.578442e-16, 7.58701e-16, 7.583786e-16, 
    7.58965e-16, 7.590828e-16, 7.581878e-16, 7.587394e-16, 7.569542e-16, 
    7.572464e-16, 7.570708e-16, 7.564314e-16, 7.58449e-16, 7.574218e-16, 
    7.593011e-16, 7.587544e-16, 7.603307e-16, 7.595534e-16, 7.610698e-16, 
    7.61709e-16, 7.622967e-16, 7.629814e-16, 7.569194e-16, 7.566959e-16, 
    7.570918e-16, 7.576388e-16, 7.581367e-16, 7.58796e-16, 7.588615e-16, 
    7.589833e-16, 7.59298e-16, 7.595626e-16, 7.590217e-16, 7.596267e-16, 
    7.57316e-16, 7.585365e-16, 7.56604e-16, 7.571942e-16, 7.575969e-16, 
    7.574188e-16, 7.583329e-16, 7.585459e-16, 7.594066e-16, 7.589623e-16, 
    7.615512e-16, 7.604209e-16, 7.634918e-16, 7.626528e-16, 7.566175e-16, 
    7.569153e-16, 7.579446e-16, 7.574567e-16, 7.588372e-16, 7.59173e-16, 
    7.594419e-16, 7.597876e-16, 7.598224e-16, 7.60026e-16, 7.596909e-16, 
    7.600111e-16, 7.587903e-16, 7.593385e-16, 7.578191e-16, 7.581922e-16, 
    7.580197e-16, 7.578301e-16, 7.584094e-16, 7.590232e-16, 7.590334e-16, 
    7.592281e-16, 7.59779e-16, 7.588306e-16, 7.616965e-16, 7.599468e-16, 
    7.572388e-16, 7.578088e-16, 7.578866e-16, 7.57667e-16, 7.591376e-16, 
    7.58609e-16, 7.600207e-16, 7.596411e-16, 7.602588e-16, 7.599526e-16, 
    7.59906e-16, 7.595095e-16, 7.592601e-16, 7.586285e-16, 7.581072e-16, 
    7.576909e-16, 7.577864e-16, 7.582431e-16, 7.590581e-16, 7.598185e-16, 
    7.596523e-16, 7.602038e-16, 7.587247e-16, 7.593506e-16, 7.591088e-16, 
    7.597331e-16, 7.583678e-16, 7.595503e-16, 7.580615e-16, 7.581921e-16, 
    7.585965e-16, 7.59404e-16, 7.595766e-16, 7.597656e-16, 7.596473e-16, 
    7.590832e-16, 7.589885e-16, 7.585819e-16, 7.584695e-16, 7.581574e-16, 
    7.578971e-16, 7.581343e-16, 7.583812e-16, 7.590775e-16, 7.596978e-16, 
    7.603652e-16, 7.605266e-16, 7.612988e-16, 7.606726e-16, 7.617032e-16, 
    7.608313e-16, 7.623279e-16, 7.596133e-16, 7.608148e-16, 7.586144e-16, 
    7.588541e-16, 7.592887e-16, 7.602683e-16, 7.597382e-16, 7.603558e-16, 
    7.589842e-16, 7.582609e-16, 7.580692e-16, 7.577157e-16, 7.58076e-16, 
    7.580467e-16, 7.583902e-16, 7.582786e-16, 7.590985e-16, 7.586592e-16, 
    7.598968e-16, 7.603427e-16, 7.615787e-16, 7.623227e-16, 7.630666e-16, 
    7.633915e-16, 7.634899e-16, 7.635304e-16 ;

 F_N2O_NIT =
  2.408225e-14, 2.42901e-14, 2.424961e-14, 2.441779e-14, 2.432442e-14, 
    2.443464e-14, 2.41243e-14, 2.429835e-14, 2.418716e-14, 2.41009e-14, 
    2.474585e-14, 2.442528e-14, 2.50811e-14, 2.487497e-14, 2.539442e-14, 
    2.504896e-14, 2.546437e-14, 2.53844e-14, 2.562544e-14, 2.555626e-14, 
    2.586586e-14, 2.565739e-14, 2.602709e-14, 2.581599e-14, 2.584895e-14, 
    2.565052e-14, 2.448963e-14, 2.470584e-14, 2.447685e-14, 2.450761e-14, 
    2.44938e-14, 2.432634e-14, 2.424217e-14, 2.406637e-14, 2.409824e-14, 
    2.422737e-14, 2.452143e-14, 2.44214e-14, 2.467389e-14, 2.466818e-14, 
    2.495082e-14, 2.482317e-14, 2.530072e-14, 2.516451e-14, 2.555914e-14, 
    2.54596e-14, 2.555446e-14, 2.552567e-14, 2.555483e-14, 2.540892e-14, 
    2.547137e-14, 2.534317e-14, 2.484708e-14, 2.499237e-14, 2.456034e-14, 
    2.430244e-14, 2.413191e-14, 2.401128e-14, 2.402831e-14, 2.40608e-14, 
    2.422813e-14, 2.438598e-14, 2.450664e-14, 2.458752e-14, 2.466735e-14, 
    2.490981e-14, 2.503863e-14, 2.532831e-14, 2.527589e-14, 2.536471e-14, 
    2.54497e-14, 2.559273e-14, 2.556916e-14, 2.563227e-14, 2.536235e-14, 
    2.554158e-14, 2.524605e-14, 2.53267e-14, 2.468912e-14, 2.444838e-14, 
    2.434644e-14, 2.425737e-14, 2.404141e-14, 2.419044e-14, 2.413163e-14, 
    2.427165e-14, 2.436084e-14, 2.43167e-14, 2.458973e-14, 2.448339e-14, 
    2.504627e-14, 2.480301e-14, 2.543978e-14, 2.528664e-14, 2.547655e-14, 
    2.537955e-14, 2.554587e-14, 2.539615e-14, 2.565578e-14, 2.57125e-14, 
    2.567373e-14, 2.58228e-14, 2.538785e-14, 2.555444e-14, 2.431548e-14, 
    2.432267e-14, 2.43562e-14, 2.420898e-14, 2.419998e-14, 2.406549e-14, 
    2.418513e-14, 2.423618e-14, 2.4366e-14, 2.444296e-14, 2.451624e-14, 
    2.467775e-14, 2.485877e-14, 2.511305e-14, 2.529655e-14, 2.541994e-14, 
    2.534424e-14, 2.541106e-14, 2.533636e-14, 2.530138e-14, 2.569123e-14, 
    2.547195e-14, 2.580132e-14, 2.578304e-14, 2.563376e-14, 2.578509e-14, 
    2.432772e-14, 2.428632e-14, 2.41429e-14, 2.42551e-14, 2.405086e-14, 
    2.416507e-14, 2.423087e-14, 2.448561e-14, 2.454176e-14, 2.459389e-14, 
    2.469701e-14, 2.482968e-14, 2.506331e-14, 2.526749e-14, 2.545464e-14, 
    2.54409e-14, 2.544573e-14, 2.548763e-14, 2.538391e-14, 2.550467e-14, 
    2.552497e-14, 2.547191e-14, 2.578058e-14, 2.56922e-14, 2.578264e-14, 
    2.572507e-14, 2.429977e-14, 2.436946e-14, 2.433178e-14, 2.440265e-14, 
    2.435271e-14, 2.457515e-14, 2.464204e-14, 2.49563e-14, 2.482707e-14, 
    2.503289e-14, 2.484793e-14, 2.488065e-14, 2.503962e-14, 2.48579e-14, 
    2.525621e-14, 2.498581e-14, 2.548925e-14, 2.521795e-14, 2.55063e-14, 
    2.545381e-14, 2.554074e-14, 2.561873e-14, 2.571702e-14, 2.589889e-14, 
    2.585671e-14, 2.600919e-14, 2.447354e-14, 2.456428e-14, 2.455628e-14, 
    2.46514e-14, 2.472188e-14, 2.487499e-14, 2.512158e-14, 2.50287e-14, 
    2.519934e-14, 2.523367e-14, 2.497447e-14, 2.513345e-14, 2.462508e-14, 
    2.470685e-14, 2.465814e-14, 2.448065e-14, 2.505007e-14, 2.4757e-14, 
    2.529956e-14, 2.513975e-14, 2.56076e-14, 2.537437e-14, 2.583351e-14, 
    2.60311e-14, 2.621775e-14, 2.643677e-14, 2.461387e-14, 2.455212e-14, 
    2.466272e-14, 2.481618e-14, 2.495899e-14, 2.514952e-14, 2.516905e-14, 
    2.520483e-14, 2.529766e-14, 2.537585e-14, 2.521616e-14, 2.539546e-14, 
    2.472584e-14, 2.507559e-14, 2.452877e-14, 2.469278e-14, 2.480709e-14, 
    2.475691e-14, 2.501806e-14, 2.507982e-14, 2.53316e-14, 2.520128e-14, 
    2.598226e-14, 2.563521e-14, 2.660415e-14, 2.63315e-14, 2.453057e-14, 
    2.461364e-14, 2.490393e-14, 2.476559e-14, 2.516225e-14, 2.526039e-14, 
    2.534031e-14, 2.544267e-14, 2.545373e-14, 2.551449e-14, 2.541495e-14, 
    2.551055e-14, 2.51499e-14, 2.531073e-14, 2.487062e-14, 2.497738e-14, 
    2.492823e-14, 2.487438e-14, 2.504075e-14, 2.521864e-14, 2.522244e-14, 
    2.527961e-14, 2.544112e-14, 2.516382e-14, 2.602723e-14, 2.549224e-14, 
    2.47044e-14, 2.486515e-14, 2.488814e-14, 2.482578e-14, 2.525054e-14, 
    2.50962e-14, 2.551301e-14, 2.54e-14, 2.558528e-14, 2.549313e-14, 
    2.547958e-14, 2.53615e-14, 2.528812e-14, 2.510325e-14, 2.495333e-14, 
    2.483479e-14, 2.486232e-14, 2.499263e-14, 2.522953e-14, 2.54547e-14, 
    2.540529e-14, 2.557115e-14, 2.513333e-14, 2.531644e-14, 2.524558e-14, 
    2.543054e-14, 2.502623e-14, 2.537038e-14, 2.493865e-14, 2.497634e-14, 
    2.509314e-14, 2.532893e-14, 2.538123e-14, 2.543716e-14, 2.540264e-14, 
    2.523558e-14, 2.520826e-14, 2.509028e-14, 2.505775e-14, 2.496811e-14, 
    2.489402e-14, 2.496171e-14, 2.503289e-14, 2.523563e-14, 2.541905e-14, 
    2.561981e-14, 2.566907e-14, 2.590492e-14, 2.571285e-14, 2.603021e-14, 
    2.576027e-14, 2.622846e-14, 2.539038e-14, 2.57524e-14, 2.509846e-14, 
    2.516848e-14, 2.529541e-14, 2.558776e-14, 2.54297e-14, 2.561459e-14, 
    2.520718e-14, 2.499714e-14, 2.494294e-14, 2.484198e-14, 2.494524e-14, 
    2.493683e-14, 2.503583e-14, 2.500399e-14, 2.524236e-14, 2.511417e-14, 
    2.547921e-14, 2.56131e-14, 2.599316e-14, 2.622759e-14, 2.646733e-14, 
    2.657353e-14, 2.66059e-14, 2.661943e-14 ;

 F_NIT =
  4.013708e-11, 4.04835e-11, 4.041602e-11, 4.069631e-11, 4.05407e-11, 
    4.07244e-11, 4.020716e-11, 4.049725e-11, 4.031193e-11, 4.016816e-11, 
    4.124308e-11, 4.07088e-11, 4.180183e-11, 4.145828e-11, 4.232403e-11, 
    4.174826e-11, 4.244061e-11, 4.230734e-11, 4.270907e-11, 4.259377e-11, 
    4.310976e-11, 4.276232e-11, 4.337848e-11, 4.302664e-11, 4.308158e-11, 
    4.275086e-11, 4.081606e-11, 4.11764e-11, 4.079475e-11, 4.084602e-11, 
    4.0823e-11, 4.054389e-11, 4.040362e-11, 4.011063e-11, 4.016373e-11, 
    4.037896e-11, 4.086906e-11, 4.070233e-11, 4.112315e-11, 4.111363e-11, 
    4.15847e-11, 4.137196e-11, 4.216787e-11, 4.194085e-11, 4.259857e-11, 
    4.243266e-11, 4.259077e-11, 4.254279e-11, 4.259138e-11, 4.234819e-11, 
    4.245229e-11, 4.223862e-11, 4.141181e-11, 4.165395e-11, 4.09339e-11, 
    4.050408e-11, 4.021985e-11, 4.00188e-11, 4.004718e-11, 4.010134e-11, 
    4.038021e-11, 4.06433e-11, 4.08444e-11, 4.09792e-11, 4.111224e-11, 
    4.151636e-11, 4.173105e-11, 4.221384e-11, 4.212649e-11, 4.227451e-11, 
    4.241617e-11, 4.265455e-11, 4.261526e-11, 4.272046e-11, 4.227058e-11, 
    4.25693e-11, 4.207674e-11, 4.221117e-11, 4.114853e-11, 4.074729e-11, 
    4.057739e-11, 4.042895e-11, 4.006902e-11, 4.03174e-11, 4.021939e-11, 
    4.045275e-11, 4.060139e-11, 4.052783e-11, 4.098288e-11, 4.080565e-11, 
    4.174378e-11, 4.133835e-11, 4.239964e-11, 4.21444e-11, 4.246092e-11, 
    4.229925e-11, 4.257645e-11, 4.232692e-11, 4.275963e-11, 4.285416e-11, 
    4.278954e-11, 4.3038e-11, 4.231309e-11, 4.259073e-11, 4.052579e-11, 
    4.053779e-11, 4.059367e-11, 4.034829e-11, 4.03333e-11, 4.010915e-11, 
    4.030856e-11, 4.039363e-11, 4.061e-11, 4.073827e-11, 4.086039e-11, 
    4.112958e-11, 4.143129e-11, 4.185508e-11, 4.216092e-11, 4.236657e-11, 
    4.22404e-11, 4.235177e-11, 4.222727e-11, 4.216897e-11, 4.281872e-11, 
    4.245325e-11, 4.30022e-11, 4.297173e-11, 4.272293e-11, 4.297515e-11, 
    4.05462e-11, 4.04772e-11, 4.023816e-11, 4.042516e-11, 4.008477e-11, 
    4.027512e-11, 4.038479e-11, 4.080936e-11, 4.090293e-11, 4.098982e-11, 
    4.116169e-11, 4.13828e-11, 4.177218e-11, 4.211249e-11, 4.24244e-11, 
    4.24015e-11, 4.240956e-11, 4.247938e-11, 4.230651e-11, 4.250779e-11, 
    4.254161e-11, 4.245319e-11, 4.296764e-11, 4.282033e-11, 4.297107e-11, 
    4.287511e-11, 4.049962e-11, 4.061576e-11, 4.055297e-11, 4.067108e-11, 
    4.058785e-11, 4.095858e-11, 4.107007e-11, 4.159383e-11, 4.137844e-11, 
    4.172148e-11, 4.141321e-11, 4.146775e-11, 4.17327e-11, 4.142982e-11, 
    4.209368e-11, 4.164302e-11, 4.248209e-11, 4.202992e-11, 4.25105e-11, 
    4.242301e-11, 4.25679e-11, 4.269789e-11, 4.286169e-11, 4.316482e-11, 
    4.309452e-11, 4.334865e-11, 4.078923e-11, 4.094046e-11, 4.092713e-11, 
    4.108568e-11, 4.120313e-11, 4.145832e-11, 4.186931e-11, 4.17145e-11, 
    4.19989e-11, 4.205612e-11, 4.162412e-11, 4.188909e-11, 4.104179e-11, 
    4.117808e-11, 4.10969e-11, 4.080108e-11, 4.175012e-11, 4.126166e-11, 
    4.216593e-11, 4.189959e-11, 4.267933e-11, 4.229062e-11, 4.305585e-11, 
    4.338517e-11, 4.369625e-11, 4.406129e-11, 4.102312e-11, 4.09202e-11, 
    4.110454e-11, 4.136031e-11, 4.159832e-11, 4.191586e-11, 4.194841e-11, 
    4.200806e-11, 4.216276e-11, 4.229308e-11, 4.202692e-11, 4.232576e-11, 
    4.120973e-11, 4.179266e-11, 4.088128e-11, 4.115464e-11, 4.134515e-11, 
    4.126151e-11, 4.169677e-11, 4.17997e-11, 4.221933e-11, 4.200213e-11, 
    4.330376e-11, 4.272535e-11, 4.434026e-11, 4.388584e-11, 4.088428e-11, 
    4.102274e-11, 4.150654e-11, 4.127598e-11, 4.193709e-11, 4.210066e-11, 
    4.223385e-11, 4.240445e-11, 4.242288e-11, 4.252415e-11, 4.235826e-11, 
    4.251758e-11, 4.191649e-11, 4.218455e-11, 4.145104e-11, 4.162896e-11, 
    4.154705e-11, 4.145731e-11, 4.173459e-11, 4.203106e-11, 4.203739e-11, 
    4.213269e-11, 4.240186e-11, 4.19397e-11, 4.337871e-11, 4.248706e-11, 
    4.1174e-11, 4.144191e-11, 4.148023e-11, 4.13763e-11, 4.208423e-11, 
    4.1827e-11, 4.252168e-11, 4.233334e-11, 4.264214e-11, 4.248855e-11, 
    4.246596e-11, 4.226916e-11, 4.214687e-11, 4.183875e-11, 4.158889e-11, 
    4.139131e-11, 4.14372e-11, 4.165439e-11, 4.204922e-11, 4.24245e-11, 
    4.234214e-11, 4.261858e-11, 4.188888e-11, 4.219407e-11, 4.207597e-11, 
    4.238424e-11, 4.171038e-11, 4.228396e-11, 4.156442e-11, 4.162724e-11, 
    4.182189e-11, 4.221488e-11, 4.230205e-11, 4.239527e-11, 4.233773e-11, 
    4.20593e-11, 4.201376e-11, 4.181713e-11, 4.176292e-11, 4.161351e-11, 
    4.149003e-11, 4.160284e-11, 4.172148e-11, 4.205938e-11, 4.236508e-11, 
    4.269969e-11, 4.278177e-11, 4.317487e-11, 4.285474e-11, 4.338369e-11, 
    4.293379e-11, 4.37141e-11, 4.23173e-11, 4.292066e-11, 4.183076e-11, 
    4.194747e-11, 4.215902e-11, 4.264626e-11, 4.238284e-11, 4.269099e-11, 
    4.201197e-11, 4.166191e-11, 4.157156e-11, 4.140331e-11, 4.15754e-11, 
    4.156139e-11, 4.172639e-11, 4.167332e-11, 4.20706e-11, 4.185696e-11, 
    4.246534e-11, 4.26885e-11, 4.332194e-11, 4.371265e-11, 4.411221e-11, 
    4.428921e-11, 4.434316e-11, 4.436572e-11 ;

 F_NIT_vr =
  2.343415e-10, 2.353797e-10, 2.351772e-10, 2.360152e-10, 2.3555e-10, 
    2.360984e-10, 2.345507e-10, 2.354192e-10, 2.348644e-10, 2.344329e-10, 
    2.376411e-10, 2.360507e-10, 2.392953e-10, 2.382788e-10, 2.408325e-10, 
    2.391364e-10, 2.411746e-10, 2.407829e-10, 2.419608e-10, 2.416229e-10, 
    2.431305e-10, 2.42116e-10, 2.439125e-10, 2.428878e-10, 2.430477e-10, 
    2.420814e-10, 2.363722e-10, 2.374447e-10, 2.363083e-10, 2.364612e-10, 
    2.363923e-10, 2.355586e-10, 2.351388e-10, 2.3426e-10, 2.344191e-10, 
    2.350644e-10, 2.365282e-10, 2.360306e-10, 2.372838e-10, 2.372556e-10, 
    2.386522e-10, 2.380221e-10, 2.403726e-10, 2.397037e-10, 2.416367e-10, 
    2.411498e-10, 2.416133e-10, 2.414724e-10, 2.416145e-10, 2.409011e-10, 
    2.412062e-10, 2.405787e-10, 2.381429e-10, 2.388595e-10, 2.367226e-10, 
    2.354393e-10, 2.345877e-10, 2.339842e-10, 2.34069e-10, 2.342317e-10, 
    2.350676e-10, 2.358542e-10, 2.364541e-10, 2.368553e-10, 2.372508e-10, 
    2.384498e-10, 2.390845e-10, 2.405073e-10, 2.402502e-10, 2.406852e-10, 
    2.411012e-10, 2.417997e-10, 2.416845e-10, 2.419921e-10, 2.406724e-10, 
    2.415492e-10, 2.401019e-10, 2.404973e-10, 2.373608e-10, 2.361658e-10, 
    2.356582e-10, 2.35214e-10, 2.341344e-10, 2.348796e-10, 2.345855e-10, 
    2.352843e-10, 2.357287e-10, 2.355085e-10, 2.36866e-10, 2.363376e-10, 
    2.391218e-10, 2.379217e-10, 2.410529e-10, 2.403024e-10, 2.412321e-10, 
    2.407575e-10, 2.415704e-10, 2.408383e-10, 2.421063e-10, 2.423827e-10, 
    2.421933e-10, 2.429191e-10, 2.407963e-10, 2.416109e-10, 2.355037e-10, 
    2.355396e-10, 2.357064e-10, 2.349718e-10, 2.349269e-10, 2.342542e-10, 
    2.348521e-10, 2.351069e-10, 2.357538e-10, 2.361365e-10, 2.365003e-10, 
    2.373016e-10, 2.381967e-10, 2.394497e-10, 2.403507e-10, 2.409549e-10, 
    2.405841e-10, 2.40911e-10, 2.40545e-10, 2.403732e-10, 2.422784e-10, 
    2.412081e-10, 2.42814e-10, 2.427251e-10, 2.419976e-10, 2.427344e-10, 
    2.355643e-10, 2.353576e-10, 2.346415e-10, 2.352014e-10, 2.341805e-10, 
    2.347517e-10, 2.3508e-10, 2.363483e-10, 2.366269e-10, 2.368857e-10, 
    2.373966e-10, 2.380525e-10, 2.392047e-10, 2.402077e-10, 2.411244e-10, 
    2.410568e-10, 2.410804e-10, 2.412849e-10, 2.407773e-10, 2.413678e-10, 
    2.414666e-10, 2.412074e-10, 2.427125e-10, 2.422822e-10, 2.427222e-10, 
    2.424416e-10, 2.354244e-10, 2.357713e-10, 2.355833e-10, 2.359362e-10, 
    2.356871e-10, 2.36793e-10, 2.371244e-10, 2.386778e-10, 2.380396e-10, 
    2.39055e-10, 2.381422e-10, 2.383039e-10, 2.390874e-10, 2.381909e-10, 
    2.401517e-10, 2.388215e-10, 2.412926e-10, 2.39963e-10, 2.413754e-10, 
    2.411184e-10, 2.415431e-10, 2.419238e-10, 2.424024e-10, 2.43287e-10, 
    2.430816e-10, 2.438217e-10, 2.362888e-10, 2.367392e-10, 2.366994e-10, 
    2.371709e-10, 2.375196e-10, 2.382767e-10, 2.394916e-10, 2.390341e-10, 
    2.398731e-10, 2.400417e-10, 2.387661e-10, 2.395489e-10, 2.370384e-10, 
    2.374432e-10, 2.372019e-10, 2.363207e-10, 2.391374e-10, 2.376905e-10, 
    2.403627e-10, 2.395779e-10, 2.418688e-10, 2.407287e-10, 2.429686e-10, 
    2.439276e-10, 2.448305e-10, 2.458864e-10, 2.36985e-10, 2.366782e-10, 
    2.372265e-10, 2.37986e-10, 2.386905e-10, 2.396286e-10, 2.397243e-10, 
    2.398997e-10, 2.403549e-10, 2.407381e-10, 2.399548e-10, 2.408335e-10, 
    2.375369e-10, 2.39263e-10, 2.365593e-10, 2.373727e-10, 2.379378e-10, 
    2.376897e-10, 2.389787e-10, 2.392825e-10, 2.405185e-10, 2.398793e-10, 
    2.436902e-10, 2.420024e-10, 2.466908e-10, 2.453788e-10, 2.36571e-10, 
    2.369829e-10, 2.384187e-10, 2.377352e-10, 2.396905e-10, 2.401725e-10, 
    2.405638e-10, 2.41065e-10, 2.411186e-10, 2.414157e-10, 2.409285e-10, 
    2.41396e-10, 2.39628e-10, 2.404175e-10, 2.382518e-10, 2.387781e-10, 
    2.385357e-10, 2.382696e-10, 2.390897e-10, 2.399644e-10, 2.399828e-10, 
    2.402629e-10, 2.410538e-10, 2.39694e-10, 2.439072e-10, 2.41303e-10, 
    2.374324e-10, 2.382269e-10, 2.383402e-10, 2.380322e-10, 2.401235e-10, 
    2.393652e-10, 2.414085e-10, 2.408554e-10, 2.417608e-10, 2.413107e-10, 
    2.41244e-10, 2.406662e-10, 2.40306e-10, 2.39398e-10, 2.386591e-10, 
    2.38074e-10, 2.382095e-10, 2.388525e-10, 2.400172e-10, 2.411205e-10, 
    2.408784e-10, 2.416889e-10, 2.395437e-10, 2.404426e-10, 2.400946e-10, 
    2.41001e-10, 2.390209e-10, 2.407111e-10, 2.38589e-10, 2.387746e-10, 
    2.393494e-10, 2.405073e-10, 2.40763e-10, 2.410369e-10, 2.408674e-10, 
    2.400486e-10, 2.399141e-10, 2.393339e-10, 2.391735e-10, 2.387319e-10, 
    2.383659e-10, 2.386999e-10, 2.390501e-10, 2.40047e-10, 2.409457e-10, 
    2.419263e-10, 2.421663e-10, 2.433133e-10, 2.423791e-10, 2.439205e-10, 
    2.426094e-10, 2.448793e-10, 2.408085e-10, 2.425759e-10, 2.393757e-10, 
    2.397196e-10, 2.403424e-10, 2.417724e-10, 2.409997e-10, 2.419031e-10, 
    2.399087e-10, 2.388751e-10, 2.386076e-10, 2.381093e-10, 2.386185e-10, 
    2.385771e-10, 2.390647e-10, 2.389075e-10, 2.400794e-10, 2.394497e-10, 
    2.412391e-10, 2.418931e-10, 2.437413e-10, 2.448755e-10, 2.460313e-10, 
    2.465415e-10, 2.466969e-10, 2.467616e-10,
  1.334684e-10, 1.344761e-10, 1.3428e-10, 1.350943e-10, 1.346424e-10, 
    1.351759e-10, 1.336725e-10, 1.345161e-10, 1.339774e-10, 1.33559e-10, 
    1.366798e-10, 1.351307e-10, 1.382958e-10, 1.373029e-10, 1.398022e-10, 
    1.381411e-10, 1.40138e-10, 1.397542e-10, 1.409105e-10, 1.405789e-10, 
    1.420616e-10, 1.410637e-10, 1.428324e-10, 1.41823e-10, 1.419807e-10, 
    1.410308e-10, 1.35442e-10, 1.364866e-10, 1.353802e-10, 1.355289e-10, 
    1.354622e-10, 1.346517e-10, 1.342439e-10, 1.333915e-10, 1.335461e-10, 
    1.341723e-10, 1.355958e-10, 1.35112e-10, 1.363326e-10, 1.36305e-10, 
    1.376685e-10, 1.370531e-10, 1.393522e-10, 1.386974e-10, 1.405927e-10, 
    1.401152e-10, 1.405703e-10, 1.404322e-10, 1.405721e-10, 1.39872e-10, 
    1.401718e-10, 1.395563e-10, 1.371683e-10, 1.378686e-10, 1.357839e-10, 
    1.345359e-10, 1.337094e-10, 1.331241e-10, 1.332068e-10, 1.333645e-10, 
    1.341759e-10, 1.349406e-10, 1.355244e-10, 1.359154e-10, 1.363011e-10, 
    1.374708e-10, 1.380915e-10, 1.394848e-10, 1.39233e-10, 1.396596e-10, 
    1.400677e-10, 1.407538e-10, 1.406408e-10, 1.409434e-10, 1.396484e-10, 
    1.405085e-10, 1.390896e-10, 1.394772e-10, 1.364059e-10, 1.352425e-10, 
    1.34749e-10, 1.343177e-10, 1.332704e-10, 1.339933e-10, 1.337081e-10, 
    1.343869e-10, 1.348189e-10, 1.346052e-10, 1.359261e-10, 1.35412e-10, 
    1.381283e-10, 1.369559e-10, 1.400201e-10, 1.392846e-10, 1.401966e-10, 
    1.39731e-10, 1.405291e-10, 1.398107e-10, 1.41056e-10, 1.413277e-10, 
    1.41142e-10, 1.418558e-10, 1.397709e-10, 1.405703e-10, 1.345992e-10, 
    1.34634e-10, 1.347964e-10, 1.340831e-10, 1.340396e-10, 1.333873e-10, 
    1.339676e-10, 1.342151e-10, 1.348439e-10, 1.352164e-10, 1.355708e-10, 
    1.363513e-10, 1.372249e-10, 1.384498e-10, 1.393323e-10, 1.399249e-10, 
    1.395614e-10, 1.398823e-10, 1.395236e-10, 1.393556e-10, 1.412259e-10, 
    1.401746e-10, 1.41753e-10, 1.416655e-10, 1.409505e-10, 1.416754e-10, 
    1.346585e-10, 1.34458e-10, 1.337628e-10, 1.343068e-10, 1.333163e-10, 
    1.338704e-10, 1.341893e-10, 1.354227e-10, 1.356943e-10, 1.359462e-10, 
    1.364444e-10, 1.370846e-10, 1.382104e-10, 1.391926e-10, 1.400915e-10, 
    1.400256e-10, 1.400488e-10, 1.402498e-10, 1.39752e-10, 1.403316e-10, 
    1.40429e-10, 1.401745e-10, 1.416538e-10, 1.412306e-10, 1.416637e-10, 
    1.413881e-10, 1.345232e-10, 1.348606e-10, 1.346782e-10, 1.350213e-10, 
    1.347796e-10, 1.358556e-10, 1.361788e-10, 1.376949e-10, 1.37072e-10, 
    1.380639e-10, 1.371726e-10, 1.373304e-10, 1.380963e-10, 1.372208e-10, 
    1.391384e-10, 1.378372e-10, 1.402576e-10, 1.389545e-10, 1.403394e-10, 
    1.400876e-10, 1.405047e-10, 1.408786e-10, 1.413495e-10, 1.422198e-10, 
    1.420181e-10, 1.427471e-10, 1.353643e-10, 1.35803e-10, 1.357644e-10, 
    1.362241e-10, 1.365644e-10, 1.373031e-10, 1.384909e-10, 1.380438e-10, 
    1.38865e-10, 1.390301e-10, 1.377827e-10, 1.385481e-10, 1.36097e-10, 
    1.364919e-10, 1.362567e-10, 1.353989e-10, 1.381468e-10, 1.36734e-10, 
    1.393469e-10, 1.385785e-10, 1.408252e-10, 1.397062e-10, 1.419071e-10, 
    1.428517e-10, 1.437427e-10, 1.447864e-10, 1.360427e-10, 1.357444e-10, 
    1.362788e-10, 1.370195e-10, 1.37708e-10, 1.386253e-10, 1.387193e-10, 
    1.388915e-10, 1.393377e-10, 1.397133e-10, 1.389459e-10, 1.398075e-10, 
    1.365835e-10, 1.382697e-10, 1.356316e-10, 1.36424e-10, 1.369758e-10, 
    1.367337e-10, 1.379928e-10, 1.382901e-10, 1.395008e-10, 1.388745e-10, 
    1.426183e-10, 1.409576e-10, 1.455829e-10, 1.44285e-10, 1.356402e-10, 
    1.360417e-10, 1.374426e-10, 1.367754e-10, 1.386867e-10, 1.391586e-10, 
    1.395426e-10, 1.400341e-10, 1.400872e-10, 1.403787e-10, 1.399011e-10, 
    1.403598e-10, 1.386273e-10, 1.394006e-10, 1.372823e-10, 1.377968e-10, 
    1.3756e-10, 1.373004e-10, 1.381021e-10, 1.389579e-10, 1.389763e-10, 
    1.392511e-10, 1.400266e-10, 1.386944e-10, 1.428331e-10, 1.402719e-10, 
    1.364801e-10, 1.372556e-10, 1.373666e-10, 1.370659e-10, 1.391112e-10, 
    1.383689e-10, 1.403716e-10, 1.398293e-10, 1.407183e-10, 1.402763e-10, 
    1.402113e-10, 1.396444e-10, 1.39292e-10, 1.384029e-10, 1.376809e-10, 
    1.371095e-10, 1.372423e-10, 1.378703e-10, 1.390104e-10, 1.40092e-10, 
    1.398548e-10, 1.406506e-10, 1.385478e-10, 1.394281e-10, 1.390876e-10, 
    1.399761e-10, 1.380319e-10, 1.396868e-10, 1.376101e-10, 1.377917e-10, 
    1.383541e-10, 1.394879e-10, 1.397392e-10, 1.400077e-10, 1.39842e-10, 
    1.390393e-10, 1.38908e-10, 1.383405e-10, 1.381839e-10, 1.377522e-10, 
    1.373951e-10, 1.377213e-10, 1.380642e-10, 1.390397e-10, 1.399209e-10, 
    1.408839e-10, 1.411199e-10, 1.422487e-10, 1.413295e-10, 1.428474e-10, 
    1.415565e-10, 1.437938e-10, 1.397829e-10, 1.415187e-10, 1.383798e-10, 
    1.387167e-10, 1.393269e-10, 1.407301e-10, 1.399719e-10, 1.408587e-10, 
    1.389029e-10, 1.37892e-10, 1.376309e-10, 1.371442e-10, 1.37642e-10, 
    1.376015e-10, 1.380784e-10, 1.379251e-10, 1.390721e-10, 1.384556e-10, 
    1.402096e-10, 1.408517e-10, 1.426706e-10, 1.437897e-10, 1.449321e-10, 
    1.454374e-10, 1.455913e-10, 1.456556e-10,
  1.248466e-10, 1.259502e-10, 1.257353e-10, 1.266278e-10, 1.261324e-10, 
    1.267172e-10, 1.2507e-10, 1.25994e-10, 1.254038e-10, 1.249458e-10, 
    1.283672e-10, 1.266676e-10, 1.301429e-10, 1.290516e-10, 1.318004e-10, 
    1.299728e-10, 1.321703e-10, 1.317476e-10, 1.330215e-10, 1.32656e-10, 
    1.342909e-10, 1.331903e-10, 1.351417e-10, 1.340277e-10, 1.342017e-10, 
    1.331541e-10, 1.270089e-10, 1.281551e-10, 1.269412e-10, 1.271043e-10, 
    1.270311e-10, 1.261426e-10, 1.256958e-10, 1.247624e-10, 1.249317e-10, 
    1.256173e-10, 1.271777e-10, 1.266471e-10, 1.279861e-10, 1.279558e-10, 
    1.294533e-10, 1.287772e-10, 1.313051e-10, 1.305846e-10, 1.326713e-10, 
    1.321452e-10, 1.326465e-10, 1.324944e-10, 1.326485e-10, 1.318773e-10, 
    1.322075e-10, 1.315297e-10, 1.289037e-10, 1.296732e-10, 1.27384e-10, 
    1.260157e-10, 1.251105e-10, 1.244697e-10, 1.245602e-10, 1.247328e-10, 
    1.256214e-10, 1.264592e-10, 1.270993e-10, 1.275283e-10, 1.279515e-10, 
    1.292361e-10, 1.299182e-10, 1.31451e-10, 1.311738e-10, 1.316435e-10, 
    1.320929e-10, 1.328488e-10, 1.327242e-10, 1.330577e-10, 1.316311e-10, 
    1.325785e-10, 1.310161e-10, 1.314426e-10, 1.280665e-10, 1.267902e-10, 
    1.262492e-10, 1.257766e-10, 1.246298e-10, 1.254213e-10, 1.25109e-10, 
    1.258525e-10, 1.263258e-10, 1.260916e-10, 1.2754e-10, 1.269761e-10, 
    1.299587e-10, 1.286704e-10, 1.320404e-10, 1.312307e-10, 1.322348e-10, 
    1.317221e-10, 1.326012e-10, 1.318099e-10, 1.331819e-10, 1.334814e-10, 
    1.332767e-10, 1.340638e-10, 1.317661e-10, 1.326465e-10, 1.26085e-10, 
    1.261232e-10, 1.263012e-10, 1.255197e-10, 1.25472e-10, 1.247578e-10, 
    1.253932e-10, 1.256642e-10, 1.263533e-10, 1.267616e-10, 1.271503e-10, 
    1.280066e-10, 1.289659e-10, 1.303122e-10, 1.312831e-10, 1.319356e-10, 
    1.315354e-10, 1.318887e-10, 1.314937e-10, 1.313088e-10, 1.333691e-10, 
    1.322106e-10, 1.339505e-10, 1.33854e-10, 1.330656e-10, 1.338649e-10, 
    1.2615e-10, 1.259304e-10, 1.251689e-10, 1.257646e-10, 1.246801e-10, 
    1.252867e-10, 1.25636e-10, 1.269878e-10, 1.272857e-10, 1.275621e-10, 
    1.281088e-10, 1.288118e-10, 1.30049e-10, 1.311294e-10, 1.321191e-10, 
    1.320465e-10, 1.32072e-10, 1.322935e-10, 1.317452e-10, 1.323836e-10, 
    1.324908e-10, 1.322105e-10, 1.338411e-10, 1.333744e-10, 1.338519e-10, 
    1.33548e-10, 1.260018e-10, 1.263716e-10, 1.261717e-10, 1.265477e-10, 
    1.262827e-10, 1.274626e-10, 1.278173e-10, 1.294824e-10, 1.287979e-10, 
    1.298879e-10, 1.289085e-10, 1.290818e-10, 1.299235e-10, 1.289614e-10, 
    1.310698e-10, 1.296387e-10, 1.323021e-10, 1.308674e-10, 1.323922e-10, 
    1.321148e-10, 1.325742e-10, 1.329863e-10, 1.335055e-10, 1.344655e-10, 
    1.34243e-10, 1.350475e-10, 1.269238e-10, 1.27405e-10, 1.273626e-10, 
    1.27867e-10, 1.282406e-10, 1.290518e-10, 1.303574e-10, 1.298658e-10, 
    1.30769e-10, 1.309506e-10, 1.295788e-10, 1.304203e-10, 1.277275e-10, 
    1.28161e-10, 1.279029e-10, 1.269617e-10, 1.29979e-10, 1.284268e-10, 
    1.312992e-10, 1.304538e-10, 1.329275e-10, 1.316948e-10, 1.341205e-10, 
    1.35163e-10, 1.361473e-10, 1.373011e-10, 1.27668e-10, 1.273407e-10, 
    1.279271e-10, 1.287402e-10, 1.294967e-10, 1.305053e-10, 1.306087e-10, 
    1.30798e-10, 1.312891e-10, 1.317025e-10, 1.308579e-10, 1.318063e-10, 
    1.282615e-10, 1.301141e-10, 1.27217e-10, 1.280864e-10, 1.286923e-10, 
    1.284264e-10, 1.298097e-10, 1.301367e-10, 1.314687e-10, 1.307794e-10, 
    1.349054e-10, 1.330734e-10, 1.381825e-10, 1.367467e-10, 1.272264e-10, 
    1.276669e-10, 1.292051e-10, 1.284723e-10, 1.305727e-10, 1.310919e-10, 
    1.315147e-10, 1.320558e-10, 1.321143e-10, 1.324355e-10, 1.319094e-10, 
    1.324147e-10, 1.305074e-10, 1.313583e-10, 1.290289e-10, 1.295943e-10, 
    1.293341e-10, 1.290489e-10, 1.299299e-10, 1.308712e-10, 1.308914e-10, 
    1.311938e-10, 1.320476e-10, 1.305813e-10, 1.351425e-10, 1.323178e-10, 
    1.28148e-10, 1.289997e-10, 1.291215e-10, 1.287912e-10, 1.310398e-10, 
    1.302232e-10, 1.324276e-10, 1.318303e-10, 1.328096e-10, 1.323226e-10, 
    1.32251e-10, 1.316268e-10, 1.312388e-10, 1.302606e-10, 1.29467e-10, 
    1.288391e-10, 1.28985e-10, 1.296751e-10, 1.309289e-10, 1.321196e-10, 
    1.318584e-10, 1.327351e-10, 1.3042e-10, 1.313886e-10, 1.310139e-10, 
    1.31992e-10, 1.298528e-10, 1.316734e-10, 1.293891e-10, 1.295887e-10, 
    1.30207e-10, 1.314544e-10, 1.317311e-10, 1.320268e-10, 1.318443e-10, 
    1.309608e-10, 1.308163e-10, 1.30192e-10, 1.300198e-10, 1.295452e-10, 
    1.291529e-10, 1.295113e-10, 1.298882e-10, 1.309611e-10, 1.319312e-10, 
    1.329922e-10, 1.332524e-10, 1.344974e-10, 1.334835e-10, 1.351583e-10, 
    1.337337e-10, 1.362037e-10, 1.317793e-10, 1.33692e-10, 1.302352e-10, 
    1.306058e-10, 1.312772e-10, 1.328226e-10, 1.319874e-10, 1.329644e-10, 
    1.308106e-10, 1.296989e-10, 1.29412e-10, 1.288772e-10, 1.294242e-10, 
    1.293797e-10, 1.299039e-10, 1.297353e-10, 1.309968e-10, 1.303186e-10, 
    1.322492e-10, 1.329567e-10, 1.349631e-10, 1.361992e-10, 1.374623e-10, 
    1.380214e-10, 1.381918e-10, 1.38263e-10,
  1.280646e-10, 1.2928e-10, 1.290433e-10, 1.300267e-10, 1.294807e-10, 
    1.301253e-10, 1.283106e-10, 1.293284e-10, 1.286782e-10, 1.281738e-10, 
    1.319455e-10, 1.300707e-10, 1.339064e-10, 1.327008e-10, 1.357393e-10, 
    1.337184e-10, 1.361485e-10, 1.356807e-10, 1.370908e-10, 1.366861e-10, 
    1.384973e-10, 1.372778e-10, 1.394407e-10, 1.382056e-10, 1.383985e-10, 
    1.372376e-10, 1.304469e-10, 1.317114e-10, 1.303722e-10, 1.305521e-10, 
    1.304713e-10, 1.29492e-10, 1.289998e-10, 1.279719e-10, 1.281583e-10, 
    1.289134e-10, 1.30633e-10, 1.30048e-10, 1.315247e-10, 1.314913e-10, 
    1.331445e-10, 1.323979e-10, 1.351912e-10, 1.343945e-10, 1.36703e-10, 
    1.361207e-10, 1.366756e-10, 1.365072e-10, 1.366778e-10, 1.358243e-10, 
    1.361897e-10, 1.354397e-10, 1.325375e-10, 1.333873e-10, 1.308605e-10, 
    1.293523e-10, 1.283551e-10, 1.276498e-10, 1.277494e-10, 1.279394e-10, 
    1.289178e-10, 1.298409e-10, 1.305466e-10, 1.310196e-10, 1.314865e-10, 
    1.329046e-10, 1.336581e-10, 1.353526e-10, 1.35046e-10, 1.355656e-10, 
    1.360628e-10, 1.368996e-10, 1.367617e-10, 1.371309e-10, 1.355519e-10, 
    1.366003e-10, 1.348716e-10, 1.353434e-10, 1.316136e-10, 1.302057e-10, 
    1.296096e-10, 1.290888e-10, 1.27826e-10, 1.286974e-10, 1.283536e-10, 
    1.291723e-10, 1.296939e-10, 1.294358e-10, 1.310325e-10, 1.304107e-10, 
    1.337028e-10, 1.3228e-10, 1.360048e-10, 1.351089e-10, 1.362199e-10, 
    1.356525e-10, 1.366254e-10, 1.357496e-10, 1.372685e-10, 1.376003e-10, 
    1.373735e-10, 1.382456e-10, 1.357011e-10, 1.366756e-10, 1.294286e-10, 
    1.294706e-10, 1.296667e-10, 1.288058e-10, 1.287532e-10, 1.279668e-10, 
    1.286665e-10, 1.289649e-10, 1.297241e-10, 1.301742e-10, 1.306028e-10, 
    1.315474e-10, 1.326061e-10, 1.340935e-10, 1.351669e-10, 1.358888e-10, 
    1.354459e-10, 1.358369e-10, 1.353999e-10, 1.351953e-10, 1.374759e-10, 
    1.361931e-10, 1.3812e-10, 1.38013e-10, 1.371397e-10, 1.380251e-10, 
    1.295002e-10, 1.292581e-10, 1.284194e-10, 1.290756e-10, 1.278813e-10, 
    1.285492e-10, 1.289339e-10, 1.304237e-10, 1.30752e-10, 1.310569e-10, 
    1.3166e-10, 1.32436e-10, 1.338025e-10, 1.34997e-10, 1.360918e-10, 
    1.360114e-10, 1.360397e-10, 1.362848e-10, 1.356781e-10, 1.363845e-10, 
    1.365033e-10, 1.361929e-10, 1.379987e-10, 1.374817e-10, 1.380108e-10, 
    1.37674e-10, 1.293368e-10, 1.297443e-10, 1.29524e-10, 1.299384e-10, 
    1.296464e-10, 1.309473e-10, 1.313385e-10, 1.331766e-10, 1.324207e-10, 
    1.336246e-10, 1.325428e-10, 1.327342e-10, 1.33664e-10, 1.326011e-10, 
    1.34931e-10, 1.333493e-10, 1.362943e-10, 1.347073e-10, 1.363941e-10, 
    1.36087e-10, 1.365956e-10, 1.370518e-10, 1.376269e-10, 1.386909e-10, 
    1.384442e-10, 1.393362e-10, 1.30353e-10, 1.308837e-10, 1.308369e-10, 
    1.313933e-10, 1.318055e-10, 1.32701e-10, 1.341434e-10, 1.336002e-10, 
    1.345983e-10, 1.347991e-10, 1.33283e-10, 1.342129e-10, 1.312394e-10, 
    1.317177e-10, 1.314328e-10, 1.303948e-10, 1.337253e-10, 1.320111e-10, 
    1.351847e-10, 1.342499e-10, 1.369868e-10, 1.356224e-10, 1.383084e-10, 
    1.394644e-10, 1.405564e-10, 1.418378e-10, 1.311738e-10, 1.308127e-10, 
    1.314595e-10, 1.323571e-10, 1.331924e-10, 1.343068e-10, 1.344211e-10, 
    1.346305e-10, 1.351735e-10, 1.356309e-10, 1.346967e-10, 1.357456e-10, 
    1.318288e-10, 1.338746e-10, 1.306763e-10, 1.316355e-10, 1.323041e-10, 
    1.320106e-10, 1.335381e-10, 1.338994e-10, 1.353722e-10, 1.346099e-10, 
    1.391787e-10, 1.371483e-10, 1.428172e-10, 1.41222e-10, 1.306866e-10, 
    1.311725e-10, 1.328703e-10, 1.320612e-10, 1.343814e-10, 1.349555e-10, 
    1.35423e-10, 1.360218e-10, 1.360865e-10, 1.36442e-10, 1.358597e-10, 
    1.364189e-10, 1.343092e-10, 1.352501e-10, 1.326757e-10, 1.333001e-10, 
    1.330127e-10, 1.326978e-10, 1.336709e-10, 1.347114e-10, 1.347337e-10, 
    1.350681e-10, 1.360129e-10, 1.343908e-10, 1.394418e-10, 1.36312e-10, 
    1.317033e-10, 1.326435e-10, 1.32778e-10, 1.324133e-10, 1.348979e-10, 
    1.339951e-10, 1.364333e-10, 1.357723e-10, 1.368562e-10, 1.36317e-10, 
    1.362378e-10, 1.355471e-10, 1.351178e-10, 1.340364e-10, 1.331595e-10, 
    1.324661e-10, 1.326272e-10, 1.333894e-10, 1.347752e-10, 1.360924e-10, 
    1.358033e-10, 1.367736e-10, 1.342125e-10, 1.352836e-10, 1.348692e-10, 
    1.359512e-10, 1.335857e-10, 1.355988e-10, 1.330735e-10, 1.33294e-10, 
    1.339772e-10, 1.353564e-10, 1.356625e-10, 1.359897e-10, 1.357877e-10, 
    1.348104e-10, 1.346506e-10, 1.339605e-10, 1.337703e-10, 1.33246e-10, 
    1.328126e-10, 1.332085e-10, 1.336249e-10, 1.348108e-10, 1.358838e-10, 
    1.370584e-10, 1.373465e-10, 1.387263e-10, 1.376026e-10, 1.394593e-10, 
    1.378801e-10, 1.406192e-10, 1.357159e-10, 1.378337e-10, 1.340083e-10, 
    1.344179e-10, 1.351604e-10, 1.368707e-10, 1.35946e-10, 1.370277e-10, 
    1.346444e-10, 1.334158e-10, 1.330987e-10, 1.325083e-10, 1.331123e-10, 
    1.330631e-10, 1.336422e-10, 1.334559e-10, 1.348503e-10, 1.341005e-10, 
    1.362358e-10, 1.370191e-10, 1.392426e-10, 1.406141e-10, 1.420168e-10, 
    1.426382e-10, 1.428275e-10, 1.429068e-10,
  1.381447e-10, 1.394323e-10, 1.391814e-10, 1.402239e-10, 1.39645e-10, 
    1.403284e-10, 1.384051e-10, 1.394835e-10, 1.387945e-10, 1.382603e-10, 
    1.422598e-10, 1.402705e-10, 1.443428e-10, 1.430616e-10, 1.462923e-10, 
    1.44143e-10, 1.467279e-10, 1.462299e-10, 1.477313e-10, 1.473003e-10, 
    1.492306e-10, 1.479305e-10, 1.502368e-10, 1.489194e-10, 1.491251e-10, 
    1.478878e-10, 1.406694e-10, 1.420112e-10, 1.405902e-10, 1.40781e-10, 
    1.406953e-10, 1.39657e-10, 1.391354e-10, 1.380465e-10, 1.382438e-10, 
    1.390437e-10, 1.408669e-10, 1.402464e-10, 1.418129e-10, 1.417774e-10, 
    1.43533e-10, 1.427399e-10, 1.457091e-10, 1.448616e-10, 1.473183e-10, 
    1.466982e-10, 1.472891e-10, 1.471098e-10, 1.472915e-10, 1.463827e-10, 
    1.467717e-10, 1.459734e-10, 1.428883e-10, 1.43791e-10, 1.411081e-10, 
    1.39509e-10, 1.384523e-10, 1.377054e-10, 1.378108e-10, 1.38012e-10, 
    1.390484e-10, 1.400268e-10, 1.407751e-10, 1.412769e-10, 1.417723e-10, 
    1.432783e-10, 1.440788e-10, 1.458808e-10, 1.455546e-10, 1.461074e-10, 
    1.466366e-10, 1.475276e-10, 1.473807e-10, 1.477741e-10, 1.460928e-10, 
    1.47209e-10, 1.45369e-10, 1.458709e-10, 1.419075e-10, 1.404136e-10, 
    1.397817e-10, 1.392296e-10, 1.37892e-10, 1.388149e-10, 1.384507e-10, 
    1.393181e-10, 1.398709e-10, 1.395973e-10, 1.412906e-10, 1.40631e-10, 
    1.441264e-10, 1.426147e-10, 1.465748e-10, 1.456215e-10, 1.468038e-10, 
    1.461998e-10, 1.472357e-10, 1.463032e-10, 1.479206e-10, 1.482742e-10, 
    1.480325e-10, 1.48962e-10, 1.462516e-10, 1.472892e-10, 1.395897e-10, 
    1.396343e-10, 1.398422e-10, 1.389298e-10, 1.388741e-10, 1.380411e-10, 
    1.387821e-10, 1.390984e-10, 1.39903e-10, 1.403802e-10, 1.408347e-10, 
    1.41837e-10, 1.429612e-10, 1.445416e-10, 1.456832e-10, 1.464513e-10, 
    1.4598e-10, 1.463961e-10, 1.45931e-10, 1.457133e-10, 1.481417e-10, 
    1.467753e-10, 1.488281e-10, 1.487141e-10, 1.477835e-10, 1.487269e-10, 
    1.396656e-10, 1.394091e-10, 1.385205e-10, 1.392156e-10, 1.379505e-10, 
    1.386579e-10, 1.390656e-10, 1.406448e-10, 1.409931e-10, 1.413165e-10, 
    1.419566e-10, 1.427804e-10, 1.442323e-10, 1.455024e-10, 1.466674e-10, 
    1.465819e-10, 1.46612e-10, 1.468729e-10, 1.462271e-10, 1.469791e-10, 
    1.471056e-10, 1.467751e-10, 1.486988e-10, 1.481478e-10, 1.487117e-10, 
    1.483527e-10, 1.394924e-10, 1.399244e-10, 1.396909e-10, 1.401302e-10, 
    1.398206e-10, 1.412002e-10, 1.416154e-10, 1.435671e-10, 1.427642e-10, 
    1.440432e-10, 1.428938e-10, 1.430971e-10, 1.440852e-10, 1.429558e-10, 
    1.454323e-10, 1.437507e-10, 1.468831e-10, 1.451944e-10, 1.469893e-10, 
    1.466624e-10, 1.472039e-10, 1.476899e-10, 1.483025e-10, 1.494369e-10, 
    1.491738e-10, 1.501253e-10, 1.405698e-10, 1.411328e-10, 1.410831e-10, 
    1.416735e-10, 1.42111e-10, 1.430619e-10, 1.445947e-10, 1.440172e-10, 
    1.450784e-10, 1.452919e-10, 1.436801e-10, 1.446686e-10, 1.415102e-10, 
    1.420178e-10, 1.417154e-10, 1.406142e-10, 1.441502e-10, 1.423293e-10, 
    1.457021e-10, 1.447079e-10, 1.476205e-10, 1.461679e-10, 1.49029e-10, 
    1.502621e-10, 1.514278e-10, 1.52797e-10, 1.414405e-10, 1.410574e-10, 
    1.417437e-10, 1.426966e-10, 1.435839e-10, 1.447684e-10, 1.448899e-10, 
    1.451126e-10, 1.456902e-10, 1.461768e-10, 1.451831e-10, 1.46299e-10, 
    1.421358e-10, 1.443089e-10, 1.409127e-10, 1.419306e-10, 1.426403e-10, 
    1.423287e-10, 1.439512e-10, 1.443352e-10, 1.459016e-10, 1.450906e-10, 
    1.499573e-10, 1.477927e-10, 1.538441e-10, 1.521388e-10, 1.409236e-10, 
    1.414391e-10, 1.432417e-10, 1.423824e-10, 1.448477e-10, 1.454582e-10, 
    1.459556e-10, 1.46593e-10, 1.466618e-10, 1.470403e-10, 1.464204e-10, 
    1.470158e-10, 1.447709e-10, 1.457716e-10, 1.43035e-10, 1.436983e-10, 
    1.433929e-10, 1.430584e-10, 1.440923e-10, 1.451987e-10, 1.452223e-10, 
    1.455781e-10, 1.465837e-10, 1.448577e-10, 1.502382e-10, 1.469021e-10, 
    1.420025e-10, 1.430009e-10, 1.431437e-10, 1.427563e-10, 1.45397e-10, 
    1.444369e-10, 1.470311e-10, 1.463273e-10, 1.474814e-10, 1.469073e-10, 
    1.468229e-10, 1.460876e-10, 1.45631e-10, 1.444809e-10, 1.43549e-10, 
    1.428124e-10, 1.429835e-10, 1.437933e-10, 1.452665e-10, 1.466681e-10, 
    1.463604e-10, 1.473935e-10, 1.446681e-10, 1.458074e-10, 1.453665e-10, 
    1.465177e-10, 1.440019e-10, 1.46143e-10, 1.434575e-10, 1.436918e-10, 
    1.444179e-10, 1.458849e-10, 1.462105e-10, 1.465588e-10, 1.463438e-10, 
    1.45304e-10, 1.45134e-10, 1.444002e-10, 1.44198e-10, 1.436408e-10, 
    1.431804e-10, 1.43601e-10, 1.440435e-10, 1.453044e-10, 1.464461e-10, 
    1.476968e-10, 1.480037e-10, 1.494748e-10, 1.482768e-10, 1.502569e-10, 
    1.485727e-10, 1.514951e-10, 1.462675e-10, 1.485231e-10, 1.44451e-10, 
    1.448865e-10, 1.456763e-10, 1.474969e-10, 1.465123e-10, 1.476641e-10, 
    1.451273e-10, 1.438213e-10, 1.434843e-10, 1.428571e-10, 1.434987e-10, 
    1.434465e-10, 1.440618e-10, 1.438639e-10, 1.453464e-10, 1.44549e-10, 
    1.468208e-10, 1.47655e-10, 1.500254e-10, 1.514895e-10, 1.529881e-10, 
    1.536525e-10, 1.538551e-10, 1.539398e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24531.77, 24551.66, 24547.76, 24564.04, 24554.97, 24565.69, 24535.77, 
    24552.46, 24541.77, 24533.54, 24596.37, 24564.77, 24630.23, 24609.29, 
    24662.33, 24626.94, 24669.6, 24661.29, 24686.51, 24679.21, 24712.26, 
    24689.9, 24729.86, 24706.87, 24710.43, 24689.17, 24571.06, 24592.39, 
    24569.81, 24572.83, 24571.47, 24555.16, 24547.05, 24530.27, 24533.29, 
    24545.63, 24574.19, 24564.4, 24589.23, 24588.66, 24616.95, 24604.09, 
    24652.66, 24638.75, 24679.52, 24669.1, 24679.03, 24676.01, 24679.07, 
    24663.83, 24670.33, 24657.03, 24606.49, 24621.17, 24578.02, 24552.86, 
    24536.5, 24525.05, 24526.66, 24529.74, 24545.7, 24560.95, 24572.73, 
    24580.7, 24588.58, 24612.81, 24625.88, 24655.5, 24650.11, 24659.25, 
    24668.07, 24683.06, 24680.57, 24687.24, 24659.01, 24677.68, 24647.06, 
    24655.33, 24590.74, 24567.03, 24557.11, 24548.51, 24527.9, 24542.09, 
    24536.47, 24549.88, 24558.51, 24554.23, 24580.92, 24570.46, 24626.66, 
    24602.07, 24667.04, 24651.21, 24670.87, 24660.79, 24678.13, 24662.51, 
    24689.73, 24695.77, 24691.64, 24707.61, 24661.65, 24679.03, 24554.11, 
    24554.81, 24558.06, 24543.86, 24543, 24530.19, 24541.58, 24546.47, 
    24559.01, 24566.5, 24573.68, 24589.61, 24607.66, 24633.51, 24652.23, 
    24664.98, 24657.14, 24664.06, 24656.33, 24652.73, 24693.5, 24670.39, 
    24705.29, 24703.33, 24687.4, 24703.55, 24555.3, 24551.3, 24537.54, 
    24548.29, 24528.8, 24539.66, 24545.96, 24570.68, 24576.19, 24581.33, 
    24591.52, 24604.74, 24628.41, 24649.25, 24668.59, 24667.16, 24667.66, 
    24672.03, 24661.24, 24673.81, 24675.94, 24670.39, 24703.06, 24693.61, 
    24703.29, 24697.12, 24552.6, 24559.34, 24555.69, 24562.57, 24557.72, 
    24579.48, 24586.09, 24617.51, 24604.48, 24625.3, 24606.58, 24609.87, 
    24625.99, 24607.58, 24648.1, 24620.51, 24672.2, 24644.19, 24673.98, 
    24668.5, 24677.59, 24685.81, 24696.25, 24715.85, 24711.28, 24727.89, 
    24569.49, 24578.41, 24577.62, 24587.01, 24593.99, 24609.29, 24634.38, 
    24624.87, 24642.29, 24645.79, 24619.35, 24635.6, 24584.41, 24592.5, 
    24587.68, 24570.19, 24627.06, 24597.48, 24652.54, 24636.24, 24684.63, 
    24660.26, 24708.77, 24730.31, 24751.01, 24775.66, 24583.31, 24577.21, 
    24588.13, 24603.39, 24617.78, 24637.23, 24639.21, 24642.85, 24652.35, 
    24660.41, 24644.01, 24662.44, 24594.39, 24629.67, 24574.92, 24591.11, 
    24602.49, 24597.47, 24623.79, 24630.1, 24655.84, 24642.49, 24724.94, 
    24687.56, 24794.64, 24763.83, 24575.09, 24583.29, 24612.21, 24598.34, 
    24638.52, 24648.52, 24656.74, 24667.34, 24668.49, 24674.84, 24664.46, 
    24674.42, 24637.27, 24653.69, 24608.86, 24619.65, 24614.67, 24609.24, 
    24626.1, 24644.26, 24644.65, 24650.5, 24667.19, 24638.68, 24729.88, 
    24672.52, 24592.25, 24608.31, 24610.62, 24604.35, 24647.52, 24631.78, 
    24674.68, 24662.91, 24682.28, 24672.6, 24671.19, 24658.93, 24651.37, 
    24632.5, 24617.21, 24605.26, 24608.03, 24621.2, 24645.37, 24668.6, 
    24663.46, 24680.79, 24635.6, 24654.28, 24647.02, 24666.09, 24624.62, 
    24659.85, 24615.72, 24619.54, 24631.46, 24655.57, 24660.97, 24666.77, 
    24663.19, 24645.99, 24643.2, 24631.17, 24627.84, 24618.71, 24611.22, 
    24618.06, 24625.3, 24646, 24664.89, 24685.93, 24691.15, 24716.51, 
    24695.81, 24730.22, 24700.89, 24752.22, 24661.92, 24700.04, 24632.01, 
    24639.15, 24652.12, 24682.54, 24666, 24685.37, 24643.09, 24621.66, 
    24616.16, 24605.98, 24616.39, 24615.54, 24625.6, 24622.36, 24646.69, 
    24633.63, 24671.15, 24685.22, 24726.14, 24752.12, 24779.11, 24791.15, 
    24794.84, 24796.39 ;

 GC_ICE1 =
  17605.52, 17637.29, 17631.06, 17657.06, 17642.58, 17659.69, 17611.9, 
    17638.56, 17621.49, 17608.35, 17708.67, 17658.23, 17762.69, 17729.29, 
    17813.81, 17757.45, 17825.38, 17812.16, 17852.29, 17840.68, 17893.26, 
    17857.68, 17921.25, 17884.69, 17890.35, 17856.52, 17668.28, 17702.33, 
    17666.28, 17671.1, 17668.93, 17642.88, 17629.92, 17603.12, 17607.95, 
    17627.65, 17673.27, 17657.63, 17697.28, 17696.38, 17741.51, 17720.99, 
    17798.42, 17776.27, 17841.16, 17824.59, 17840.38, 17835.57, 17840.44, 
    17816.21, 17826.54, 17805.38, 17724.81, 17748.23, 17679.38, 17639.19, 
    17613.06, 17594.79, 17597.36, 17602.27, 17627.76, 17652.12, 17670.95, 
    17683.67, 17696.24, 17734.9, 17755.76, 17802.94, 17794.36, 17808.92, 
    17822.95, 17846.79, 17842.84, 17853.45, 17808.53, 17838.23, 17789.5, 
    17802.67, 17699.69, 17661.83, 17645.99, 17632.25, 17599.34, 17621.99, 
    17613.02, 17634.45, 17648.22, 17641.39, 17684.02, 17667.3, 17757.01, 
    17717.77, 17821.3, 17796.12, 17827.4, 17811.36, 17838.95, 17814.1, 
    17857.41, 17867.02, 17860.45, 17885.86, 17812.73, 17840.38, 17641.2, 
    17642.31, 17647.5, 17624.83, 17623.45, 17602.98, 17621.18, 17629, 
    17649.02, 17660.99, 17672.45, 17697.89, 17726.7, 17767.93, 17797.74, 
    17818.03, 17805.55, 17816.56, 17804.26, 17798.53, 17863.41, 17826.64, 
    17882.18, 17879.04, 17853.7, 17879.4, 17643.09, 17636.71, 17614.74, 
    17631.9, 17600.77, 17618.12, 17628.19, 17667.65, 17676.46, 17684.68, 
    17700.93, 17722.04, 17759.79, 17792.99, 17823.77, 17821.49, 17822.29, 
    17829.24, 17812.08, 17832.08, 17835.46, 17826.63, 17878.63, 17863.58, 
    17878.98, 17869.16, 17638.78, 17649.56, 17643.72, 17654.71, 17646.96, 
    17681.72, 17692.26, 17742.4, 17721.62, 17754.83, 17724.96, 17730.21, 
    17755.93, 17726.55, 17791.16, 17747.18, 17829.51, 17784.94, 17832.35, 
    17823.63, 17838.09, 17851.17, 17867.79, 17898.96, 17891.69, 17918.12, 
    17665.76, 17680.01, 17678.74, 17693.73, 17704.87, 17729.29, 17769.33, 
    17754.15, 17781.91, 17787.48, 17745.34, 17771.27, 17689.6, 17702.5, 
    17694.8, 17666.88, 17757.63, 17710.45, 17798.23, 17772.29, 17849.3, 
    17810.51, 17887.7, 17921.96, 17954.88, 17994.03, 17687.83, 17678.09, 
    17695.52, 17719.88, 17742.84, 17773.86, 17777.01, 17782.8, 17797.92, 
    17810.75, 17784.64, 17813.98, 17705.51, 17761.8, 17674.43, 17700.27, 
    17718.43, 17710.44, 17752.42, 17762.49, 17803.48, 17782.23, 17913.43, 
    17853.95, 18024.12, 17975.26, 17674.7, 17687.79, 17733.95, 17711.81, 
    17775.91, 17791.84, 17804.91, 17821.79, 17823.62, 17833.71, 17817.21, 
    17833.06, 17773.92, 17800.06, 17728.6, 17745.82, 17737.87, 17729.21, 
    17756.12, 17785.05, 17785.67, 17794.98, 17821.54, 17776.17, 17921.29, 
    17830.02, 17702.1, 17727.72, 17731.41, 17721.41, 17790.23, 17765.17, 
    17833.47, 17814.74, 17845.55, 17830.16, 17827.91, 17808.39, 17796.37, 
    17766.33, 17741.93, 17722.86, 17727.27, 17748.29, 17786.82, 17823.79, 
    17815.62, 17843.19, 17771.26, 17801, 17789.43, 17819.79, 17753.74, 
    17809.86, 17739.55, 17745.65, 17764.67, 17803.04, 17811.64, 17820.88, 
    17815.17, 17787.8, 17783.36, 17764.2, 17758.89, 17744.32, 17732.36, 
    17743.28, 17754.84, 17787.81, 17817.89, 17851.36, 17859.67, 17900.01, 
    17867.09, 17921.82, 17875.17, 17956.8, 17813.15, 17873.82, 17765.54, 
    17776.92, 17797.56, 17845.97, 17819.64, 17850.48, 17783.19, 17749.03, 
    17740.25, 17724.01, 17740.62, 17739.26, 17755.31, 17750.14, 17788.91, 
    17768.12, 17827.85, 17850.23, 17915.33, 17956.64, 17999.5, 18018.58, 
    18024.43, 18026.89 ;

 GC_LIQ1 =
  5232.774, 5234.803, 5234.405, 5236.066, 5235.141, 5236.234, 5233.182, 
    5234.884, 5233.793, 5232.955, 5239.375, 5236.141, 5242.854, 5240.703, 
    5246.204, 5242.517, 5246.966, 5246.096, 5248.739, 5247.974, 5251.44, 
    5249.095, 5253.29, 5250.875, 5251.249, 5249.018, 5236.783, 5238.966, 
    5236.655, 5236.963, 5236.825, 5235.16, 5234.332, 5232.62, 5232.929, 
    5234.187, 5237.102, 5236.102, 5238.641, 5238.583, 5241.49, 5240.168, 
    5245.192, 5243.737, 5248.006, 5246.914, 5247.955, 5247.638, 5247.958, 
    5246.362, 5247.042, 5245.65, 5240.414, 5241.923, 5237.493, 5234.925, 
    5233.255, 5232.089, 5232.253, 5232.566, 5234.194, 5235.75, 5236.953, 
    5237.767, 5238.575, 5241.064, 5242.408, 5245.489, 5244.925, 5245.882, 
    5246.806, 5248.377, 5248.117, 5248.815, 5245.857, 5247.813, 5244.606, 
    5245.472, 5238.796, 5236.371, 5235.359, 5234.481, 5232.379, 5233.826, 
    5233.253, 5234.622, 5235.501, 5235.065, 5237.789, 5236.721, 5242.488, 
    5239.961, 5246.698, 5245.041, 5247.099, 5246.043, 5247.86, 5246.223, 
    5249.077, 5249.71, 5249.277, 5250.952, 5246.133, 5247.955, 5235.053, 
    5235.124, 5235.455, 5234.007, 5233.919, 5232.612, 5233.774, 5234.273, 
    5235.552, 5236.317, 5237.05, 5238.68, 5240.536, 5243.192, 5245.147, 
    5246.482, 5245.661, 5246.385, 5245.576, 5245.2, 5249.472, 5247.049, 
    5250.709, 5250.503, 5248.832, 5250.526, 5235.174, 5234.766, 5233.362, 
    5234.459, 5232.471, 5233.579, 5234.222, 5236.743, 5237.306, 5237.831, 
    5238.876, 5240.235, 5242.667, 5244.835, 5246.86, 5246.71, 5246.763, 
    5247.221, 5246.091, 5247.407, 5247.63, 5247.049, 5250.475, 5249.483, 
    5250.499, 5249.851, 5234.898, 5235.586, 5235.214, 5235.916, 5235.421, 
    5237.642, 5238.318, 5241.547, 5240.208, 5242.348, 5240.423, 5240.762, 
    5242.419, 5240.526, 5244.715, 5241.855, 5247.238, 5244.306, 5247.425, 
    5246.851, 5247.804, 5248.666, 5249.761, 5251.817, 5251.337, 5253.083, 
    5236.622, 5237.532, 5237.452, 5238.413, 5239.13, 5240.703, 5243.282, 
    5242.304, 5244.107, 5244.474, 5241.736, 5243.408, 5238.146, 5238.977, 
    5238.481, 5236.694, 5242.528, 5239.489, 5245.18, 5243.475, 5248.542, 
    5245.988, 5251.074, 5253.337, 5255.519, 5258.137, 5238.033, 5237.41, 
    5238.528, 5240.097, 5241.575, 5243.578, 5243.785, 5244.166, 5245.16, 
    5246.003, 5244.287, 5246.216, 5239.171, 5242.797, 5237.176, 5238.834, 
    5240.003, 5239.488, 5242.192, 5242.841, 5245.525, 5244.128, 5252.773, 
    5248.849, 5260.182, 5256.871, 5237.193, 5238.031, 5241.003, 5239.577, 
    5243.713, 5244.76, 5245.619, 5246.729, 5246.85, 5247.515, 5246.428, 
    5247.472, 5243.582, 5245.3, 5240.658, 5241.767, 5241.255, 5240.697, 
    5242.431, 5244.313, 5244.354, 5244.966, 5246.713, 5243.73, 5253.293, 
    5247.272, 5238.952, 5240.602, 5240.839, 5240.195, 5244.654, 5243.014, 
    5247.499, 5246.265, 5248.295, 5247.281, 5247.133, 5245.848, 5245.057, 
    5243.088, 5241.517, 5240.288, 5240.572, 5241.927, 5244.43, 5246.861, 
    5246.323, 5248.139, 5243.407, 5245.362, 5244.602, 5246.598, 5242.278, 
    5245.945, 5241.363, 5241.756, 5242.982, 5245.497, 5246.062, 5246.669, 
    5246.294, 5244.494, 5244.203, 5242.952, 5242.609, 5241.67, 5240.9, 
    5241.604, 5242.348, 5244.495, 5246.473, 5248.678, 5249.226, 5251.887, 
    5249.715, 5253.328, 5250.248, 5255.646, 5246.161, 5250.158, 5243.038, 
    5243.779, 5245.136, 5248.323, 5246.588, 5248.62, 5244.191, 5241.974, 
    5241.408, 5240.363, 5241.433, 5241.345, 5242.379, 5242.045, 5244.567, 
    5243.204, 5247.129, 5248.604, 5252.899, 5255.635, 5258.507, 5259.805, 
    5260.204, 5260.371 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.955614e-09, 8.994996e-09, 8.98734e-09, 9.019104e-09, 9.001483e-09, 
    9.022282e-09, 8.963598e-09, 8.996559e-09, 8.975517e-09, 8.959159e-09, 
    9.080747e-09, 9.02052e-09, 9.1433e-09, 9.104892e-09, 9.201374e-09, 
    9.137325e-09, 9.214289e-09, 9.199526e-09, 9.243957e-09, 9.231228e-09, 
    9.28806e-09, 9.249831e-09, 9.317519e-09, 9.27893e-09, 9.284967e-09, 
    9.248571e-09, 9.03264e-09, 9.073249e-09, 9.030234e-09, 9.036024e-09, 
    9.033426e-09, 9.001847e-09, 8.985934e-09, 8.952603e-09, 8.958654e-09, 
    8.983134e-09, 9.038629e-09, 9.01979e-09, 9.067265e-09, 9.066193e-09, 
    9.119047e-09, 9.095216e-09, 9.184049e-09, 9.158802e-09, 9.231759e-09, 
    9.213411e-09, 9.230898e-09, 9.225595e-09, 9.230966e-09, 9.204057e-09, 
    9.215587e-09, 9.191908e-09, 9.09968e-09, 9.126786e-09, 9.045943e-09, 
    8.997334e-09, 8.965044e-09, 8.942131e-09, 8.945371e-09, 8.951545e-09, 
    8.983277e-09, 9.013111e-09, 9.035847e-09, 9.051054e-09, 9.066039e-09, 
    9.111399e-09, 9.135404e-09, 9.189155e-09, 9.179454e-09, 9.195888e-09, 
    9.211586e-09, 9.237944e-09, 9.233605e-09, 9.245217e-09, 9.195453e-09, 
    9.228527e-09, 9.173928e-09, 9.188861e-09, 9.070117e-09, 9.024872e-09, 
    9.005644e-09, 8.988811e-09, 8.947861e-09, 8.976141e-09, 8.964992e-09, 
    8.991513e-09, 9.008366e-09, 9.000031e-09, 9.051471e-09, 9.031472e-09, 
    9.136826e-09, 9.091448e-09, 9.209755e-09, 9.181445e-09, 9.21654e-09, 
    9.198631e-09, 9.229317e-09, 9.201701e-09, 9.249539e-09, 9.259956e-09, 
    9.252838e-09, 9.280182e-09, 9.20017e-09, 9.230898e-09, 8.999797e-09, 
    9.001157e-09, 9.00749e-09, 8.979653e-09, 8.977949e-09, 8.952438e-09, 
    8.975138e-09, 8.984804e-09, 9.009343e-09, 9.023857e-09, 9.037655e-09, 
    9.067991e-09, 9.101871e-09, 9.149246e-09, 9.18328e-09, 9.206094e-09, 
    9.192104e-09, 9.204455e-09, 9.190648e-09, 9.184177e-09, 9.256053e-09, 
    9.215694e-09, 9.276248e-09, 9.272898e-09, 9.245494e-09, 9.273275e-09, 
    9.002111e-09, 8.994289e-09, 8.96713e-09, 8.988384e-09, 8.94966e-09, 
    8.971337e-09, 8.9838e-09, 9.031891e-09, 9.042456e-09, 9.052254e-09, 
    9.071603e-09, 9.096436e-09, 9.139998e-09, 9.1779e-09, 9.212499e-09, 
    9.209963e-09, 9.210856e-09, 9.218586e-09, 9.19944e-09, 9.221729e-09, 
    9.22547e-09, 9.215689e-09, 9.272449e-09, 9.256233e-09, 9.272827e-09, 
    9.262268e-09, 8.996832e-09, 9.009994e-09, 9.002881e-09, 9.016256e-09, 
    9.006834e-09, 9.048732e-09, 9.061294e-09, 9.120071e-09, 9.095948e-09, 
    9.134339e-09, 9.099847e-09, 9.105959e-09, 9.135593e-09, 9.10171e-09, 
    9.175811e-09, 9.125575e-09, 9.218886e-09, 9.168723e-09, 9.22203e-09, 
    9.212349e-09, 9.228377e-09, 9.242732e-09, 9.26079e-09, 9.294112e-09, 
    9.286396e-09, 9.314261e-09, 9.029616e-09, 9.046689e-09, 9.045185e-09, 
    9.063051e-09, 9.076264e-09, 9.104902e-09, 9.150832e-09, 9.13356e-09, 
    9.165268e-09, 9.171634e-09, 9.123461e-09, 9.153039e-09, 9.058114e-09, 
    9.073451e-09, 9.064319e-09, 9.030964e-09, 9.137541e-09, 9.082846e-09, 
    9.183842e-09, 9.154213e-09, 9.240686e-09, 9.197682e-09, 9.282148e-09, 
    9.318259e-09, 9.35224e-09, 9.391956e-09, 9.056006e-09, 9.044405e-09, 
    9.065175e-09, 9.093913e-09, 9.120575e-09, 9.156021e-09, 9.159647e-09, 
    9.166287e-09, 9.183487e-09, 9.197949e-09, 9.168388e-09, 9.201575e-09, 
    9.07701e-09, 9.142289e-09, 9.04002e-09, 9.070817e-09, 9.092219e-09, 
    9.08283e-09, 9.131586e-09, 9.143077e-09, 9.189773e-09, 9.165634e-09, 
    9.309347e-09, 9.245765e-09, 9.422193e-09, 9.37289e-09, 9.040352e-09, 
    9.055965e-09, 9.110305e-09, 9.08445e-09, 9.158387e-09, 9.176586e-09, 
    9.19138e-09, 9.210292e-09, 9.212334e-09, 9.223539e-09, 9.205177e-09, 
    9.222814e-09, 9.156096e-09, 9.185911e-09, 9.104093e-09, 9.124007e-09, 
    9.114845e-09, 9.104796e-09, 9.13581e-09, 9.168853e-09, 9.169558e-09, 
    9.180154e-09, 9.210012e-09, 9.158686e-09, 9.317556e-09, 9.219444e-09, 
    9.07299e-09, 9.103065e-09, 9.107358e-09, 9.095709e-09, 9.174761e-09, 
    9.146119e-09, 9.223266e-09, 9.202416e-09, 9.236578e-09, 9.219602e-09, 
    9.217104e-09, 9.195301e-09, 9.181726e-09, 9.147432e-09, 9.119527e-09, 
    9.097398e-09, 9.102544e-09, 9.126851e-09, 9.170875e-09, 9.212519e-09, 
    9.203397e-09, 9.233982e-09, 9.153026e-09, 9.186973e-09, 9.173853e-09, 
    9.208063e-09, 9.133101e-09, 9.196939e-09, 9.116784e-09, 9.123812e-09, 
    9.14555e-09, 9.189276e-09, 9.198948e-09, 9.209278e-09, 9.202903e-09, 
    9.171992e-09, 9.166927e-09, 9.145021e-09, 9.138973e-09, 9.122282e-09, 
    9.108462e-09, 9.121089e-09, 9.134348e-09, 9.172004e-09, 9.205939e-09, 
    9.242936e-09, 9.25199e-09, 9.295221e-09, 9.260031e-09, 9.318102e-09, 
    9.268733e-09, 9.354192e-09, 9.200637e-09, 9.267279e-09, 9.146539e-09, 
    9.159546e-09, 9.183074e-09, 9.237034e-09, 9.207902e-09, 9.241972e-09, 
    9.166729e-09, 9.127691e-09, 9.117589e-09, 9.098744e-09, 9.11802e-09, 
    9.116452e-09, 9.134897e-09, 9.12897e-09, 9.173254e-09, 9.149467e-09, 
    9.217042e-09, 9.241703e-09, 9.311342e-09, 9.354033e-09, 9.397487e-09, 
    9.416673e-09, 9.422512e-09, 9.424952e-09 ;

 H2OCAN =
  0.0599289, 0.05991397, 0.05991681, 0.05990487, 0.05991139, 0.05990365, 
    0.05992574, 0.05991349, 0.05992124, 0.05992737, 0.05988196, 0.05990431, 
    0.05985762, 0.05987198, 0.05983538, 0.05986004, 0.05983032, 0.05983579, 
    0.05981853, 0.05982347, 0.05980191, 0.05981624, 0.05979014, 0.05980518, 
    0.05980295, 0.05981677, 0.05989953, 0.05988485, 0.05990047, 0.05989837, 
    0.05989924, 0.05991136, 0.05991764, 0.05992983, 0.05992756, 0.0599185, 
    0.05989741, 0.05990439, 0.05988617, 0.05988657, 0.05986657, 0.05987556, 
    0.05984174, 0.05985131, 0.05982326, 0.0598304, 0.05982365, 0.05982566, 
    0.05982362, 0.05983406, 0.05982961, 0.05983868, 0.05987393, 0.05986371, 
    0.05989452, 0.0599135, 0.05992526, 0.0599338, 0.0599326, 0.05993036, 
    0.05991845, 0.05990693, 0.05989821, 0.05989241, 0.05988664, 0.05987005, 
    0.05986063, 0.05983995, 0.05984343, 0.05983732, 0.05983109, 0.05982095, 
    0.05982259, 0.05981817, 0.05983729, 0.0598247, 0.05984547, 0.05983984, 
    0.05988612, 0.05990246, 0.05991027, 0.0599163, 0.05993169, 0.05992113, 
    0.05992532, 0.05991511, 0.05990875, 0.05991185, 0.05989225, 0.05989993, 
    0.05986007, 0.05987716, 0.05983182, 0.05984269, 0.05982916, 0.05983603, 
    0.05982434, 0.05983486, 0.05981643, 0.05981253, 0.05981522, 0.05980449, 
    0.05983547, 0.05982375, 0.05991199, 0.05991149, 0.05990904, 0.05991982, 
    0.05992042, 0.05992994, 0.05992137, 0.0599178, 0.0599083, 0.05990285, 
    0.0598976, 0.05988599, 0.05987325, 0.05985519, 0.05984201, 0.05983316, 
    0.05983852, 0.0598338, 0.05983911, 0.05984155, 0.05981406, 0.05982963, 
    0.05980604, 0.05980731, 0.0598181, 0.05980717, 0.05991112, 0.05991403, 
    0.05992443, 0.0599163, 0.05993096, 0.05992289, 0.05991832, 0.0599, 
    0.0598957, 0.05989204, 0.05988455, 0.0598751, 0.05985868, 0.05984417, 
    0.05983068, 0.05983165, 0.05983132, 0.05982841, 0.05983577, 0.05982719, 
    0.05982585, 0.05982951, 0.05980749, 0.05981379, 0.05980734, 0.05981142, 
    0.05991306, 0.05990811, 0.0599108, 0.0599058, 0.05990941, 0.05989362, 
    0.05988888, 0.05986645, 0.05987535, 0.05986089, 0.05987379, 0.05987157, 
    0.05986086, 0.05987303, 0.05984517, 0.05986448, 0.05982829, 0.05984813, 
    0.05982707, 0.05983074, 0.05982455, 0.05981911, 0.05981204, 0.05979925, 
    0.05980217, 0.05979126, 0.05990063, 0.05989427, 0.05989464, 0.05988783, 
    0.05988283, 0.05987184, 0.05985446, 0.05986095, 0.05984882, 0.05984645, 
    0.05986475, 0.05985371, 0.05988986, 0.05988419, 0.05988742, 0.05990024, 
    0.05985972, 0.05988055, 0.05984182, 0.05985313, 0.05981991, 0.0598367, 
    0.05980383, 0.05979015, 0.05977625, 0.05976101, 0.05989058, 0.05989493, 
    0.05988697, 0.05987632, 0.05986597, 0.05985247, 0.05985098, 0.05984851, 
    0.05984184, 0.05983631, 0.05984791, 0.0598349, 0.05988327, 0.05985782, 
    0.05989676, 0.05988524, 0.05987686, 0.05988031, 0.05986164, 0.05985729, 
    0.05983965, 0.05984867, 0.05979371, 0.05981823, 0.05974865, 0.05976845, 
    0.0598965, 0.05989051, 0.05987, 0.05987967, 0.05985147, 0.05984458, 
    0.05983879, 0.0598317, 0.05983078, 0.05982654, 0.05983351, 0.05982674, 
    0.05985244, 0.05984097, 0.05987209, 0.05986466, 0.05986802, 0.05987183, 
    0.05986005, 0.05984778, 0.0598472, 0.05984331, 0.05983286, 0.05985135, 
    0.05979111, 0.05982907, 0.05988398, 0.05987292, 0.05987096, 0.05987529, 
    0.05984528, 0.05985622, 0.0598266, 0.05983458, 0.0598214, 0.05982799, 
    0.05982897, 0.05983732, 0.05984259, 0.05985578, 0.0598664, 0.05987462, 
    0.05987269, 0.05986364, 0.05984696, 0.05983084, 0.05983443, 0.0598224, 
    0.05985353, 0.0598407, 0.05984577, 0.05983246, 0.05986119, 0.05983771, 
    0.05986727, 0.05986463, 0.05985644, 0.05984004, 0.05983592, 0.05983209, 
    0.05983439, 0.05984647, 0.0598483, 0.05985656, 0.059859, 0.05986518, 
    0.05987044, 0.05986571, 0.05986081, 0.05984633, 0.0598334, 0.05981908, 
    0.05981543, 0.05979936, 0.0598129, 0.05979097, 0.0598103, 0.0597764, 
    0.05983588, 0.05981021, 0.05985596, 0.059851, 0.05984235, 0.05982166, 
    0.05983252, 0.05981966, 0.05984835, 0.05986349, 0.05986699, 0.05987418, 
    0.05986683, 0.05986742, 0.05986038, 0.05986262, 0.05984585, 0.05985485, 
    0.05982908, 0.05981968, 0.05979252, 0.05977591, 0.05975834, 0.05975072, 
    0.05974837, 0.0597474 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.78002, 3.793108, 3.790562, 3.801136, 3.795269, 3.802197, 3.782672, 
    3.793626, 3.786632, 3.781199, 3.821721, 3.801609, 3.842721, 3.829824, 
    3.862291, 3.840709, 3.866655, 3.861671, 3.876696, 3.872387, 3.891646, 
    3.878686, 3.901665, 3.888551, 3.890598, 3.878258, 3.805654, 3.819211, 
    3.804851, 3.806782, 3.805916, 3.795389, 3.79009, 3.779024, 3.781032, 
    3.789162, 3.80765, 3.801369, 3.817224, 3.816865, 3.834575, 3.826582, 
    3.856449, 3.847942, 3.872567, 3.866362, 3.872275, 3.870482, 3.872298, 
    3.863201, 3.867096, 3.8591, 3.828077, 3.837173, 3.810094, 3.79388, 
    3.783152, 3.775551, 3.776624, 3.778671, 3.789209, 3.799143, 3.806725, 
    3.811804, 3.816814, 3.831999, 3.840066, 3.858168, 3.8549, 3.860441, 
    3.865745, 3.874659, 3.873191, 3.877121, 3.860297, 3.871471, 3.853039, 
    3.858073, 3.818162, 3.803063, 3.796648, 3.79105, 3.77745, 3.786837, 
    3.783134, 3.791952, 3.797561, 3.794787, 3.811943, 3.805265, 3.840544, 
    3.825316, 3.865126, 3.855571, 3.86742, 3.861371, 3.871739, 3.862407, 
    3.878586, 3.882114, 3.879703, 3.888978, 3.86189, 3.872273, 3.794708, 
    3.795161, 3.79727, 3.788004, 3.787439, 3.778969, 3.786506, 3.789718, 
    3.797888, 3.802725, 3.807328, 3.817465, 3.82881, 3.844723, 3.85619, 
    3.863891, 3.859168, 3.863337, 3.858676, 3.856494, 3.880791, 3.867132, 
    3.887643, 3.886506, 3.877214, 3.886634, 3.795479, 3.792876, 3.783845, 
    3.790911, 3.778047, 3.785241, 3.789382, 3.805401, 3.808932, 3.812203, 
    3.818674, 3.82699, 3.841613, 3.854374, 3.866055, 3.865198, 3.8655, 
    3.868111, 3.861643, 3.869174, 3.870437, 3.867132, 3.886354, 3.880855, 
    3.886482, 3.882901, 3.793722, 3.798104, 3.795735, 3.80019, 3.79705, 
    3.811023, 3.815221, 3.834915, 3.826826, 3.83971, 3.828134, 3.830182, 
    3.840125, 3.82876, 3.853667, 3.836761, 3.868212, 3.851275, 3.869276, 
    3.866004, 3.871423, 3.87628, 3.8824, 3.893707, 3.891087, 3.900559, 
    3.804646, 3.810343, 3.809843, 3.815814, 3.820233, 3.82983, 3.845258, 
    3.839452, 3.85012, 3.852264, 3.836059, 3.845999, 3.814161, 3.819288, 
    3.816236, 3.805094, 3.840785, 3.822433, 3.856379, 3.846397, 3.875587, 
    3.861046, 3.889644, 3.901913, 3.913499, 3.927058, 3.813457, 3.809583, 
    3.816525, 3.826141, 3.835088, 3.847005, 3.848227, 3.850462, 3.856261, 
    3.86114, 3.851167, 3.862365, 3.820472, 3.842383, 3.808117, 3.818405, 
    3.825575, 3.822431, 3.838789, 3.842652, 3.858378, 3.850244, 3.89888, 
    3.877303, 3.937414, 3.920543, 3.808229, 3.813445, 3.831639, 3.822974, 
    3.847803, 3.853932, 3.858924, 3.865307, 3.865998, 3.869785, 3.863581, 
    3.869541, 3.84703, 3.857077, 3.829559, 3.836241, 3.833167, 3.829795, 
    3.840209, 3.851323, 3.851565, 3.855134, 3.865197, 3.847903, 3.901664, 
    3.868387, 3.819139, 3.829208, 3.830653, 3.826748, 3.853317, 3.843673, 
    3.869694, 3.862648, 3.874198, 3.868455, 3.86761, 3.860246, 3.855666, 
    3.844114, 3.834736, 3.827315, 3.82904, 3.837195, 3.852005, 3.866059, 
    3.862976, 3.873319, 3.845998, 3.857434, 3.853009, 3.864555, 3.839296, 
    3.860784, 3.833818, 3.836177, 3.843482, 3.858207, 3.861478, 3.864964, 
    3.862813, 3.852382, 3.850677, 3.843305, 3.841269, 3.835664, 3.831025, 
    3.835262, 3.839714, 3.852388, 3.863836, 3.876348, 3.879417, 3.894075, 
    3.882134, 3.901849, 3.885074, 3.914152, 3.862039, 3.88459, 3.843816, 
    3.848193, 3.856116, 3.874346, 3.864501, 3.876019, 3.850611, 3.837475, 
    3.834087, 3.827765, 3.834232, 3.833706, 3.839902, 3.83791, 3.85281, 
    3.844801, 3.867588, 3.875929, 3.899564, 3.914106, 3.928957, 3.935525, 
    3.937526, 3.938362,
  3.295895, 3.308631, 3.306154, 3.316445, 3.310736, 3.317477, 3.298478, 
    3.309134, 3.30233, 3.297045, 3.336163, 3.316905, 3.356097, 3.343864, 
    3.374674, 3.354186, 3.378819, 3.374091, 3.388361, 3.384268, 3.402553, 
    3.390251, 3.412076, 3.399617, 3.40156, 3.389844, 3.320845, 3.333782, 
    3.320063, 3.321941, 3.3211, 3.310851, 3.305691, 3.294929, 3.296882, 
    3.30479, 3.322786, 3.316674, 3.331913, 3.331573, 3.348372, 3.340789, 
    3.369133, 3.361059, 3.384439, 3.378546, 3.384161, 3.382458, 3.384183, 
    3.375543, 3.379242, 3.371651, 3.342206, 3.350835, 3.325147, 3.309377, 
    3.298943, 3.291549, 3.292593, 3.294584, 3.304837, 3.314507, 3.321889, 
    3.326771, 3.331524, 3.345918, 3.353577, 3.370763, 3.367664, 3.372921, 
    3.37796, 3.386424, 3.385031, 3.388762, 3.372788, 3.383395, 3.365898, 
    3.370675, 3.332786, 3.318323, 3.312072, 3.306629, 3.293396, 3.302528, 
    3.298925, 3.307508, 3.312968, 3.310268, 3.326903, 3.320467, 3.354032, 
    3.339586, 3.377372, 3.3683, 3.379551, 3.373808, 3.38365, 3.374791, 
    3.390154, 3.393503, 3.391214, 3.400026, 3.3743, 3.384157, 3.310191, 
    3.310631, 3.312685, 3.303664, 3.303114, 3.294874, 3.302208, 3.305332, 
    3.313286, 3.317993, 3.322474, 3.33214, 3.342899, 3.358, 3.368887, 3.3762, 
    3.371716, 3.375674, 3.371249, 3.369178, 3.392246, 3.379275, 3.398757, 
    3.397678, 3.38885, 3.3978, 3.31094, 3.308408, 3.299618, 3.306495, 
    3.293978, 3.300976, 3.305004, 3.320596, 3.324037, 3.327149, 3.333288, 
    3.341176, 3.355049, 3.367162, 3.378255, 3.377442, 3.377728, 3.380206, 
    3.374065, 3.381216, 3.382414, 3.379277, 3.397533, 3.39231, 3.397655, 
    3.394254, 3.309232, 3.313496, 3.311191, 3.315525, 3.312469, 3.326026, 
    3.330006, 3.34869, 3.341019, 3.353242, 3.342262, 3.344203, 3.353628, 
    3.342856, 3.366488, 3.35044, 3.380303, 3.364213, 3.381312, 3.378207, 
    3.383353, 3.387964, 3.393777, 3.404515, 3.402028, 3.411028, 3.319864, 
    3.325382, 3.324913, 3.330574, 3.334765, 3.343871, 3.35851, 3.353001, 
    3.363127, 3.365161, 3.349782, 3.359212, 3.329005, 3.333864, 3.330974, 
    3.320298, 3.354262, 3.336848, 3.369066, 3.359592, 3.387305, 3.373494, 
    3.400657, 3.412307, 3.423327, 3.436209, 3.328339, 3.324666, 3.33125, 
    3.340366, 3.348859, 3.360168, 3.36133, 3.363451, 3.368957, 3.373589, 
    3.364116, 3.374751, 3.33498, 3.355779, 3.323241, 3.333026, 3.339831, 
    3.33685, 3.352373, 3.356038, 3.370963, 3.363244, 3.409424, 3.38893, 
    3.446062, 3.430017, 3.323353, 3.328329, 3.345584, 3.337366, 3.360927, 
    3.366744, 3.371485, 3.377542, 3.378201, 3.381795, 3.375906, 3.381565, 
    3.360192, 3.36973, 3.343615, 3.349953, 3.347038, 3.343839, 3.35372, 
    3.364263, 3.364498, 3.367883, 3.37742, 3.361023, 3.412059, 3.380452, 
    3.33373, 3.343275, 3.344651, 3.340948, 3.36616, 3.357006, 3.381709, 
    3.375021, 3.385988, 3.380533, 3.379731, 3.37274, 3.36839, 3.357424, 
    3.348524, 3.341486, 3.343122, 3.350858, 3.364912, 3.378256, 3.375328, 
    3.385153, 3.359214, 3.370066, 3.365865, 3.37683, 3.352853, 3.373234, 
    3.347656, 3.349894, 3.356825, 3.370797, 3.373909, 3.377217, 3.375177, 
    3.365271, 3.363654, 3.356658, 3.354724, 3.349407, 3.345006, 3.349025, 
    3.353248, 3.365278, 3.376145, 3.388028, 3.390945, 3.404857, 3.393516, 
    3.412234, 3.396296, 3.423933, 3.374432, 3.395846, 3.357144, 3.361298, 
    3.368814, 3.386121, 3.376778, 3.387711, 3.363591, 3.35112, 3.347911, 
    3.341912, 3.348049, 3.347549, 3.353429, 3.351539, 3.365679, 3.358078, 
    3.379709, 3.387627, 3.410081, 3.423898, 3.438022, 3.444267, 3.446171, 
    3.446966,
  3.020731, 3.03483, 3.032086, 3.043485, 3.037158, 3.044627, 3.023586, 
    3.035391, 3.027851, 3.021999, 3.065695, 3.043994, 3.08836, 3.074431, 
    3.109509, 3.086189, 3.114136, 3.108835, 3.12466, 3.120142, 3.140349, 
    3.126747, 3.150863, 3.137097, 3.139247, 3.126299, 3.048353, 3.062987, 
    3.047487, 3.049571, 3.048636, 3.037288, 3.031581, 3.019656, 3.021819, 
    3.030579, 3.050508, 3.043732, 3.06083, 3.060443, 3.079559, 3.07093, 
    3.10319, 3.093996, 3.120331, 3.113827, 3.120025, 3.118145, 3.120049, 
    3.11049, 3.114597, 3.106056, 3.072544, 3.082365, 3.053142, 3.035667, 
    3.024103, 3.015916, 3.017072, 3.019278, 3.03063, 3.041332, 3.049507, 
    3.054984, 3.060388, 3.076786, 3.085492, 3.105051, 3.101515, 3.107507, 
    3.11318, 3.122525, 3.120986, 3.125108, 3.107349, 3.119184, 3.099502, 
    3.104945, 3.061856, 3.045559, 3.03865, 3.032613, 3.017962, 3.028074, 
    3.024085, 3.033582, 3.039628, 3.036637, 3.055134, 3.047933, 3.086009, 
    3.069566, 3.112532, 3.102241, 3.114935, 3.10851, 3.119464, 3.10963, 
    3.126643, 3.130345, 3.127815, 3.137544, 3.109071, 3.120025, 3.036553, 
    3.037041, 3.039314, 3.029331, 3.028722, 3.019597, 3.027715, 3.031177, 
    3.039979, 3.045194, 3.050158, 3.061092, 3.073337, 3.090521, 3.10291, 
    3.111234, 3.106128, 3.110636, 3.105597, 3.103237, 3.128957, 3.114635, 
    3.136143, 3.13495, 3.125205, 3.135085, 3.037383, 3.034577, 3.024849, 
    3.03246, 3.018604, 3.026354, 3.030817, 3.048083, 3.051887, 3.055416, 
    3.062396, 3.071371, 3.087161, 3.100949, 3.113504, 3.112606, 3.112922, 
    3.11566, 3.108804, 3.116774, 3.1181, 3.114634, 3.13479, 3.129022, 
    3.134925, 3.131168, 3.035489, 3.040213, 3.03766, 3.042462, 3.039078, 
    3.054146, 3.058674, 3.07993, 3.071194, 3.085106, 3.072605, 3.074817, 
    3.08556, 3.07328, 3.100187, 3.081925, 3.115767, 3.097605, 3.116881, 
    3.113451, 3.119131, 3.124225, 3.130642, 3.142508, 3.139758, 3.1497, 
    3.047265, 3.05341, 3.052869, 3.059309, 3.064079, 3.074435, 3.091098, 
    3.084824, 3.096349, 3.098666, 3.08116, 3.0919, 3.057528, 3.063062, 
    3.059767, 3.047749, 3.086268, 3.066456, 3.103114, 3.092327, 3.123498, 
    3.108162, 3.138244, 3.151127, 3.16329, 3.177544, 3.056768, 3.052588, 
    3.060076, 3.070457, 3.080113, 3.092984, 3.094304, 3.09672, 3.102985, 
    3.10826, 3.097484, 3.109584, 3.064346, 3.087993, 3.051009, 3.062111, 
    3.069845, 3.066451, 3.084108, 3.08828, 3.105277, 3.096482, 3.147943, 
    3.125301, 3.188432, 3.170695, 3.051129, 3.056754, 3.076391, 3.067036, 
    3.093845, 3.10047, 3.105863, 3.112722, 3.113446, 3.117415, 3.110899, 
    3.117159, 3.093012, 3.103868, 3.074142, 3.081358, 3.078037, 3.074397, 
    3.085641, 3.097653, 3.097911, 3.10177, 3.112618, 3.093954, 3.150872, 
    3.11596, 3.062897, 3.073769, 3.075325, 3.071108, 3.099805, 3.089385, 
    3.117319, 3.109891, 3.122041, 3.11602, 3.115135, 3.107294, 3.102343, 
    3.089862, 3.079733, 3.071719, 3.073581, 3.082389, 3.098389, 3.11351, 
    3.110248, 3.121119, 3.091895, 3.104255, 3.099474, 3.111933, 3.084657, 
    3.107888, 3.07874, 3.081287, 3.089178, 3.105095, 3.108625, 3.112363, 
    3.110069, 3.098796, 3.096952, 3.088986, 3.086789, 3.080733, 3.075725, 
    3.0803, 3.08511, 3.098801, 3.111177, 3.124297, 3.127514, 3.142901, 
    3.13037, 3.151067, 3.133462, 3.163985, 3.109239, 3.132947, 3.089538, 
    3.094267, 3.102834, 3.122201, 3.111876, 3.123954, 3.09688, 3.082693, 
    3.079031, 3.072206, 3.079187, 3.078619, 3.08531, 3.083158, 3.099257, 
    3.090602, 3.115113, 3.123858, 3.148657, 3.16393, 3.179536, 3.186443, 
    3.188547, 3.189427,
  2.893865, 2.909182, 2.906199, 2.91859, 2.911711, 2.919832, 2.896965, 
    2.909792, 2.901598, 2.895241, 2.942754, 2.919143, 2.967429, 2.952258, 
    2.990482, 2.965065, 2.995516, 2.989746, 3.006982, 3.002058, 3.024093, 
    3.009256, 3.035564, 3.020544, 3.02289, 3.008768, 2.923882, 2.939806, 
    2.922941, 2.925207, 2.92419, 2.911854, 2.905653, 2.892696, 2.895045, 
    2.904562, 2.926226, 2.918858, 2.937454, 2.937033, 2.957842, 2.948445, 
    2.98359, 2.973568, 3.002263, 2.995177, 3.00193, 2.999881, 3.001957, 
    2.99155, 2.996017, 2.986714, 2.950204, 2.960898, 2.929091, 2.910094, 
    2.897527, 2.888635, 2.889891, 2.892286, 2.904618, 2.916249, 2.925137, 
    2.931094, 2.936972, 2.954825, 2.964305, 2.98562, 2.981764, 2.988298, 
    2.994473, 3.004655, 3.002977, 3.00747, 2.988125, 3.001014, 2.979569, 
    2.985503, 2.938576, 2.920844, 2.913336, 2.906773, 2.890857, 2.901841, 
    2.897507, 2.907825, 2.914396, 2.911145, 2.931257, 2.923425, 2.964868, 
    2.946962, 2.993767, 2.982555, 2.996385, 2.989389, 3.00132, 2.990611, 
    3.009143, 3.01318, 3.010421, 3.021029, 2.990002, 3.001931, 2.911054, 
    2.911584, 2.914054, 2.903207, 2.902544, 2.892632, 2.901451, 2.905212, 
    2.914777, 2.920447, 2.925845, 2.937739, 2.951068, 2.969783, 2.983284, 
    2.992355, 2.986792, 2.991708, 2.986213, 2.98364, 3.011667, 2.996058, 
    3.019502, 3.018201, 3.007577, 3.018347, 2.911956, 2.908906, 2.898338, 
    2.906606, 2.891554, 2.899973, 2.904822, 2.923589, 2.927724, 2.931564, 
    2.939157, 2.948926, 2.966122, 2.981147, 2.994825, 2.993847, 2.994191, 
    2.997175, 2.989711, 2.998388, 2.999833, 2.996056, 3.018027, 3.011737, 
    3.018173, 3.014076, 2.909897, 2.915032, 2.912256, 2.917477, 2.913799, 
    2.930184, 2.935111, 2.958247, 2.948733, 2.963884, 2.950269, 2.952678, 
    2.964381, 2.951004, 2.980318, 2.960421, 2.99729, 2.977504, 2.998504, 
    2.994767, 3.000956, 3.006508, 3.013503, 3.026446, 3.023445, 3.034294, 
    2.922699, 2.929383, 2.928793, 2.935799, 2.940989, 2.952261, 2.970411, 
    2.963575, 2.976132, 2.978658, 2.959584, 2.971285, 2.933862, 2.939885, 
    2.936297, 2.923226, 2.96515, 2.943578, 2.983508, 2.97175, 3.005716, 
    2.989012, 3.021794, 3.035853, 3.049129, 3.064706, 2.933035, 2.928488, 
    2.936633, 2.947933, 2.958445, 2.972466, 2.973903, 2.976537, 2.983366, 
    2.989118, 2.977371, 2.990561, 2.941284, 2.967028, 2.926771, 2.938849, 
    2.947265, 2.94357, 2.962795, 2.96734, 2.985866, 2.976277, 3.032379, 
    3.007683, 3.076607, 3.057221, 2.9269, 2.933019, 2.954392, 2.944208, 
    2.973403, 2.980625, 2.986504, 2.993974, 2.994761, 2.999087, 2.991996, 
    2.998807, 2.972496, 2.984329, 2.951942, 2.9598, 2.956183, 2.952219, 
    2.964465, 2.977556, 2.977834, 2.982042, 2.993869, 2.973522, 3.035581, 
    2.997508, 2.939702, 2.951538, 2.95323, 2.948639, 2.9799, 2.968544, 
    2.998981, 2.990896, 3.004127, 2.997567, 2.996603, 2.988064, 2.982667, 
    2.969064, 2.958031, 2.949305, 2.951332, 2.960924, 2.978358, 2.994833, 
    2.991287, 3.003123, 2.971279, 2.984752, 2.97954, 2.993114, 2.963394, 
    2.988719, 2.956948, 2.959723, 2.968319, 2.985669, 2.989516, 2.993583, 
    2.99109, 2.978801, 2.976791, 2.968109, 2.965717, 2.959118, 2.953665, 
    2.958648, 2.963887, 2.978806, 2.992295, 3.006587, 3.010092, 3.026879, 
    3.01321, 3.035794, 3.016587, 3.049895, 2.990189, 3.016021, 2.96871, 
    2.973863, 2.983203, 3.004304, 2.993052, 3.006214, 2.976712, 2.961256, 
    2.957266, 2.949835, 2.957436, 2.956817, 2.964104, 2.961761, 2.979302, 
    2.969869, 2.996579, 3.00611, 3.033156, 3.049832, 3.06688, 3.074431, 
    3.076732, 3.077694,
  2.944312, 2.960424, 2.957285, 2.970329, 2.963086, 2.971637, 2.947571, 
    2.961066, 2.952444, 2.945758, 2.995805, 2.970912, 3.021869, 3.005837, 
    3.046266, 3.01937, 3.051717, 3.045485, 3.064275, 3.058881, 3.082962, 
    3.066768, 3.095155, 3.079147, 3.081684, 3.066233, 2.975904, 2.992695, 
    2.974912, 2.9773, 2.976228, 2.963236, 2.95671, 2.943083, 2.945552, 
    2.955562, 2.978375, 2.970611, 2.990212, 2.989768, 3.011735, 3.001812, 
    3.038966, 3.028361, 3.059106, 3.051345, 3.058741, 3.056496, 3.05877, 
    3.047397, 3.052265, 3.042274, 3.003668, 3.014965, 2.981394, 2.961385, 
    2.948162, 2.938815, 2.940135, 2.942652, 2.955621, 2.967863, 2.977226, 
    2.983505, 2.989704, 3.008549, 3.018566, 3.041116, 3.037033, 3.043952, 
    3.050574, 3.061726, 3.059887, 3.064811, 3.043768, 3.057738, 3.03471, 
    3.040992, 2.991397, 2.972703, 2.964796, 2.957888, 2.94115, 2.952699, 
    2.948141, 2.958995, 2.965913, 2.962489, 2.983677, 2.975423, 3.019161, 
    3.000246, 3.049801, 3.037871, 3.052667, 3.045108, 3.058072, 3.046402, 
    3.066644, 3.07107, 3.068045, 3.079679, 3.045757, 3.058741, 2.962394, 
    2.962952, 2.965553, 2.954137, 2.953439, 2.943016, 2.952288, 2.956246, 
    2.966314, 2.972285, 2.977972, 2.990513, 3.00458, 3.024357, 3.038643, 
    3.048255, 3.042357, 3.047564, 3.041744, 3.03902, 3.069412, 3.05231, 
    3.078003, 3.076576, 3.064928, 3.076737, 2.963344, 2.960133, 2.949014, 
    2.957712, 2.941883, 2.950734, 2.955835, 2.975596, 2.979954, 2.984001, 
    2.99201, 3.002319, 3.020487, 3.036381, 3.05096, 3.049889, 3.050266, 
    3.053532, 3.045449, 3.054861, 3.056444, 3.052308, 3.076385, 3.069487, 
    3.076546, 3.072052, 2.961176, 2.966582, 2.96366, 2.969157, 2.965284, 
    2.982547, 2.987741, 3.012163, 3.002116, 3.018121, 3.003737, 3.006281, 
    3.018646, 3.004513, 3.035503, 3.014461, 3.053659, 3.032526, 3.054988, 
    3.050897, 3.057673, 3.063756, 3.071424, 3.085462, 3.082273, 3.093804, 
    2.974658, 2.981702, 2.98108, 2.988467, 2.993942, 3.005841, 3.025021, 
    3.017794, 3.031074, 3.033746, 3.013577, 3.025946, 2.986425, 2.992777, 
    2.988992, 2.975213, 3.019459, 2.996674, 3.03888, 3.026438, 3.062888, 
    3.044709, 3.080518, 3.095463, 3.109589, 3.126186, 2.985552, 2.980758, 
    2.989347, 3.001271, 3.012372, 3.027195, 3.028715, 3.031502, 3.03873, 
    3.04482, 3.032384, 3.046349, 2.994254, 3.021445, 2.978948, 2.991685, 
    3.000566, 2.996666, 3.016969, 3.021774, 3.041377, 3.031227, 3.091769, 
    3.065044, 3.13888, 3.118207, 2.979085, 2.985535, 3.008091, 2.997339, 
    3.028187, 3.035828, 3.042052, 3.050029, 3.05089, 3.055627, 3.047869, 
    3.05532, 3.027227, 3.03975, 3.005503, 3.013805, 3.009983, 3.005797, 
    3.018735, 3.03258, 3.032875, 3.037328, 3.049915, 3.028312, 3.095174, 
    3.053899, 2.992584, 3.005077, 3.006864, 3.002016, 3.035061, 3.023047, 
    3.055511, 3.046704, 3.061147, 3.053962, 3.052906, 3.043704, 3.037989, 
    3.023597, 3.011936, 3.002718, 3.004859, 3.014992, 3.033428, 3.050969, 
    3.047118, 3.060047, 3.02594, 3.040197, 3.034679, 3.049087, 3.017603, 
    3.044398, 3.010791, 3.013723, 3.022809, 3.041168, 3.045241, 3.0496, 
    3.04691, 3.033898, 3.03177, 3.022588, 3.020058, 3.013084, 3.007323, 
    3.012587, 3.018124, 3.033902, 3.048191, 3.063843, 3.067685, 3.085922, 
    3.071104, 3.095401, 3.074808, 3.110406, 3.045956, 3.074187, 3.023223, 
    3.028673, 3.038557, 3.061342, 3.049019, 3.063435, 3.031687, 3.015343, 
    3.011127, 3.003278, 3.011307, 3.010653, 3.018353, 3.015876, 3.034428, 
    3.024449, 3.05288, 3.06332, 3.092594, 3.110337, 3.128503, 3.136557, 
    3.139013, 3.14004,
  2.969938, 2.988338, 2.98475, 2.999671, 2.991382, 3.001169, 2.973656, 
    2.989072, 2.979219, 2.971587, 3.028894, 3.000339, 3.058904, 3.040431, 
    3.087099, 3.056021, 3.093413, 3.086195, 3.107979, 3.101718, 3.129798, 
    3.110874, 3.144477, 3.125264, 3.128261, 3.110252, 3.006057, 3.025321, 
    3.00492, 3.007657, 3.006428, 2.991553, 2.984093, 2.968536, 2.971352, 
    2.982781, 3.008888, 2.999994, 3.022469, 3.021959, 3.047222, 3.0358, 
    3.078652, 3.066396, 3.101979, 3.092982, 3.101557, 3.098953, 3.10159, 
    3.088408, 3.094048, 3.082479, 3.037935, 3.050943, 3.01235, 2.989436, 
    2.97433, 2.963669, 2.965173, 2.968044, 2.982848, 2.996848, 3.007572, 
    3.014771, 3.021886, 3.043553, 3.055095, 3.081139, 3.076417, 3.084421, 
    3.092089, 3.10502, 3.102887, 3.108601, 3.084208, 3.100393, 3.073731, 
    3.080995, 3.02383, 3.00239, 2.993339, 2.985439, 2.966331, 2.979511, 
    2.974307, 2.986705, 2.994616, 2.9907, 3.014969, 3.005505, 3.05578, 
    3.033998, 3.091193, 3.077385, 3.094514, 3.085758, 3.100781, 3.087257, 
    3.11073, 3.115872, 3.112357, 3.125884, 3.086509, 3.101557, 2.99059, 
    2.991229, 2.994204, 2.981153, 2.980356, 2.968459, 2.979042, 2.983563, 
    2.995075, 3.001911, 3.008427, 3.022815, 3.038985, 3.061775, 3.078278, 
    3.089403, 3.082575, 3.088602, 3.081866, 3.078714, 3.113945, 3.094101, 
    3.123934, 3.122273, 3.108737, 3.12246, 2.991677, 2.988005, 2.975303, 
    2.985238, 2.967166, 2.977267, 2.983093, 3.005704, 3.010698, 3.015341, 
    3.024534, 3.036383, 3.057309, 3.075662, 3.092536, 3.091295, 3.091732, 
    3.095517, 3.086153, 3.097057, 3.098893, 3.094098, 3.122051, 3.114032, 
    3.122238, 3.117013, 2.989198, 2.995382, 2.992038, 2.998329, 2.993896, 
    3.013672, 3.019632, 3.047715, 3.03615, 3.05458, 3.038015, 3.040942, 
    3.055187, 3.038907, 3.074648, 3.050362, 3.095664, 3.071208, 3.097205, 
    3.092462, 3.100318, 3.107376, 3.116283, 3.132805, 3.128969, 3.142848, 
    3.004628, 3.012703, 3.01199, 3.020466, 3.026753, 3.040435, 3.062541, 
    3.054204, 3.069529, 3.072618, 3.049343, 3.063608, 3.018121, 3.025415, 
    3.021069, 3.005265, 3.056125, 3.029892, 3.078552, 3.064176, 3.106369, 
    3.085296, 3.12686, 3.144848, 3.161419, 3.180853, 3.01712, 3.011621, 
    3.021475, 3.035177, 3.047956, 3.06505, 3.066805, 3.070024, 3.078378, 
    3.085426, 3.071044, 3.087195, 3.027112, 3.058414, 3.009546, 3.024161, 
    3.034367, 3.029883, 3.053253, 3.058794, 3.08144, 3.069707, 3.140397, 
    3.108872, 3.195752, 3.171504, 3.009703, 3.017101, 3.043026, 3.030656, 
    3.066195, 3.075023, 3.082222, 3.091457, 3.092455, 3.097945, 3.088955, 
    3.097589, 3.065087, 3.079558, 3.040047, 3.049606, 3.045204, 3.040385, 
    3.055289, 3.07127, 3.07161, 3.076758, 3.091325, 3.06634, 3.1445, 
    3.095942, 3.025193, 3.039557, 3.041613, 3.036035, 3.074136, 3.060263, 
    3.097811, 3.087606, 3.104348, 3.096014, 3.094791, 3.084134, 3.077522, 
    3.060898, 3.047453, 3.036843, 3.039306, 3.050975, 3.07225, 3.092546, 
    3.088086, 3.103072, 3.063601, 3.080076, 3.073696, 3.090366, 3.053984, 
    3.084937, 3.046134, 3.049512, 3.059988, 3.081199, 3.085913, 3.090961, 
    3.087844, 3.072792, 3.070334, 3.059732, 3.056814, 3.048776, 3.042142, 
    3.048203, 3.054585, 3.072798, 3.089328, 3.107477, 3.111938, 3.133359, 
    3.115911, 3.144773, 3.120218, 3.162374, 3.08674, 3.119495, 3.060465, 
    3.066756, 3.078179, 3.104575, 3.090287, 3.107003, 3.070238, 3.051379, 
    3.046521, 3.037487, 3.046728, 3.045975, 3.054848, 3.051993, 3.073405, 
    3.06188, 3.094761, 3.10687, 3.141391, 3.162294, 3.18357, 3.193024, 
    3.195909, 3.197116,
  3.254741, 3.278218, 3.27363, 3.292737, 3.282113, 3.29466, 3.259476, 
    3.279157, 3.266568, 3.256841, 3.329907, 3.293594, 3.367681, 3.34439, 
    3.403476, 3.364038, 3.411533, 3.402324, 3.430179, 3.422155, 3.458265, 
    3.433895, 3.477267, 3.452414, 3.45628, 3.433097, 3.300939, 3.325432, 
    3.299479, 3.302996, 3.301416, 3.282333, 3.272791, 3.252957, 3.256542, 
    3.271116, 3.30458, 3.293151, 3.321862, 3.321224, 3.352938, 3.33857, 
    3.392721, 3.377164, 3.422489, 3.410983, 3.421947, 3.418616, 3.421991, 
    3.405146, 3.412344, 3.397591, 3.341253, 3.357629, 3.309036, 3.279623, 
    3.260335, 3.24677, 3.248682, 3.252332, 3.271201, 3.289116, 3.302887, 
    3.312155, 3.321133, 3.348318, 3.362868, 3.395885, 3.389879, 3.400063, 
    3.409842, 3.426385, 3.423651, 3.430977, 3.399792, 3.420458, 3.386468, 
    3.395701, 3.323565, 3.296227, 3.284619, 3.274511, 3.250153, 3.266941, 
    3.260305, 3.276129, 3.286255, 3.28124, 3.31241, 3.30023, 3.363734, 
    3.336309, 3.408699, 3.39111, 3.41294, 3.401767, 3.420955, 3.403677, 
    3.43371, 3.440318, 3.4358, 3.453213, 3.402724, 3.421948, 3.2811, 
    3.281917, 3.285727, 3.269036, 3.268019, 3.25286, 3.266342, 3.272114, 
    3.286843, 3.295613, 3.303987, 3.322295, 3.342572, 3.371312, 3.392245, 
    3.406414, 3.397712, 3.405393, 3.396809, 3.3928, 3.43784, 3.412412, 
    3.450698, 3.448558, 3.431152, 3.448799, 3.28249, 3.277792, 3.261575, 
    3.274255, 3.251216, 3.264078, 3.271514, 3.300485, 3.306909, 3.312889, 
    3.324445, 3.339303, 3.365666, 3.388921, 3.410413, 3.408829, 3.409386, 
    3.414221, 3.40227, 3.416191, 3.418538, 3.412408, 3.448272, 3.437953, 
    3.448513, 3.441786, 3.279318, 3.287236, 3.282954, 3.291016, 3.285333, 
    3.310739, 3.318315, 3.353559, 3.339009, 3.362219, 3.341353, 3.345033, 
    3.362985, 3.342474, 3.387632, 3.356896, 3.414409, 3.383265, 3.416379, 
    3.410319, 3.420363, 3.429406, 3.440847, 3.462151, 3.457195, 3.475155, 
    3.299103, 3.309491, 3.308573, 3.319357, 3.327225, 3.344395, 3.372282, 
    3.361744, 3.381135, 3.385054, 3.355611, 3.373633, 3.316427, 3.325549, 
    3.320111, 3.299921, 3.364169, 3.331158, 3.392593, 3.374351, 3.428114, 
    3.401179, 3.454473, 3.477749, 3.499924, 3.526197, 3.315176, 3.308097, 
    3.320619, 3.337789, 3.353863, 3.375459, 3.377682, 3.381763, 3.392373, 
    3.401343, 3.383056, 3.403599, 3.327674, 3.367062, 3.305427, 3.323979, 
    3.336771, 3.331147, 3.360543, 3.367542, 3.396268, 3.38136, 3.471978, 
    3.431325, 3.546064, 3.513538, 3.305628, 3.315152, 3.347654, 3.332116, 
    3.376909, 3.388108, 3.397263, 3.409035, 3.41031, 3.417326, 3.405843, 
    3.41687, 3.375505, 3.393873, 3.343907, 3.355943, 3.350395, 3.344331, 
    3.363113, 3.383343, 3.383775, 3.390312, 3.408867, 3.377093, 3.477297, 
    3.414765, 3.325272, 3.343291, 3.345876, 3.338865, 3.386982, 3.3694, 
    3.417154, 3.404122, 3.425524, 3.414857, 3.413294, 3.399697, 3.391284, 
    3.370203, 3.353229, 3.33988, 3.342975, 3.357669, 3.384588, 3.410426, 
    3.404735, 3.423888, 3.373624, 3.394532, 3.386423, 3.407643, 3.361465, 
    3.400721, 3.351568, 3.355824, 3.369052, 3.395961, 3.401964, 3.408402, 
    3.404426, 3.385276, 3.382156, 3.368729, 3.365041, 3.354896, 3.346541, 
    3.354174, 3.362225, 3.385283, 3.406319, 3.429536, 3.435262, 3.462867, 
    3.440368, 3.477652, 3.44591, 3.501212, 3.403018, 3.44498, 3.369656, 
    3.37762, 3.392119, 3.425814, 3.407542, 3.428928, 3.382034, 3.358179, 
    3.352055, 3.340689, 3.352316, 3.351367, 3.362557, 3.358953, 3.386053, 
    3.371446, 3.413255, 3.428757, 3.473265, 3.501104, 3.529883, 3.542462, 
    3.546271, 3.547866,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016907, 3.972589, 
    4.084889, 4.009923, 4.100391, 4.082681, 4.136661, 4.120984, 4.192374, 
    4.143956, 4.230835, 4.180657, 4.188393, 4.142387, 3.892786, 3.937096, 
    3.890205, 3.896428, 3.893631, 3.860096, 3.843497, 3.80934, 3.815479, 
    3.840594, 3.899235, 3.879052, 3.93047, 3.929288, 3.988761, 3.961638, 
    4.064354, 4.034963, 4.121634, 4.099329, 4.12058, 4.114101, 4.120664, 
    4.088093, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821992, 3.798779, 3.802038, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078353, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077835, 4.117682, 4.052496, 
    4.070027, 3.93363, 3.884468, 3.86409, 3.846481, 3.804549, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085275, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083448, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835237, 3.809173, 3.832339, 3.842323, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023889, 4.06345, 
    4.09053, 4.073862, 4.088568, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846036, 3.806363, 3.828434, 3.841284, 3.891984, 3.903368, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095177, 4.096251, 
    4.105585, 4.082578, 4.109398, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172878, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865339, 
    3.910178, 3.923903, 3.989941, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007906, 3.968978, 4.0547, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226529, 
    3.889542, 3.907957, 3.906323, 3.92583, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937314, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132617, 
    4.080488, 4.184773, 4.231818, 4.277538, 4.332246, 3.918106, 3.905478, 
    3.928167, 3.960172, 3.990517, 4.031764, 4.035937, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941268, 4.015719, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071107, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034485, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971679, 3.994471, 3.98394, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.09525, 4.03483, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975394, 3.962193, 4.053471, 4.020208, 
    4.111266, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021753, 3.989313, 3.964099, 3.969922, 3.997757, 4.048943, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.0678, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994245, 4.019541, 4.070521, 4.081992, 4.094354, 
    4.086712, 4.050242, 4.044355, 4.018919, 4.011842, 3.992481, 3.976649, 
    3.991108, 4.006452, 4.050256, 4.090347, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084012, 4.165855, 4.020701, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044125, 3.99873, 
    3.987085, 3.965621, 3.98758, 3.985781, 4.007088, 4.000206, 4.051713, 
    4.024146, 4.103716, 4.133875, 4.222682, 4.279996, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24813.8, 24834.23, 24830.23, 24846.96, 24837.64, 24848.64, 24817.91, 
    24835.05, 24824.07, 24815.62, 24880.17, 24847.71, 24914.96, 24893.45, 
    24947.95, 24911.58, 24955.42, 24946.88, 24972.81, 24965.31, 24999.27, 
    24976.29, 25017.36, 24993.73, 24997.39, 24975.54, 24854.17, 24876.09, 
    24852.88, 24855.98, 24854.59, 24837.83, 24829.5, 24812.25, 24815.36, 
    24828.04, 24857.38, 24847.32, 24872.83, 24872.25, 24901.32, 24888.11, 
    24938.01, 24923.72, 24965.62, 24954.91, 24965.12, 24962.01, 24965.15, 
    24949.5, 24956.18, 24942.51, 24890.57, 24905.65, 24861.31, 24835.46, 
    24818.65, 24806.9, 24808.55, 24811.71, 24828.11, 24843.78, 24855.89, 
    24864.07, 24872.17, 24897.06, 24910.5, 24940.93, 24935.39, 24944.79, 
    24953.85, 24969.26, 24966.71, 24973.55, 24944.54, 24963.73, 24932.26, 
    24940.76, 24874.39, 24850.02, 24839.83, 24831, 24809.83, 24824.4, 
    24818.63, 24832.41, 24841.27, 24836.88, 24864.3, 24853.55, 24911.3, 
    24886.03, 24952.79, 24936.53, 24956.73, 24946.37, 24964.19, 24948.14, 
    24976.12, 24982.32, 24978.08, 24994.49, 24947.26, 24965.12, 24836.75, 
    24837.47, 24840.8, 24826.22, 24825.34, 24812.17, 24823.88, 24828.9, 
    24841.78, 24849.48, 24856.86, 24873.23, 24891.78, 24918.33, 24937.57, 
    24950.68, 24942.62, 24949.73, 24941.79, 24938.09, 24979.99, 24956.24, 
    24992.11, 24990.09, 24973.72, 24990.32, 24837.97, 24833.86, 24819.73, 
    24830.77, 24810.75, 24821.91, 24828.38, 24853.77, 24859.44, 24864.72, 
    24875.19, 24888.78, 24913.09, 24934.51, 24954.38, 24952.91, 24953.43, 
    24957.92, 24946.84, 24959.75, 24961.94, 24956.23, 24989.82, 24980.1, 
    24990.04, 24983.7, 24835.2, 24842.13, 24838.38, 24845.44, 24840.46, 
    24862.82, 24869.61, 24901.89, 24888.51, 24909.9, 24890.66, 24894.04, 
    24910.61, 24891.69, 24933.33, 24904.97, 24958.1, 24929.31, 24959.93, 
    24954.3, 24963.64, 24972.08, 24982.82, 25002.96, 24998.26, 25015.34, 
    24852.55, 24861.72, 24860.91, 24870.55, 24877.72, 24893.45, 24919.23, 
    24909.46, 24927.36, 24930.96, 24903.79, 24920.49, 24867.89, 24876.2, 
    24871.24, 24853.28, 24911.7, 24881.32, 24937.9, 24921.14, 24970.88, 
    24945.83, 24995.68, 25017.82, 25039.1, 25064.44, 24866.75, 24860.49, 
    24871.7, 24887.39, 24902.17, 24922.16, 24924.19, 24927.93, 24937.69, 
    24945.98, 24929.12, 24948.07, 24878.13, 24914.39, 24858.13, 24874.76, 
    24886.46, 24881.31, 24908.35, 24914.83, 24941.29, 24927.56, 25012.3, 
    24973.88, 25083.95, 25052.28, 24858.31, 24866.73, 24896.45, 24882.2, 
    24923.48, 24933.77, 24942.21, 24953.11, 24954.29, 24960.81, 24950.15, 
    24960.38, 24922.2, 24939.08, 24893.01, 24904.09, 24898.98, 24893.4, 
    24910.73, 24929.38, 24929.78, 24935.79, 24952.95, 24923.65, 25017.38, 
    24958.42, 24875.94, 24892.44, 24894.82, 24888.38, 24932.73, 24916.56, 
    24960.65, 24948.55, 24968.45, 24958.51, 24957.06, 24944.46, 24936.69, 
    24917.3, 24901.59, 24889.31, 24892.15, 24905.69, 24930.53, 24954.39, 
    24949.12, 24966.93, 24920.48, 24939.68, 24932.21, 24951.81, 24909.2, 
    24945.4, 24900.06, 24903.98, 24916.23, 24941, 24946.55, 24952.52, 
    24948.83, 24931.16, 24928.29, 24915.93, 24912.51, 24903.13, 24895.43, 
    24902.46, 24909.9, 24931.17, 24950.59, 24972.21, 24977.57, 25003.63, 
    24982.37, 25017.72, 24987.59, 25040.34, 24947.53, 24986.71, 24916.79, 
    24924.14, 24937.46, 24968.72, 24951.72, 24971.63, 24928.18, 24906.16, 
    24900.51, 24890.05, 24900.75, 24899.87, 24910.21, 24906.88, 24931.88, 
    24918.46, 24957.02, 24971.48, 25013.53, 25040.23, 25067.98, 25080.36, 
    25084.15, 25085.74 ;

 HCSOI =
  24813.8, 24834.23, 24830.23, 24846.96, 24837.64, 24848.64, 24817.91, 
    24835.05, 24824.07, 24815.62, 24880.17, 24847.71, 24914.96, 24893.45, 
    24947.95, 24911.58, 24955.42, 24946.88, 24972.81, 24965.31, 24999.27, 
    24976.29, 25017.36, 24993.73, 24997.39, 24975.54, 24854.17, 24876.09, 
    24852.88, 24855.98, 24854.59, 24837.83, 24829.5, 24812.25, 24815.36, 
    24828.04, 24857.38, 24847.32, 24872.83, 24872.25, 24901.32, 24888.11, 
    24938.01, 24923.72, 24965.62, 24954.91, 24965.12, 24962.01, 24965.15, 
    24949.5, 24956.18, 24942.51, 24890.57, 24905.65, 24861.31, 24835.46, 
    24818.65, 24806.9, 24808.55, 24811.71, 24828.11, 24843.78, 24855.89, 
    24864.07, 24872.17, 24897.06, 24910.5, 24940.93, 24935.39, 24944.79, 
    24953.85, 24969.26, 24966.71, 24973.55, 24944.54, 24963.73, 24932.26, 
    24940.76, 24874.39, 24850.02, 24839.83, 24831, 24809.83, 24824.4, 
    24818.63, 24832.41, 24841.27, 24836.88, 24864.3, 24853.55, 24911.3, 
    24886.03, 24952.79, 24936.53, 24956.73, 24946.37, 24964.19, 24948.14, 
    24976.12, 24982.32, 24978.08, 24994.49, 24947.26, 24965.12, 24836.75, 
    24837.47, 24840.8, 24826.22, 24825.34, 24812.17, 24823.88, 24828.9, 
    24841.78, 24849.48, 24856.86, 24873.23, 24891.78, 24918.33, 24937.57, 
    24950.68, 24942.62, 24949.73, 24941.79, 24938.09, 24979.99, 24956.24, 
    24992.11, 24990.09, 24973.72, 24990.32, 24837.97, 24833.86, 24819.73, 
    24830.77, 24810.75, 24821.91, 24828.38, 24853.77, 24859.44, 24864.72, 
    24875.19, 24888.78, 24913.09, 24934.51, 24954.38, 24952.91, 24953.43, 
    24957.92, 24946.84, 24959.75, 24961.94, 24956.23, 24989.82, 24980.1, 
    24990.04, 24983.7, 24835.2, 24842.13, 24838.38, 24845.44, 24840.46, 
    24862.82, 24869.61, 24901.89, 24888.51, 24909.9, 24890.66, 24894.04, 
    24910.61, 24891.69, 24933.33, 24904.97, 24958.1, 24929.31, 24959.93, 
    24954.3, 24963.64, 24972.08, 24982.82, 25002.96, 24998.26, 25015.34, 
    24852.55, 24861.72, 24860.91, 24870.55, 24877.72, 24893.45, 24919.23, 
    24909.46, 24927.36, 24930.96, 24903.79, 24920.49, 24867.89, 24876.2, 
    24871.24, 24853.28, 24911.7, 24881.32, 24937.9, 24921.14, 24970.88, 
    24945.83, 24995.68, 25017.82, 25039.1, 25064.44, 24866.75, 24860.49, 
    24871.7, 24887.39, 24902.17, 24922.16, 24924.19, 24927.93, 24937.69, 
    24945.98, 24929.12, 24948.07, 24878.13, 24914.39, 24858.13, 24874.76, 
    24886.46, 24881.31, 24908.35, 24914.83, 24941.29, 24927.56, 25012.3, 
    24973.88, 25083.95, 25052.28, 24858.31, 24866.73, 24896.45, 24882.2, 
    24923.48, 24933.77, 24942.21, 24953.11, 24954.29, 24960.81, 24950.15, 
    24960.38, 24922.2, 24939.08, 24893.01, 24904.09, 24898.98, 24893.4, 
    24910.73, 24929.38, 24929.78, 24935.79, 24952.95, 24923.65, 25017.38, 
    24958.42, 24875.94, 24892.44, 24894.82, 24888.38, 24932.73, 24916.56, 
    24960.65, 24948.55, 24968.45, 24958.51, 24957.06, 24944.46, 24936.69, 
    24917.3, 24901.59, 24889.31, 24892.15, 24905.69, 24930.53, 24954.39, 
    24949.12, 24966.93, 24920.48, 24939.68, 24932.21, 24951.81, 24909.2, 
    24945.4, 24900.06, 24903.98, 24916.23, 24941, 24946.55, 24952.52, 
    24948.83, 24931.16, 24928.29, 24915.93, 24912.51, 24903.13, 24895.43, 
    24902.46, 24909.9, 24931.17, 24950.59, 24972.21, 24977.57, 25003.63, 
    24982.37, 25017.72, 24987.59, 25040.34, 24947.53, 24986.71, 24916.79, 
    24924.14, 24937.46, 24968.72, 24951.72, 24971.63, 24928.18, 24906.16, 
    24900.51, 24890.05, 24900.75, 24899.87, 24910.21, 24906.88, 24931.88, 
    24918.46, 24957.02, 24971.48, 25013.53, 25040.23, 25067.98, 25080.36, 
    25084.15, 25085.74 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.356978e-08, 6.384934e-08, 6.379499e-08, 6.402048e-08, 6.389539e-08, 
    6.404304e-08, 6.362645e-08, 6.386044e-08, 6.371106e-08, 6.359494e-08, 
    6.445807e-08, 6.403054e-08, 6.490213e-08, 6.462948e-08, 6.531439e-08, 
    6.485971e-08, 6.540607e-08, 6.530126e-08, 6.561668e-08, 6.552632e-08, 
    6.592977e-08, 6.565838e-08, 6.61389e-08, 6.586495e-08, 6.590781e-08, 
    6.564943e-08, 6.411657e-08, 6.440485e-08, 6.409949e-08, 6.41406e-08, 
    6.412215e-08, 6.389798e-08, 6.378502e-08, 6.354841e-08, 6.359136e-08, 
    6.376514e-08, 6.415908e-08, 6.402535e-08, 6.436237e-08, 6.435476e-08, 
    6.472996e-08, 6.456079e-08, 6.51914e-08, 6.501217e-08, 6.553009e-08, 
    6.539984e-08, 6.552398e-08, 6.548633e-08, 6.552447e-08, 6.533344e-08, 
    6.541529e-08, 6.524719e-08, 6.459248e-08, 6.478489e-08, 6.421101e-08, 
    6.386593e-08, 6.363672e-08, 6.347406e-08, 6.349706e-08, 6.35409e-08, 
    6.376616e-08, 6.397794e-08, 6.413933e-08, 6.42473e-08, 6.435366e-08, 
    6.467567e-08, 6.484608e-08, 6.522765e-08, 6.515878e-08, 6.527544e-08, 
    6.538689e-08, 6.557399e-08, 6.55432e-08, 6.562563e-08, 6.527236e-08, 
    6.550714e-08, 6.511956e-08, 6.522556e-08, 6.438261e-08, 6.406143e-08, 
    6.392494e-08, 6.380544e-08, 6.351474e-08, 6.371549e-08, 6.363636e-08, 
    6.382462e-08, 6.394425e-08, 6.388508e-08, 6.425024e-08, 6.410828e-08, 
    6.485618e-08, 6.453404e-08, 6.537388e-08, 6.517291e-08, 6.542206e-08, 
    6.529492e-08, 6.551276e-08, 6.53167e-08, 6.565631e-08, 6.573026e-08, 
    6.567973e-08, 6.587384e-08, 6.530584e-08, 6.552398e-08, 6.388343e-08, 
    6.389308e-08, 6.393803e-08, 6.374042e-08, 6.372833e-08, 6.354723e-08, 
    6.370837e-08, 6.377699e-08, 6.395118e-08, 6.405422e-08, 6.415217e-08, 
    6.436752e-08, 6.460803e-08, 6.494434e-08, 6.518594e-08, 6.53479e-08, 
    6.524859e-08, 6.533626e-08, 6.523825e-08, 6.519231e-08, 6.570255e-08, 
    6.541605e-08, 6.584592e-08, 6.582213e-08, 6.562759e-08, 6.582481e-08, 
    6.389985e-08, 6.384432e-08, 6.365153e-08, 6.38024e-08, 6.352751e-08, 
    6.368138e-08, 6.376987e-08, 6.411125e-08, 6.418625e-08, 6.425581e-08, 
    6.439316e-08, 6.456945e-08, 6.487869e-08, 6.514775e-08, 6.539337e-08, 
    6.537537e-08, 6.538171e-08, 6.543657e-08, 6.530066e-08, 6.545889e-08, 
    6.548544e-08, 6.541601e-08, 6.581894e-08, 6.570383e-08, 6.582162e-08, 
    6.574668e-08, 6.386237e-08, 6.395581e-08, 6.390532e-08, 6.400027e-08, 
    6.393338e-08, 6.42308e-08, 6.431998e-08, 6.473723e-08, 6.456598e-08, 
    6.483852e-08, 6.459366e-08, 6.463705e-08, 6.484741e-08, 6.460689e-08, 
    6.513292e-08, 6.47763e-08, 6.543871e-08, 6.50826e-08, 6.546102e-08, 
    6.53923e-08, 6.550608e-08, 6.560798e-08, 6.573618e-08, 6.597273e-08, 
    6.591795e-08, 6.611577e-08, 6.40951e-08, 6.42163e-08, 6.420562e-08, 
    6.433245e-08, 6.442625e-08, 6.462955e-08, 6.49556e-08, 6.483299e-08, 
    6.505808e-08, 6.510327e-08, 6.476129e-08, 6.497127e-08, 6.42974e-08, 
    6.440629e-08, 6.434146e-08, 6.410467e-08, 6.486125e-08, 6.447298e-08, 
    6.518994e-08, 6.49796e-08, 6.559345e-08, 6.528818e-08, 6.58878e-08, 
    6.614415e-08, 6.638538e-08, 6.666732e-08, 6.428244e-08, 6.420009e-08, 
    6.434753e-08, 6.455154e-08, 6.47408e-08, 6.499243e-08, 6.501818e-08, 
    6.506531e-08, 6.518741e-08, 6.529008e-08, 6.508023e-08, 6.531582e-08, 
    6.443155e-08, 6.489495e-08, 6.416896e-08, 6.438758e-08, 6.453951e-08, 
    6.447286e-08, 6.481897e-08, 6.490055e-08, 6.523204e-08, 6.506068e-08, 
    6.608088e-08, 6.562952e-08, 6.688197e-08, 6.653197e-08, 6.417132e-08, 
    6.428215e-08, 6.466789e-08, 6.448436e-08, 6.500922e-08, 6.513842e-08, 
    6.524344e-08, 6.53777e-08, 6.539219e-08, 6.547174e-08, 6.534139e-08, 
    6.546659e-08, 6.499297e-08, 6.520462e-08, 6.46238e-08, 6.476517e-08, 
    6.470013e-08, 6.46288e-08, 6.484896e-08, 6.508353e-08, 6.508854e-08, 
    6.516375e-08, 6.537572e-08, 6.501136e-08, 6.613915e-08, 6.544267e-08, 
    6.440301e-08, 6.461651e-08, 6.464699e-08, 6.456429e-08, 6.512547e-08, 
    6.492213e-08, 6.54698e-08, 6.532179e-08, 6.55643e-08, 6.544379e-08, 
    6.542606e-08, 6.527128e-08, 6.517492e-08, 6.493146e-08, 6.473337e-08, 
    6.457628e-08, 6.461281e-08, 6.478536e-08, 6.509788e-08, 6.539351e-08, 
    6.532875e-08, 6.554587e-08, 6.497117e-08, 6.521216e-08, 6.511902e-08, 
    6.536187e-08, 6.482973e-08, 6.52829e-08, 6.471389e-08, 6.476378e-08, 
    6.49181e-08, 6.522851e-08, 6.529717e-08, 6.53705e-08, 6.532525e-08, 
    6.510581e-08, 6.506986e-08, 6.491435e-08, 6.487141e-08, 6.475292e-08, 
    6.465483e-08, 6.474446e-08, 6.483858e-08, 6.51059e-08, 6.53468e-08, 
    6.560944e-08, 6.567371e-08, 6.59806e-08, 6.573079e-08, 6.614304e-08, 
    6.579257e-08, 6.639924e-08, 6.530915e-08, 6.578225e-08, 6.492512e-08, 
    6.501746e-08, 6.518448e-08, 6.556754e-08, 6.536073e-08, 6.560259e-08, 
    6.506844e-08, 6.479132e-08, 6.471961e-08, 6.458583e-08, 6.472267e-08, 
    6.471154e-08, 6.484247e-08, 6.48004e-08, 6.511478e-08, 6.494591e-08, 
    6.542562e-08, 6.560068e-08, 6.609504e-08, 6.63981e-08, 6.670659e-08, 
    6.684278e-08, 6.688423e-08, 6.690156e-08 ;

 HR_vr =
  2.666893e-07, 2.673978e-07, 2.672601e-07, 2.678311e-07, 2.675144e-07, 
    2.678882e-07, 2.66833e-07, 2.674259e-07, 2.670475e-07, 2.667531e-07, 
    2.689377e-07, 2.678565e-07, 2.700584e-07, 2.693704e-07, 2.710969e-07, 
    2.699514e-07, 2.713276e-07, 2.710638e-07, 2.718573e-07, 2.716301e-07, 
    2.726438e-07, 2.719621e-07, 2.731686e-07, 2.724811e-07, 2.725887e-07, 
    2.719396e-07, 2.680742e-07, 2.688032e-07, 2.68031e-07, 2.68135e-07, 
    2.680883e-07, 2.675209e-07, 2.672349e-07, 2.666351e-07, 2.66744e-07, 
    2.671845e-07, 2.681818e-07, 2.678434e-07, 2.686957e-07, 2.686765e-07, 
    2.696241e-07, 2.69197e-07, 2.707872e-07, 2.703357e-07, 2.716396e-07, 
    2.713119e-07, 2.716242e-07, 2.715295e-07, 2.716254e-07, 2.711448e-07, 
    2.713508e-07, 2.709277e-07, 2.69277e-07, 2.697627e-07, 2.683131e-07, 
    2.674398e-07, 2.66859e-07, 2.664466e-07, 2.665049e-07, 2.666161e-07, 
    2.671871e-07, 2.677234e-07, 2.681318e-07, 2.684048e-07, 2.686737e-07, 
    2.694871e-07, 2.69917e-07, 2.708785e-07, 2.707051e-07, 2.709989e-07, 
    2.712793e-07, 2.7175e-07, 2.716725e-07, 2.718798e-07, 2.709911e-07, 
    2.715819e-07, 2.706063e-07, 2.708733e-07, 2.68747e-07, 2.679347e-07, 
    2.675892e-07, 2.672866e-07, 2.665497e-07, 2.670587e-07, 2.668581e-07, 
    2.673351e-07, 2.676381e-07, 2.674883e-07, 2.684123e-07, 2.680532e-07, 
    2.699425e-07, 2.691295e-07, 2.712466e-07, 2.707407e-07, 2.713678e-07, 
    2.710479e-07, 2.71596e-07, 2.711027e-07, 2.719569e-07, 2.721428e-07, 
    2.720157e-07, 2.725034e-07, 2.710754e-07, 2.716242e-07, 2.674841e-07, 
    2.675085e-07, 2.676223e-07, 2.671219e-07, 2.670912e-07, 2.666321e-07, 
    2.670406e-07, 2.672145e-07, 2.676556e-07, 2.679164e-07, 2.681643e-07, 
    2.687088e-07, 2.693163e-07, 2.701648e-07, 2.707735e-07, 2.711812e-07, 
    2.709312e-07, 2.711519e-07, 2.709052e-07, 2.707895e-07, 2.720731e-07, 
    2.713527e-07, 2.724333e-07, 2.723735e-07, 2.718847e-07, 2.723802e-07, 
    2.675257e-07, 2.67385e-07, 2.668966e-07, 2.672789e-07, 2.665821e-07, 
    2.669723e-07, 2.671965e-07, 2.680608e-07, 2.682505e-07, 2.684264e-07, 
    2.687736e-07, 2.692189e-07, 2.699992e-07, 2.706773e-07, 2.712956e-07, 
    2.712503e-07, 2.712663e-07, 2.714044e-07, 2.710623e-07, 2.714605e-07, 
    2.715273e-07, 2.713526e-07, 2.723655e-07, 2.720763e-07, 2.723722e-07, 
    2.72184e-07, 2.674307e-07, 2.676674e-07, 2.675395e-07, 2.677799e-07, 
    2.676106e-07, 2.683632e-07, 2.685886e-07, 2.696424e-07, 2.692101e-07, 
    2.698979e-07, 2.6928e-07, 2.693895e-07, 2.699204e-07, 2.693134e-07, 
    2.7064e-07, 2.69741e-07, 2.714097e-07, 2.705133e-07, 2.714659e-07, 
    2.712929e-07, 2.715792e-07, 2.718354e-07, 2.721576e-07, 2.727516e-07, 
    2.726141e-07, 2.731105e-07, 2.680199e-07, 2.683265e-07, 2.682995e-07, 
    2.686201e-07, 2.688572e-07, 2.693706e-07, 2.701931e-07, 2.698839e-07, 
    2.704514e-07, 2.705653e-07, 2.697031e-07, 2.702326e-07, 2.685316e-07, 
    2.688068e-07, 2.686429e-07, 2.680441e-07, 2.699553e-07, 2.689752e-07, 
    2.707835e-07, 2.702537e-07, 2.717989e-07, 2.710309e-07, 2.725384e-07, 
    2.731817e-07, 2.737864e-07, 2.744923e-07, 2.684937e-07, 2.682854e-07, 
    2.686582e-07, 2.691737e-07, 2.696514e-07, 2.70286e-07, 2.703509e-07, 
    2.704697e-07, 2.707772e-07, 2.710357e-07, 2.705073e-07, 2.711005e-07, 
    2.688706e-07, 2.700402e-07, 2.682067e-07, 2.687595e-07, 2.691433e-07, 
    2.689749e-07, 2.698486e-07, 2.700543e-07, 2.708896e-07, 2.70458e-07, 
    2.730231e-07, 2.718896e-07, 2.750291e-07, 2.741535e-07, 2.682127e-07, 
    2.68493e-07, 2.694674e-07, 2.69004e-07, 2.703283e-07, 2.706539e-07, 
    2.709183e-07, 2.712562e-07, 2.712927e-07, 2.714928e-07, 2.711648e-07, 
    2.714798e-07, 2.702873e-07, 2.708205e-07, 2.693561e-07, 2.697129e-07, 
    2.695488e-07, 2.693687e-07, 2.699242e-07, 2.705156e-07, 2.705282e-07, 
    2.707176e-07, 2.712513e-07, 2.703337e-07, 2.731693e-07, 2.714198e-07, 
    2.687984e-07, 2.693377e-07, 2.694146e-07, 2.692058e-07, 2.706212e-07, 
    2.701088e-07, 2.714879e-07, 2.711155e-07, 2.717256e-07, 2.714225e-07, 
    2.713779e-07, 2.709884e-07, 2.707457e-07, 2.701323e-07, 2.696326e-07, 
    2.692361e-07, 2.693283e-07, 2.697638e-07, 2.705517e-07, 2.71296e-07, 
    2.71133e-07, 2.716793e-07, 2.702324e-07, 2.708395e-07, 2.70605e-07, 
    2.712164e-07, 2.698757e-07, 2.710177e-07, 2.695835e-07, 2.697094e-07, 
    2.700986e-07, 2.708807e-07, 2.710535e-07, 2.712381e-07, 2.711242e-07, 
    2.705717e-07, 2.704811e-07, 2.700891e-07, 2.699809e-07, 2.69682e-07, 
    2.694344e-07, 2.696606e-07, 2.698981e-07, 2.705719e-07, 2.711785e-07, 
    2.718391e-07, 2.720006e-07, 2.727714e-07, 2.721441e-07, 2.73179e-07, 
    2.722994e-07, 2.738212e-07, 2.710838e-07, 2.722734e-07, 2.701163e-07, 
    2.703491e-07, 2.707698e-07, 2.717338e-07, 2.712135e-07, 2.718219e-07, 
    2.704776e-07, 2.697789e-07, 2.695979e-07, 2.692602e-07, 2.696056e-07, 
    2.695776e-07, 2.699079e-07, 2.698017e-07, 2.705943e-07, 2.701687e-07, 
    2.713768e-07, 2.718171e-07, 2.730585e-07, 2.738183e-07, 2.745905e-07, 
    2.749311e-07, 2.750347e-07, 2.75078e-07,
  2.414476e-07, 2.42358e-07, 2.421811e-07, 2.429149e-07, 2.425079e-07, 
    2.429883e-07, 2.416322e-07, 2.423941e-07, 2.419078e-07, 2.415296e-07, 
    2.443372e-07, 2.429476e-07, 2.457786e-07, 2.44894e-07, 2.471145e-07, 
    2.45641e-07, 2.474114e-07, 2.470721e-07, 2.480929e-07, 2.478006e-07, 
    2.491049e-07, 2.482278e-07, 2.497804e-07, 2.488956e-07, 2.49034e-07, 
    2.481989e-07, 2.432275e-07, 2.441643e-07, 2.431719e-07, 2.433056e-07, 
    2.432456e-07, 2.425163e-07, 2.421486e-07, 2.41378e-07, 2.415179e-07, 
    2.420839e-07, 2.433657e-07, 2.429308e-07, 2.440265e-07, 2.440018e-07, 
    2.452201e-07, 2.44671e-07, 2.467162e-07, 2.461354e-07, 2.478128e-07, 
    2.473912e-07, 2.47793e-07, 2.476712e-07, 2.477946e-07, 2.471762e-07, 
    2.474412e-07, 2.468969e-07, 2.447738e-07, 2.453983e-07, 2.435345e-07, 
    2.424119e-07, 2.416656e-07, 2.411357e-07, 2.412106e-07, 2.413535e-07, 
    2.420872e-07, 2.427765e-07, 2.433015e-07, 2.436525e-07, 2.439982e-07, 
    2.450438e-07, 2.455968e-07, 2.468336e-07, 2.466105e-07, 2.469884e-07, 
    2.473493e-07, 2.479548e-07, 2.478552e-07, 2.481218e-07, 2.469785e-07, 
    2.477385e-07, 2.464835e-07, 2.468269e-07, 2.440921e-07, 2.430481e-07, 
    2.42604e-07, 2.422151e-07, 2.412683e-07, 2.419222e-07, 2.416645e-07, 
    2.422776e-07, 2.426669e-07, 2.424744e-07, 2.436621e-07, 2.432005e-07, 
    2.456295e-07, 2.445841e-07, 2.473072e-07, 2.466563e-07, 2.474632e-07, 
    2.470516e-07, 2.477567e-07, 2.471221e-07, 2.482211e-07, 2.484602e-07, 
    2.482968e-07, 2.489243e-07, 2.470869e-07, 2.47793e-07, 2.42469e-07, 
    2.425004e-07, 2.426467e-07, 2.420034e-07, 2.41964e-07, 2.413741e-07, 
    2.41899e-07, 2.421225e-07, 2.426895e-07, 2.430247e-07, 2.433432e-07, 
    2.440432e-07, 2.448243e-07, 2.459155e-07, 2.466985e-07, 2.472231e-07, 
    2.469015e-07, 2.471854e-07, 2.46868e-07, 2.467192e-07, 2.483706e-07, 
    2.474437e-07, 2.488341e-07, 2.487572e-07, 2.481282e-07, 2.487659e-07, 
    2.425224e-07, 2.423417e-07, 2.417139e-07, 2.422053e-07, 2.413099e-07, 
    2.418112e-07, 2.420992e-07, 2.432102e-07, 2.434541e-07, 2.436802e-07, 
    2.441266e-07, 2.446991e-07, 2.457026e-07, 2.465748e-07, 2.473703e-07, 
    2.47312e-07, 2.473325e-07, 2.475101e-07, 2.470701e-07, 2.475824e-07, 
    2.476683e-07, 2.474436e-07, 2.487469e-07, 2.483748e-07, 2.487556e-07, 
    2.485133e-07, 2.424005e-07, 2.427045e-07, 2.425402e-07, 2.428492e-07, 
    2.426315e-07, 2.435989e-07, 2.438887e-07, 2.452436e-07, 2.446878e-07, 
    2.455723e-07, 2.447777e-07, 2.449186e-07, 2.456011e-07, 2.448207e-07, 
    2.465267e-07, 2.453704e-07, 2.475171e-07, 2.463636e-07, 2.475893e-07, 
    2.473668e-07, 2.477351e-07, 2.480648e-07, 2.484794e-07, 2.492438e-07, 
    2.490668e-07, 2.497057e-07, 2.431577e-07, 2.435517e-07, 2.435171e-07, 
    2.439293e-07, 2.44234e-07, 2.448942e-07, 2.45952e-07, 2.455544e-07, 
    2.462843e-07, 2.464307e-07, 2.453218e-07, 2.460028e-07, 2.438154e-07, 
    2.441691e-07, 2.439585e-07, 2.431888e-07, 2.45646e-07, 2.443857e-07, 
    2.467115e-07, 2.460298e-07, 2.480178e-07, 2.470296e-07, 2.489694e-07, 
    2.497972e-07, 2.505757e-07, 2.514845e-07, 2.437667e-07, 2.434991e-07, 
    2.439783e-07, 2.446409e-07, 2.452553e-07, 2.460714e-07, 2.461549e-07, 
    2.463077e-07, 2.467033e-07, 2.470359e-07, 2.46356e-07, 2.471192e-07, 
    2.442511e-07, 2.457553e-07, 2.433978e-07, 2.441083e-07, 2.446019e-07, 
    2.443854e-07, 2.455089e-07, 2.457735e-07, 2.468478e-07, 2.462927e-07, 
    2.49593e-07, 2.481344e-07, 2.521758e-07, 2.510483e-07, 2.434055e-07, 
    2.437658e-07, 2.450187e-07, 2.444228e-07, 2.461259e-07, 2.465446e-07, 
    2.468848e-07, 2.473195e-07, 2.473665e-07, 2.476239e-07, 2.47202e-07, 
    2.476073e-07, 2.460732e-07, 2.46759e-07, 2.448756e-07, 2.453343e-07, 
    2.451233e-07, 2.448918e-07, 2.456062e-07, 2.463667e-07, 2.463829e-07, 
    2.466266e-07, 2.473129e-07, 2.461328e-07, 2.49781e-07, 2.475297e-07, 
    2.441585e-07, 2.448518e-07, 2.449508e-07, 2.446824e-07, 2.465026e-07, 
    2.458435e-07, 2.476177e-07, 2.471385e-07, 2.479235e-07, 2.475335e-07, 
    2.474761e-07, 2.46975e-07, 2.466628e-07, 2.458737e-07, 2.452311e-07, 
    2.447213e-07, 2.448399e-07, 2.453999e-07, 2.464132e-07, 2.473707e-07, 
    2.47161e-07, 2.478639e-07, 2.460025e-07, 2.467834e-07, 2.464817e-07, 
    2.472683e-07, 2.455438e-07, 2.470124e-07, 2.45168e-07, 2.453299e-07, 
    2.458304e-07, 2.468364e-07, 2.470588e-07, 2.472962e-07, 2.471498e-07, 
    2.464389e-07, 2.463224e-07, 2.458183e-07, 2.45679e-07, 2.452946e-07, 
    2.449763e-07, 2.452672e-07, 2.455725e-07, 2.464392e-07, 2.472195e-07, 
    2.480695e-07, 2.482774e-07, 2.492691e-07, 2.484618e-07, 2.497935e-07, 
    2.486614e-07, 2.506202e-07, 2.470975e-07, 2.486281e-07, 2.458532e-07, 
    2.461526e-07, 2.466938e-07, 2.479339e-07, 2.472646e-07, 2.480473e-07, 
    2.463178e-07, 2.454192e-07, 2.451866e-07, 2.447523e-07, 2.451965e-07, 
    2.451604e-07, 2.455852e-07, 2.454487e-07, 2.46468e-07, 2.459206e-07, 
    2.474747e-07, 2.480411e-07, 2.496388e-07, 2.506167e-07, 2.516111e-07, 
    2.520497e-07, 2.521831e-07, 2.522389e-07,
  2.259466e-07, 2.269439e-07, 2.267501e-07, 2.275541e-07, 2.271082e-07, 
    2.276345e-07, 2.261489e-07, 2.269835e-07, 2.264508e-07, 2.260365e-07, 
    2.29113e-07, 2.275899e-07, 2.306936e-07, 2.297234e-07, 2.321593e-07, 
    2.305427e-07, 2.324851e-07, 2.321127e-07, 2.332332e-07, 2.329123e-07, 
    2.343444e-07, 2.333813e-07, 2.350862e-07, 2.341145e-07, 2.342665e-07, 
    2.333495e-07, 2.278966e-07, 2.289235e-07, 2.278357e-07, 2.279822e-07, 
    2.279165e-07, 2.271174e-07, 2.267144e-07, 2.258704e-07, 2.260237e-07, 
    2.266436e-07, 2.280481e-07, 2.275715e-07, 2.287724e-07, 2.287453e-07, 
    2.300811e-07, 2.29479e-07, 2.317223e-07, 2.310851e-07, 2.329257e-07, 
    2.32463e-07, 2.32904e-07, 2.327703e-07, 2.329057e-07, 2.322271e-07, 
    2.325179e-07, 2.319206e-07, 2.295917e-07, 2.302765e-07, 2.282331e-07, 
    2.27003e-07, 2.261855e-07, 2.256051e-07, 2.256871e-07, 2.258436e-07, 
    2.266472e-07, 2.274025e-07, 2.279778e-07, 2.283624e-07, 2.287414e-07, 
    2.298877e-07, 2.304942e-07, 2.318511e-07, 2.316063e-07, 2.320209e-07, 
    2.32417e-07, 2.330816e-07, 2.329722e-07, 2.33265e-07, 2.3201e-07, 
    2.328442e-07, 2.314669e-07, 2.318437e-07, 2.288443e-07, 2.277001e-07, 
    2.272134e-07, 2.267873e-07, 2.257502e-07, 2.264665e-07, 2.261842e-07, 
    2.268558e-07, 2.272824e-07, 2.270714e-07, 2.28373e-07, 2.278671e-07, 
    2.305301e-07, 2.293837e-07, 2.323708e-07, 2.316566e-07, 2.325419e-07, 
    2.320902e-07, 2.328641e-07, 2.321676e-07, 2.333739e-07, 2.336364e-07, 
    2.33457e-07, 2.34146e-07, 2.32129e-07, 2.329039e-07, 2.270655e-07, 
    2.270999e-07, 2.272602e-07, 2.265554e-07, 2.265123e-07, 2.258662e-07, 
    2.264411e-07, 2.266859e-07, 2.273071e-07, 2.276744e-07, 2.280235e-07, 
    2.287907e-07, 2.296471e-07, 2.308438e-07, 2.317029e-07, 2.322785e-07, 
    2.319255e-07, 2.322371e-07, 2.318888e-07, 2.317255e-07, 2.33538e-07, 
    2.325206e-07, 2.340469e-07, 2.339625e-07, 2.332719e-07, 2.33972e-07, 
    2.271241e-07, 2.269261e-07, 2.262383e-07, 2.267766e-07, 2.257958e-07, 
    2.263449e-07, 2.266604e-07, 2.278776e-07, 2.28145e-07, 2.283928e-07, 
    2.288821e-07, 2.295098e-07, 2.306103e-07, 2.315671e-07, 2.3244e-07, 
    2.323761e-07, 2.323986e-07, 2.325935e-07, 2.321106e-07, 2.326728e-07, 
    2.327671e-07, 2.325205e-07, 2.339512e-07, 2.335426e-07, 2.339607e-07, 
    2.336947e-07, 2.269904e-07, 2.273236e-07, 2.271436e-07, 2.274821e-07, 
    2.272436e-07, 2.283036e-07, 2.286213e-07, 2.301069e-07, 2.294974e-07, 
    2.304673e-07, 2.29596e-07, 2.297504e-07, 2.304989e-07, 2.296431e-07, 
    2.315143e-07, 2.302459e-07, 2.326011e-07, 2.313354e-07, 2.326804e-07, 
    2.324362e-07, 2.328404e-07, 2.332023e-07, 2.336575e-07, 2.344969e-07, 
    2.343025e-07, 2.350042e-07, 2.278201e-07, 2.28252e-07, 2.28214e-07, 
    2.286658e-07, 2.289999e-07, 2.297237e-07, 2.308838e-07, 2.304477e-07, 
    2.312483e-07, 2.31409e-07, 2.301926e-07, 2.309395e-07, 2.28541e-07, 
    2.289287e-07, 2.286979e-07, 2.278542e-07, 2.305482e-07, 2.291662e-07, 
    2.317171e-07, 2.309692e-07, 2.331507e-07, 2.320662e-07, 2.341955e-07, 
    2.351048e-07, 2.3596e-07, 2.369587e-07, 2.284877e-07, 2.281943e-07, 
    2.287195e-07, 2.294459e-07, 2.301197e-07, 2.310148e-07, 2.311064e-07, 
    2.31274e-07, 2.317081e-07, 2.32073e-07, 2.31327e-07, 2.321645e-07, 
    2.290186e-07, 2.306681e-07, 2.280833e-07, 2.288621e-07, 2.294032e-07, 
    2.291659e-07, 2.303978e-07, 2.30688e-07, 2.318667e-07, 2.312575e-07, 
    2.348804e-07, 2.332787e-07, 2.377187e-07, 2.364794e-07, 2.280917e-07, 
    2.284866e-07, 2.298602e-07, 2.292068e-07, 2.310746e-07, 2.315339e-07, 
    2.319073e-07, 2.323843e-07, 2.324358e-07, 2.327184e-07, 2.322553e-07, 
    2.327001e-07, 2.310167e-07, 2.317692e-07, 2.297033e-07, 2.302064e-07, 
    2.29975e-07, 2.297211e-07, 2.305045e-07, 2.313387e-07, 2.313566e-07, 
    2.316239e-07, 2.32377e-07, 2.310821e-07, 2.350869e-07, 2.32615e-07, 
    2.289171e-07, 2.296772e-07, 2.297858e-07, 2.294914e-07, 2.314879e-07, 
    2.307648e-07, 2.327115e-07, 2.321857e-07, 2.330472e-07, 2.326191e-07, 
    2.325562e-07, 2.320062e-07, 2.316637e-07, 2.30798e-07, 2.300932e-07, 
    2.295341e-07, 2.296641e-07, 2.302782e-07, 2.313897e-07, 2.324405e-07, 
    2.322104e-07, 2.329817e-07, 2.309392e-07, 2.31796e-07, 2.314649e-07, 
    2.323281e-07, 2.304361e-07, 2.320473e-07, 2.300239e-07, 2.302015e-07, 
    2.307505e-07, 2.318541e-07, 2.320982e-07, 2.323587e-07, 2.32198e-07, 
    2.31418e-07, 2.312901e-07, 2.307371e-07, 2.305844e-07, 2.301628e-07, 
    2.298137e-07, 2.301327e-07, 2.304676e-07, 2.314183e-07, 2.322745e-07, 
    2.332074e-07, 2.334357e-07, 2.345247e-07, 2.336382e-07, 2.351007e-07, 
    2.338573e-07, 2.360089e-07, 2.321407e-07, 2.338208e-07, 2.307754e-07, 
    2.311039e-07, 2.316976e-07, 2.330586e-07, 2.323241e-07, 2.331831e-07, 
    2.312851e-07, 2.302994e-07, 2.300443e-07, 2.295681e-07, 2.300552e-07, 
    2.300155e-07, 2.304815e-07, 2.303318e-07, 2.314499e-07, 2.308494e-07, 
    2.325546e-07, 2.331763e-07, 2.349307e-07, 2.360051e-07, 2.370979e-07, 
    2.3758e-07, 2.377267e-07, 2.377881e-07,
  2.166375e-07, 2.17664e-07, 2.174645e-07, 2.182923e-07, 2.178331e-07, 
    2.183752e-07, 2.168456e-07, 2.177048e-07, 2.171563e-07, 2.167299e-07, 
    2.198986e-07, 2.183292e-07, 2.215282e-07, 2.205277e-07, 2.230406e-07, 
    2.213725e-07, 2.233769e-07, 2.229925e-07, 2.241493e-07, 2.238179e-07, 
    2.252974e-07, 2.243023e-07, 2.260641e-07, 2.250597e-07, 2.252169e-07, 
    2.242694e-07, 2.186451e-07, 2.197032e-07, 2.185824e-07, 2.187333e-07, 
    2.186656e-07, 2.178426e-07, 2.174278e-07, 2.16559e-07, 2.167168e-07, 
    2.173549e-07, 2.188011e-07, 2.183102e-07, 2.195474e-07, 2.195194e-07, 
    2.208964e-07, 2.202756e-07, 2.225894e-07, 2.219319e-07, 2.238317e-07, 
    2.23354e-07, 2.238093e-07, 2.236713e-07, 2.238111e-07, 2.231105e-07, 
    2.234107e-07, 2.227941e-07, 2.203919e-07, 2.21098e-07, 2.189918e-07, 
    2.177249e-07, 2.168833e-07, 2.16286e-07, 2.163705e-07, 2.165314e-07, 
    2.173586e-07, 2.181362e-07, 2.187287e-07, 2.19125e-07, 2.195154e-07, 
    2.206971e-07, 2.213225e-07, 2.227224e-07, 2.224698e-07, 2.228977e-07, 
    2.233065e-07, 2.239928e-07, 2.238798e-07, 2.241821e-07, 2.228864e-07, 
    2.237476e-07, 2.223259e-07, 2.227148e-07, 2.196216e-07, 2.184427e-07, 
    2.179415e-07, 2.175028e-07, 2.164354e-07, 2.171726e-07, 2.16882e-07, 
    2.175733e-07, 2.180125e-07, 2.177953e-07, 2.191358e-07, 2.186147e-07, 
    2.213595e-07, 2.201774e-07, 2.232588e-07, 2.225216e-07, 2.234355e-07, 
    2.229692e-07, 2.237682e-07, 2.230491e-07, 2.242947e-07, 2.245658e-07, 
    2.243805e-07, 2.250923e-07, 2.230092e-07, 2.238093e-07, 2.177892e-07, 
    2.178246e-07, 2.179897e-07, 2.172641e-07, 2.172197e-07, 2.165547e-07, 
    2.171464e-07, 2.173984e-07, 2.18038e-07, 2.184162e-07, 2.187758e-07, 
    2.195663e-07, 2.20449e-07, 2.21683e-07, 2.225694e-07, 2.231635e-07, 
    2.227992e-07, 2.231208e-07, 2.227613e-07, 2.225928e-07, 2.244642e-07, 
    2.234135e-07, 2.249899e-07, 2.249027e-07, 2.241893e-07, 2.249126e-07, 
    2.178495e-07, 2.176456e-07, 2.169377e-07, 2.174917e-07, 2.164823e-07, 
    2.170473e-07, 2.173722e-07, 2.186256e-07, 2.189009e-07, 2.191562e-07, 
    2.196604e-07, 2.203074e-07, 2.214421e-07, 2.224293e-07, 2.233303e-07, 
    2.232643e-07, 2.232875e-07, 2.234888e-07, 2.229902e-07, 2.235706e-07, 
    2.23668e-07, 2.234133e-07, 2.248911e-07, 2.244689e-07, 2.249009e-07, 
    2.24626e-07, 2.177119e-07, 2.180549e-07, 2.178696e-07, 2.182181e-07, 
    2.179726e-07, 2.190644e-07, 2.193917e-07, 2.209231e-07, 2.202946e-07, 
    2.212947e-07, 2.203962e-07, 2.205554e-07, 2.213274e-07, 2.204448e-07, 
    2.223749e-07, 2.210664e-07, 2.234966e-07, 2.221903e-07, 2.235784e-07, 
    2.233264e-07, 2.237437e-07, 2.241174e-07, 2.245876e-07, 2.254549e-07, 
    2.252541e-07, 2.259793e-07, 2.185663e-07, 2.190112e-07, 2.18972e-07, 
    2.194376e-07, 2.197818e-07, 2.205279e-07, 2.217243e-07, 2.212744e-07, 
    2.221003e-07, 2.222661e-07, 2.210114e-07, 2.217818e-07, 2.193089e-07, 
    2.197085e-07, 2.194706e-07, 2.186014e-07, 2.213781e-07, 2.199533e-07, 
    2.22584e-07, 2.218124e-07, 2.240641e-07, 2.229444e-07, 2.251435e-07, 
    2.260833e-07, 2.269677e-07, 2.28001e-07, 2.19254e-07, 2.189517e-07, 
    2.194929e-07, 2.202416e-07, 2.209362e-07, 2.218595e-07, 2.219539e-07, 
    2.221269e-07, 2.225748e-07, 2.229514e-07, 2.221816e-07, 2.230458e-07, 
    2.198012e-07, 2.215018e-07, 2.188374e-07, 2.196399e-07, 2.201975e-07, 
    2.199529e-07, 2.21223e-07, 2.215224e-07, 2.227385e-07, 2.221099e-07, 
    2.258514e-07, 2.241964e-07, 2.287875e-07, 2.275049e-07, 2.188461e-07, 
    2.192529e-07, 2.206686e-07, 2.199951e-07, 2.219211e-07, 2.223951e-07, 
    2.227803e-07, 2.232728e-07, 2.23326e-07, 2.236177e-07, 2.231396e-07, 
    2.235988e-07, 2.218614e-07, 2.226379e-07, 2.205068e-07, 2.210256e-07, 
    2.20787e-07, 2.205252e-07, 2.213331e-07, 2.221937e-07, 2.222121e-07, 
    2.22488e-07, 2.232655e-07, 2.219289e-07, 2.26065e-07, 2.235111e-07, 
    2.196965e-07, 2.2048e-07, 2.205919e-07, 2.202884e-07, 2.223476e-07, 
    2.216016e-07, 2.236106e-07, 2.230677e-07, 2.239572e-07, 2.235152e-07, 
    2.234502e-07, 2.228824e-07, 2.22529e-07, 2.216358e-07, 2.209089e-07, 
    2.203325e-07, 2.204665e-07, 2.210997e-07, 2.222463e-07, 2.233308e-07, 
    2.230933e-07, 2.238896e-07, 2.217815e-07, 2.226656e-07, 2.223239e-07, 
    2.232148e-07, 2.212625e-07, 2.229251e-07, 2.208375e-07, 2.210205e-07, 
    2.215867e-07, 2.227255e-07, 2.229774e-07, 2.232464e-07, 2.230804e-07, 
    2.222754e-07, 2.221435e-07, 2.21573e-07, 2.214154e-07, 2.209807e-07, 
    2.206207e-07, 2.209496e-07, 2.21295e-07, 2.222757e-07, 2.231594e-07, 
    2.241227e-07, 2.243585e-07, 2.254837e-07, 2.245678e-07, 2.260792e-07, 
    2.247942e-07, 2.270184e-07, 2.230214e-07, 2.247564e-07, 2.216125e-07, 
    2.219513e-07, 2.22564e-07, 2.239691e-07, 2.232106e-07, 2.240976e-07, 
    2.221383e-07, 2.211216e-07, 2.208584e-07, 2.203675e-07, 2.208697e-07, 
    2.208288e-07, 2.213093e-07, 2.211549e-07, 2.223083e-07, 2.216888e-07, 
    2.234486e-07, 2.240906e-07, 2.259033e-07, 2.270143e-07, 2.281449e-07, 
    2.286439e-07, 2.287958e-07, 2.288593e-07,
  2.081375e-07, 2.091063e-07, 2.089179e-07, 2.096997e-07, 2.092659e-07, 
    2.097779e-07, 2.083338e-07, 2.091448e-07, 2.08627e-07, 2.082246e-07, 
    2.112182e-07, 2.097346e-07, 2.127607e-07, 2.118133e-07, 2.141943e-07, 
    2.126132e-07, 2.145133e-07, 2.141486e-07, 2.152464e-07, 2.149318e-07, 
    2.163371e-07, 2.153916e-07, 2.17066e-07, 2.161112e-07, 2.162605e-07, 
    2.153604e-07, 2.100329e-07, 2.110334e-07, 2.099737e-07, 2.101163e-07, 
    2.100523e-07, 2.092749e-07, 2.088833e-07, 2.080634e-07, 2.082122e-07, 
    2.088144e-07, 2.101804e-07, 2.097165e-07, 2.108858e-07, 2.108594e-07, 
    2.121623e-07, 2.115747e-07, 2.137664e-07, 2.131431e-07, 2.149449e-07, 
    2.144916e-07, 2.149236e-07, 2.147926e-07, 2.149253e-07, 2.142605e-07, 
    2.145453e-07, 2.139604e-07, 2.116848e-07, 2.123532e-07, 2.103606e-07, 
    2.091639e-07, 2.083694e-07, 2.078059e-07, 2.078856e-07, 2.080374e-07, 
    2.088179e-07, 2.095521e-07, 2.101119e-07, 2.104865e-07, 2.108556e-07, 
    2.119738e-07, 2.125658e-07, 2.138925e-07, 2.136529e-07, 2.140587e-07, 
    2.144465e-07, 2.150978e-07, 2.149905e-07, 2.152776e-07, 2.14048e-07, 
    2.148651e-07, 2.135165e-07, 2.138852e-07, 2.109562e-07, 2.098417e-07, 
    2.093684e-07, 2.089541e-07, 2.079468e-07, 2.086424e-07, 2.083681e-07, 
    2.090206e-07, 2.094353e-07, 2.092302e-07, 2.104967e-07, 2.100042e-07, 
    2.126009e-07, 2.114818e-07, 2.144012e-07, 2.137021e-07, 2.145689e-07, 
    2.141265e-07, 2.148846e-07, 2.142023e-07, 2.153844e-07, 2.156419e-07, 
    2.154659e-07, 2.161421e-07, 2.141645e-07, 2.149236e-07, 2.092244e-07, 
    2.092579e-07, 2.094137e-07, 2.087287e-07, 2.086868e-07, 2.080593e-07, 
    2.086177e-07, 2.088555e-07, 2.094593e-07, 2.098167e-07, 2.101564e-07, 
    2.109037e-07, 2.117388e-07, 2.129073e-07, 2.137474e-07, 2.143108e-07, 
    2.139653e-07, 2.142703e-07, 2.139293e-07, 2.137695e-07, 2.155455e-07, 
    2.14548e-07, 2.160448e-07, 2.15962e-07, 2.152844e-07, 2.159713e-07, 
    2.092814e-07, 2.090889e-07, 2.084207e-07, 2.089436e-07, 2.07991e-07, 
    2.085242e-07, 2.088308e-07, 2.100145e-07, 2.102747e-07, 2.10516e-07, 
    2.109927e-07, 2.116048e-07, 2.126792e-07, 2.136146e-07, 2.14469e-07, 
    2.144064e-07, 2.144284e-07, 2.146194e-07, 2.141465e-07, 2.146971e-07, 
    2.147895e-07, 2.145478e-07, 2.159509e-07, 2.155499e-07, 2.159602e-07, 
    2.156991e-07, 2.091514e-07, 2.094754e-07, 2.093003e-07, 2.096296e-07, 
    2.093976e-07, 2.104293e-07, 2.107387e-07, 2.121876e-07, 2.115927e-07, 
    2.125395e-07, 2.116889e-07, 2.118396e-07, 2.125705e-07, 2.117348e-07, 
    2.13563e-07, 2.123234e-07, 2.146268e-07, 2.133881e-07, 2.147045e-07, 
    2.144653e-07, 2.148613e-07, 2.152161e-07, 2.156626e-07, 2.164868e-07, 
    2.162958e-07, 2.169854e-07, 2.099585e-07, 2.103789e-07, 2.103419e-07, 
    2.10782e-07, 2.111076e-07, 2.118135e-07, 2.129464e-07, 2.125203e-07, 
    2.133027e-07, 2.134598e-07, 2.122712e-07, 2.130009e-07, 2.106604e-07, 
    2.110383e-07, 2.108133e-07, 2.099917e-07, 2.126185e-07, 2.112698e-07, 
    2.137613e-07, 2.130299e-07, 2.151655e-07, 2.141031e-07, 2.161908e-07, 
    2.170844e-07, 2.179257e-07, 2.189099e-07, 2.106084e-07, 2.103227e-07, 
    2.108343e-07, 2.115426e-07, 2.122e-07, 2.130745e-07, 2.13164e-07, 
    2.133279e-07, 2.137525e-07, 2.141096e-07, 2.133798e-07, 2.141992e-07, 
    2.111261e-07, 2.127356e-07, 2.102147e-07, 2.109734e-07, 2.115008e-07, 
    2.112694e-07, 2.124716e-07, 2.127551e-07, 2.139078e-07, 2.133117e-07, 
    2.168638e-07, 2.152911e-07, 2.196596e-07, 2.184373e-07, 2.102229e-07, 
    2.106074e-07, 2.119467e-07, 2.113093e-07, 2.131329e-07, 2.135821e-07, 
    2.139474e-07, 2.144145e-07, 2.144649e-07, 2.147418e-07, 2.142881e-07, 
    2.147239e-07, 2.130763e-07, 2.138123e-07, 2.117935e-07, 2.122846e-07, 
    2.120587e-07, 2.118109e-07, 2.125758e-07, 2.133913e-07, 2.134086e-07, 
    2.136702e-07, 2.144078e-07, 2.131403e-07, 2.170671e-07, 2.146407e-07, 
    2.110269e-07, 2.117683e-07, 2.118741e-07, 2.115869e-07, 2.135371e-07, 
    2.128301e-07, 2.14735e-07, 2.142199e-07, 2.15064e-07, 2.146445e-07, 
    2.145828e-07, 2.140442e-07, 2.13709e-07, 2.128625e-07, 2.121742e-07, 
    2.116285e-07, 2.117554e-07, 2.123548e-07, 2.134411e-07, 2.144695e-07, 
    2.142442e-07, 2.149998e-07, 2.130006e-07, 2.138386e-07, 2.135147e-07, 
    2.143594e-07, 2.12509e-07, 2.140848e-07, 2.121065e-07, 2.122798e-07, 
    2.128161e-07, 2.138955e-07, 2.141343e-07, 2.143895e-07, 2.14232e-07, 
    2.134687e-07, 2.133437e-07, 2.12803e-07, 2.126538e-07, 2.122421e-07, 
    2.119013e-07, 2.122127e-07, 2.125398e-07, 2.13469e-07, 2.14307e-07, 
    2.152212e-07, 2.15445e-07, 2.165143e-07, 2.156439e-07, 2.170806e-07, 
    2.158592e-07, 2.179742e-07, 2.141761e-07, 2.158231e-07, 2.128405e-07, 
    2.131615e-07, 2.137423e-07, 2.150753e-07, 2.143555e-07, 2.151974e-07, 
    2.133388e-07, 2.123756e-07, 2.121264e-07, 2.116617e-07, 2.12137e-07, 
    2.120983e-07, 2.125533e-07, 2.12407e-07, 2.134999e-07, 2.129127e-07, 
    2.145813e-07, 2.151907e-07, 2.169131e-07, 2.179702e-07, 2.190469e-07, 
    2.195226e-07, 2.196675e-07, 2.19728e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.356978e-08, 6.384934e-08, 6.379499e-08, 6.402048e-08, 6.389539e-08, 
    6.404304e-08, 6.362645e-08, 6.386044e-08, 6.371106e-08, 6.359494e-08, 
    6.445807e-08, 6.403054e-08, 6.490213e-08, 6.462948e-08, 6.531439e-08, 
    6.485971e-08, 6.540607e-08, 6.530126e-08, 6.561668e-08, 6.552632e-08, 
    6.592977e-08, 6.565838e-08, 6.61389e-08, 6.586495e-08, 6.590781e-08, 
    6.564943e-08, 6.411657e-08, 6.440485e-08, 6.409949e-08, 6.41406e-08, 
    6.412215e-08, 6.389798e-08, 6.378502e-08, 6.354841e-08, 6.359136e-08, 
    6.376514e-08, 6.415908e-08, 6.402535e-08, 6.436237e-08, 6.435476e-08, 
    6.472996e-08, 6.456079e-08, 6.51914e-08, 6.501217e-08, 6.553009e-08, 
    6.539984e-08, 6.552398e-08, 6.548633e-08, 6.552447e-08, 6.533344e-08, 
    6.541529e-08, 6.524719e-08, 6.459248e-08, 6.478489e-08, 6.421101e-08, 
    6.386593e-08, 6.363672e-08, 6.347406e-08, 6.349706e-08, 6.35409e-08, 
    6.376616e-08, 6.397794e-08, 6.413933e-08, 6.42473e-08, 6.435366e-08, 
    6.467567e-08, 6.484608e-08, 6.522765e-08, 6.515878e-08, 6.527544e-08, 
    6.538689e-08, 6.557399e-08, 6.55432e-08, 6.562563e-08, 6.527236e-08, 
    6.550714e-08, 6.511956e-08, 6.522556e-08, 6.438261e-08, 6.406143e-08, 
    6.392494e-08, 6.380544e-08, 6.351474e-08, 6.371549e-08, 6.363636e-08, 
    6.382462e-08, 6.394425e-08, 6.388508e-08, 6.425024e-08, 6.410828e-08, 
    6.485618e-08, 6.453404e-08, 6.537388e-08, 6.517291e-08, 6.542206e-08, 
    6.529492e-08, 6.551276e-08, 6.53167e-08, 6.565631e-08, 6.573026e-08, 
    6.567973e-08, 6.587384e-08, 6.530584e-08, 6.552398e-08, 6.388343e-08, 
    6.389308e-08, 6.393803e-08, 6.374042e-08, 6.372833e-08, 6.354723e-08, 
    6.370837e-08, 6.377699e-08, 6.395118e-08, 6.405422e-08, 6.415217e-08, 
    6.436752e-08, 6.460803e-08, 6.494434e-08, 6.518594e-08, 6.53479e-08, 
    6.524859e-08, 6.533626e-08, 6.523825e-08, 6.519231e-08, 6.570255e-08, 
    6.541605e-08, 6.584592e-08, 6.582213e-08, 6.562759e-08, 6.582481e-08, 
    6.389985e-08, 6.384432e-08, 6.365153e-08, 6.38024e-08, 6.352751e-08, 
    6.368138e-08, 6.376987e-08, 6.411125e-08, 6.418625e-08, 6.425581e-08, 
    6.439316e-08, 6.456945e-08, 6.487869e-08, 6.514775e-08, 6.539337e-08, 
    6.537537e-08, 6.538171e-08, 6.543657e-08, 6.530066e-08, 6.545889e-08, 
    6.548544e-08, 6.541601e-08, 6.581894e-08, 6.570383e-08, 6.582162e-08, 
    6.574668e-08, 6.386237e-08, 6.395581e-08, 6.390532e-08, 6.400027e-08, 
    6.393338e-08, 6.42308e-08, 6.431998e-08, 6.473723e-08, 6.456598e-08, 
    6.483852e-08, 6.459366e-08, 6.463705e-08, 6.484741e-08, 6.460689e-08, 
    6.513292e-08, 6.47763e-08, 6.543871e-08, 6.50826e-08, 6.546102e-08, 
    6.53923e-08, 6.550608e-08, 6.560798e-08, 6.573618e-08, 6.597273e-08, 
    6.591795e-08, 6.611577e-08, 6.40951e-08, 6.42163e-08, 6.420562e-08, 
    6.433245e-08, 6.442625e-08, 6.462955e-08, 6.49556e-08, 6.483299e-08, 
    6.505808e-08, 6.510327e-08, 6.476129e-08, 6.497127e-08, 6.42974e-08, 
    6.440629e-08, 6.434146e-08, 6.410467e-08, 6.486125e-08, 6.447298e-08, 
    6.518994e-08, 6.49796e-08, 6.559345e-08, 6.528818e-08, 6.58878e-08, 
    6.614415e-08, 6.638538e-08, 6.666732e-08, 6.428244e-08, 6.420009e-08, 
    6.434753e-08, 6.455154e-08, 6.47408e-08, 6.499243e-08, 6.501818e-08, 
    6.506531e-08, 6.518741e-08, 6.529008e-08, 6.508023e-08, 6.531582e-08, 
    6.443155e-08, 6.489495e-08, 6.416896e-08, 6.438758e-08, 6.453951e-08, 
    6.447286e-08, 6.481897e-08, 6.490055e-08, 6.523204e-08, 6.506068e-08, 
    6.608088e-08, 6.562952e-08, 6.688197e-08, 6.653197e-08, 6.417132e-08, 
    6.428215e-08, 6.466789e-08, 6.448436e-08, 6.500922e-08, 6.513842e-08, 
    6.524344e-08, 6.53777e-08, 6.539219e-08, 6.547174e-08, 6.534139e-08, 
    6.546659e-08, 6.499297e-08, 6.520462e-08, 6.46238e-08, 6.476517e-08, 
    6.470013e-08, 6.46288e-08, 6.484896e-08, 6.508353e-08, 6.508854e-08, 
    6.516375e-08, 6.537572e-08, 6.501136e-08, 6.613915e-08, 6.544267e-08, 
    6.440301e-08, 6.461651e-08, 6.464699e-08, 6.456429e-08, 6.512547e-08, 
    6.492213e-08, 6.54698e-08, 6.532179e-08, 6.55643e-08, 6.544379e-08, 
    6.542606e-08, 6.527128e-08, 6.517492e-08, 6.493146e-08, 6.473337e-08, 
    6.457628e-08, 6.461281e-08, 6.478536e-08, 6.509788e-08, 6.539351e-08, 
    6.532875e-08, 6.554587e-08, 6.497117e-08, 6.521216e-08, 6.511902e-08, 
    6.536187e-08, 6.482973e-08, 6.52829e-08, 6.471389e-08, 6.476378e-08, 
    6.49181e-08, 6.522851e-08, 6.529717e-08, 6.53705e-08, 6.532525e-08, 
    6.510581e-08, 6.506986e-08, 6.491435e-08, 6.487141e-08, 6.475292e-08, 
    6.465483e-08, 6.474446e-08, 6.483858e-08, 6.51059e-08, 6.53468e-08, 
    6.560944e-08, 6.567371e-08, 6.59806e-08, 6.573079e-08, 6.614304e-08, 
    6.579257e-08, 6.639924e-08, 6.530915e-08, 6.578225e-08, 6.492512e-08, 
    6.501746e-08, 6.518448e-08, 6.556754e-08, 6.536073e-08, 6.560259e-08, 
    6.506844e-08, 6.479132e-08, 6.471961e-08, 6.458583e-08, 6.472267e-08, 
    6.471154e-08, 6.484247e-08, 6.48004e-08, 6.511478e-08, 6.494591e-08, 
    6.542562e-08, 6.560068e-08, 6.609504e-08, 6.63981e-08, 6.670659e-08, 
    6.684278e-08, 6.688423e-08, 6.690156e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  8.580827e-13, 8.604064e-13, 8.599551e-13, 8.618275e-13, 8.607893e-13, 
    8.620149e-13, 8.585544e-13, 8.604983e-13, 8.592577e-13, 8.582925e-13, 
    8.654558e-13, 8.619111e-13, 8.691352e-13, 8.668784e-13, 8.725437e-13, 
    8.687836e-13, 8.733013e-13, 8.724361e-13, 8.750411e-13, 8.742953e-13, 
    8.77622e-13, 8.753853e-13, 8.793459e-13, 8.770885e-13, 8.774415e-13, 
    8.753114e-13, 8.626257e-13, 8.650145e-13, 8.624839e-13, 8.628247e-13, 
    8.62672e-13, 8.608104e-13, 8.598713e-13, 8.579055e-13, 8.582627e-13, 
    8.597067e-13, 8.62978e-13, 8.618686e-13, 8.646651e-13, 8.64602e-13, 
    8.677107e-13, 8.663096e-13, 8.715281e-13, 8.700467e-13, 8.743264e-13, 
    8.732506e-13, 8.742757e-13, 8.739651e-13, 8.742798e-13, 8.727019e-13, 
    8.73378e-13, 8.719893e-13, 8.665719e-13, 8.681653e-13, 8.634091e-13, 
    8.605431e-13, 8.586395e-13, 8.572872e-13, 8.574784e-13, 8.578427e-13, 
    8.597151e-13, 8.614749e-13, 8.628148e-13, 8.637106e-13, 8.645929e-13, 
    8.672594e-13, 8.686712e-13, 8.718272e-13, 8.712586e-13, 8.722224e-13, 
    8.731436e-13, 8.746886e-13, 8.744345e-13, 8.751147e-13, 8.721974e-13, 
    8.741364e-13, 8.70935e-13, 8.718107e-13, 8.6483e-13, 8.621681e-13, 
    8.610334e-13, 8.600417e-13, 8.576253e-13, 8.592942e-13, 8.586364e-13, 
    8.602016e-13, 8.611951e-13, 8.607039e-13, 8.637351e-13, 8.62557e-13, 
    8.687549e-13, 8.660874e-13, 8.730362e-13, 8.713754e-13, 8.734342e-13, 
    8.72384e-13, 8.741829e-13, 8.72564e-13, 8.75368e-13, 8.759778e-13, 
    8.75561e-13, 8.771624e-13, 8.724741e-13, 8.742755e-13, 8.6069e-13, 
    8.607701e-13, 8.611436e-13, 8.595013e-13, 8.594009e-13, 8.578956e-13, 
    8.592354e-13, 8.598054e-13, 8.61253e-13, 8.621082e-13, 8.629211e-13, 
    8.647075e-13, 8.667004e-13, 8.694849e-13, 8.714831e-13, 8.728217e-13, 
    8.720011e-13, 8.727256e-13, 8.719156e-13, 8.71536e-13, 8.757491e-13, 
    8.733842e-13, 8.769321e-13, 8.76736e-13, 8.751308e-13, 8.767581e-13, 
    8.608264e-13, 8.603653e-13, 8.587627e-13, 8.60017e-13, 8.577317e-13, 
    8.590108e-13, 8.597458e-13, 8.625811e-13, 8.632041e-13, 8.637809e-13, 
    8.649203e-13, 8.663813e-13, 8.689417e-13, 8.711671e-13, 8.731973e-13, 
    8.730487e-13, 8.73101e-13, 8.735541e-13, 8.724313e-13, 8.737383e-13, 
    8.739573e-13, 8.733842e-13, 8.767098e-13, 8.757602e-13, 8.767318e-13, 
    8.761137e-13, 8.605153e-13, 8.612912e-13, 8.608719e-13, 8.616601e-13, 
    8.611046e-13, 8.635729e-13, 8.643124e-13, 8.677701e-13, 8.663524e-13, 
    8.686091e-13, 8.66582e-13, 8.669411e-13, 8.686814e-13, 8.666917e-13, 
    8.710443e-13, 8.680933e-13, 8.735717e-13, 8.706275e-13, 8.73756e-13, 
    8.731886e-13, 8.741282e-13, 8.749692e-13, 8.760271e-13, 8.77977e-13, 
    8.775258e-13, 8.791559e-13, 8.624476e-13, 8.634529e-13, 8.633649e-13, 
    8.644169e-13, 8.651944e-13, 8.668793e-13, 8.695784e-13, 8.68564e-13, 
    8.704265e-13, 8.708e-13, 8.679706e-13, 8.697077e-13, 8.641258e-13, 
    8.650281e-13, 8.644913e-13, 8.625267e-13, 8.687971e-13, 8.65581e-13, 
    8.71516e-13, 8.697771e-13, 8.748492e-13, 8.723274e-13, 8.772771e-13, 
    8.793883e-13, 8.813757e-13, 8.836929e-13, 8.640019e-13, 8.63319e-13, 
    8.645421e-13, 8.662322e-13, 8.678005e-13, 8.698832e-13, 8.700964e-13, 
    8.704861e-13, 8.714955e-13, 8.72344e-13, 8.706088e-13, 8.725566e-13, 
    8.652363e-13, 8.690762e-13, 8.630603e-13, 8.648729e-13, 8.661328e-13, 
    8.655807e-13, 8.684481e-13, 8.691232e-13, 8.718637e-13, 8.70448e-13, 
    8.78867e-13, 8.751459e-13, 8.854573e-13, 8.825805e-13, 8.630802e-13, 
    8.639998e-13, 8.671964e-13, 8.656761e-13, 8.700224e-13, 8.710906e-13, 
    8.719586e-13, 8.730675e-13, 8.731875e-13, 8.738443e-13, 8.727679e-13, 
    8.73802e-13, 8.698875e-13, 8.716375e-13, 8.668319e-13, 8.680023e-13, 
    8.674641e-13, 8.668733e-13, 8.686963e-13, 8.70636e-13, 8.706783e-13, 
    8.712993e-13, 8.730481e-13, 8.700399e-13, 8.793452e-13, 8.736015e-13, 
    8.65002e-13, 8.667702e-13, 8.670236e-13, 8.663388e-13, 8.709835e-13, 
    8.693016e-13, 8.738284e-13, 8.726059e-13, 8.746088e-13, 8.736137e-13, 
    8.734672e-13, 8.721886e-13, 8.713919e-13, 8.693786e-13, 8.677389e-13, 
    8.664382e-13, 8.667408e-13, 8.681694e-13, 8.707548e-13, 8.731981e-13, 
    8.726628e-13, 8.744566e-13, 8.697075e-13, 8.716995e-13, 8.709298e-13, 
    8.72937e-13, 8.685368e-13, 8.722818e-13, 8.675781e-13, 8.679911e-13, 
    8.692682e-13, 8.71834e-13, 8.724025e-13, 8.73008e-13, 8.726346e-13, 
    8.708206e-13, 8.705235e-13, 8.692374e-13, 8.688817e-13, 8.679013e-13, 
    8.670888e-13, 8.678309e-13, 8.686098e-13, 8.708217e-13, 8.728121e-13, 
    8.74981e-13, 8.755117e-13, 8.780403e-13, 8.75981e-13, 8.79377e-13, 
    8.764883e-13, 8.814871e-13, 8.724998e-13, 8.764051e-13, 8.693266e-13, 
    8.700905e-13, 8.714702e-13, 8.746343e-13, 8.729275e-13, 8.749238e-13, 
    8.70512e-13, 8.682182e-13, 8.676254e-13, 8.665172e-13, 8.676507e-13, 
    8.675586e-13, 8.686427e-13, 8.682944e-13, 8.708951e-13, 8.694985e-13, 
    8.734633e-13, 8.749083e-13, 8.789848e-13, 8.814794e-13, 8.84017e-13, 
    8.851359e-13, 8.854764e-13, 8.856186e-13 ;

 LITR1C =
  3.066807e-05, 3.066795e-05, 3.066798e-05, 3.066788e-05, 3.066794e-05, 
    3.066787e-05, 3.066805e-05, 3.066795e-05, 3.066801e-05, 3.066806e-05, 
    3.06677e-05, 3.066788e-05, 3.066752e-05, 3.066763e-05, 3.066735e-05, 
    3.066753e-05, 3.066731e-05, 3.066735e-05, 3.066722e-05, 3.066726e-05, 
    3.066709e-05, 3.06672e-05, 3.0667e-05, 3.066712e-05, 3.06671e-05, 
    3.06672e-05, 3.066784e-05, 3.066772e-05, 3.066785e-05, 3.066783e-05, 
    3.066784e-05, 3.066794e-05, 3.066798e-05, 3.066808e-05, 3.066806e-05, 
    3.066799e-05, 3.066783e-05, 3.066788e-05, 3.066774e-05, 3.066774e-05, 
    3.066759e-05, 3.066766e-05, 3.06674e-05, 3.066747e-05, 3.066726e-05, 
    3.066731e-05, 3.066726e-05, 3.066727e-05, 3.066726e-05, 3.066734e-05, 
    3.06673e-05, 3.066737e-05, 3.066764e-05, 3.066756e-05, 3.06678e-05, 
    3.066795e-05, 3.066804e-05, 3.066811e-05, 3.06681e-05, 3.066808e-05, 
    3.066799e-05, 3.06679e-05, 3.066783e-05, 3.066779e-05, 3.066774e-05, 
    3.066761e-05, 3.066754e-05, 3.066738e-05, 3.066741e-05, 3.066736e-05, 
    3.066731e-05, 3.066724e-05, 3.066725e-05, 3.066722e-05, 3.066736e-05, 
    3.066727e-05, 3.066743e-05, 3.066738e-05, 3.066773e-05, 3.066787e-05, 
    3.066792e-05, 3.066797e-05, 3.06681e-05, 3.066801e-05, 3.066804e-05, 
    3.066796e-05, 3.066791e-05, 3.066794e-05, 3.066779e-05, 3.066784e-05, 
    3.066754e-05, 3.066767e-05, 3.066732e-05, 3.06674e-05, 3.06673e-05, 
    3.066735e-05, 3.066726e-05, 3.066734e-05, 3.06672e-05, 3.066717e-05, 
    3.066719e-05, 3.066711e-05, 3.066735e-05, 3.066726e-05, 3.066794e-05, 
    3.066794e-05, 3.066792e-05, 3.0668e-05, 3.0668e-05, 3.066808e-05, 
    3.066801e-05, 3.066798e-05, 3.066791e-05, 3.066787e-05, 3.066783e-05, 
    3.066774e-05, 3.066764e-05, 3.06675e-05, 3.06674e-05, 3.066733e-05, 
    3.066737e-05, 3.066734e-05, 3.066738e-05, 3.066739e-05, 3.066718e-05, 
    3.06673e-05, 3.066712e-05, 3.066714e-05, 3.066722e-05, 3.066713e-05, 
    3.066793e-05, 3.066796e-05, 3.066804e-05, 3.066798e-05, 3.066809e-05, 
    3.066802e-05, 3.066799e-05, 3.066784e-05, 3.066782e-05, 3.066779e-05, 
    3.066773e-05, 3.066766e-05, 3.066752e-05, 3.066742e-05, 3.066731e-05, 
    3.066732e-05, 3.066732e-05, 3.06673e-05, 3.066735e-05, 3.066728e-05, 
    3.066727e-05, 3.06673e-05, 3.066714e-05, 3.066718e-05, 3.066714e-05, 
    3.066716e-05, 3.066795e-05, 3.066791e-05, 3.066793e-05, 3.066789e-05, 
    3.066792e-05, 3.066779e-05, 3.066776e-05, 3.066758e-05, 3.066766e-05, 
    3.066754e-05, 3.066764e-05, 3.066763e-05, 3.066754e-05, 3.066764e-05, 
    3.066742e-05, 3.066757e-05, 3.066729e-05, 3.066744e-05, 3.066728e-05, 
    3.066731e-05, 3.066727e-05, 3.066722e-05, 3.066717e-05, 3.066707e-05, 
    3.06671e-05, 3.066701e-05, 3.066785e-05, 3.06678e-05, 3.06678e-05, 
    3.066775e-05, 3.066771e-05, 3.066763e-05, 3.06675e-05, 3.066755e-05, 
    3.066745e-05, 3.066743e-05, 3.066758e-05, 3.066749e-05, 3.066777e-05, 
    3.066772e-05, 3.066775e-05, 3.066785e-05, 3.066753e-05, 3.06677e-05, 
    3.06674e-05, 3.066748e-05, 3.066723e-05, 3.066736e-05, 3.066711e-05, 
    3.0667e-05, 3.06669e-05, 3.066679e-05, 3.066777e-05, 3.066781e-05, 
    3.066775e-05, 3.066766e-05, 3.066758e-05, 3.066748e-05, 3.066747e-05, 
    3.066745e-05, 3.06674e-05, 3.066735e-05, 3.066744e-05, 3.066734e-05, 
    3.066771e-05, 3.066752e-05, 3.066782e-05, 3.066773e-05, 3.066767e-05, 
    3.06677e-05, 3.066755e-05, 3.066752e-05, 3.066738e-05, 3.066745e-05, 
    3.066703e-05, 3.066722e-05, 3.06667e-05, 3.066684e-05, 3.066782e-05, 
    3.066778e-05, 3.066761e-05, 3.066769e-05, 3.066747e-05, 3.066742e-05, 
    3.066738e-05, 3.066732e-05, 3.066731e-05, 3.066728e-05, 3.066733e-05, 
    3.066728e-05, 3.066748e-05, 3.066739e-05, 3.066763e-05, 3.066757e-05, 
    3.06676e-05, 3.066763e-05, 3.066754e-05, 3.066744e-05, 3.066744e-05, 
    3.066741e-05, 3.066732e-05, 3.066747e-05, 3.0667e-05, 3.066729e-05, 
    3.066772e-05, 3.066763e-05, 3.066762e-05, 3.066766e-05, 3.066742e-05, 
    3.066751e-05, 3.066728e-05, 3.066734e-05, 3.066724e-05, 3.066729e-05, 
    3.06673e-05, 3.066736e-05, 3.06674e-05, 3.06675e-05, 3.066759e-05, 
    3.066765e-05, 3.066764e-05, 3.066756e-05, 3.066743e-05, 3.066731e-05, 
    3.066734e-05, 3.066725e-05, 3.066749e-05, 3.066739e-05, 3.066743e-05, 
    3.066732e-05, 3.066755e-05, 3.066736e-05, 3.066759e-05, 3.066757e-05, 
    3.066751e-05, 3.066738e-05, 3.066735e-05, 3.066732e-05, 3.066734e-05, 
    3.066743e-05, 3.066744e-05, 3.066751e-05, 3.066753e-05, 3.066758e-05, 
    3.066762e-05, 3.066758e-05, 3.066754e-05, 3.066743e-05, 3.066733e-05, 
    3.066722e-05, 3.06672e-05, 3.066707e-05, 3.066717e-05, 3.0667e-05, 
    3.066715e-05, 3.06669e-05, 3.066735e-05, 3.066715e-05, 3.066751e-05, 
    3.066747e-05, 3.06674e-05, 3.066724e-05, 3.066732e-05, 3.066723e-05, 
    3.066745e-05, 3.066756e-05, 3.066759e-05, 3.066765e-05, 3.066759e-05, 
    3.066759e-05, 3.066754e-05, 3.066756e-05, 3.066743e-05, 3.06675e-05, 
    3.06673e-05, 3.066723e-05, 3.066702e-05, 3.06669e-05, 3.066677e-05, 
    3.066671e-05, 3.06667e-05, 3.066669e-05 ;

 LITR1C_TO_SOIL1C =
  5.715241e-13, 5.730715e-13, 5.727709e-13, 5.740178e-13, 5.733265e-13, 
    5.741426e-13, 5.718381e-13, 5.731327e-13, 5.723065e-13, 5.716638e-13, 
    5.76434e-13, 5.740735e-13, 5.788842e-13, 5.773814e-13, 5.81154e-13, 
    5.786501e-13, 5.816586e-13, 5.810824e-13, 5.828172e-13, 5.823204e-13, 
    5.845358e-13, 5.830464e-13, 5.856837e-13, 5.841805e-13, 5.844156e-13, 
    5.829971e-13, 5.745494e-13, 5.761402e-13, 5.744549e-13, 5.746819e-13, 
    5.745802e-13, 5.733406e-13, 5.727152e-13, 5.714061e-13, 5.716439e-13, 
    5.726055e-13, 5.74784e-13, 5.740452e-13, 5.759075e-13, 5.758655e-13, 
    5.779356e-13, 5.770026e-13, 5.804777e-13, 5.794912e-13, 5.823412e-13, 
    5.816248e-13, 5.823074e-13, 5.821006e-13, 5.823101e-13, 5.812594e-13, 
    5.817096e-13, 5.807849e-13, 5.771772e-13, 5.782384e-13, 5.750711e-13, 
    5.731625e-13, 5.718949e-13, 5.709943e-13, 5.711217e-13, 5.713642e-13, 
    5.726112e-13, 5.73783e-13, 5.746753e-13, 5.752718e-13, 5.758594e-13, 
    5.776351e-13, 5.785752e-13, 5.806769e-13, 5.802983e-13, 5.8094e-13, 
    5.815535e-13, 5.825824e-13, 5.824131e-13, 5.828661e-13, 5.809234e-13, 
    5.822147e-13, 5.800827e-13, 5.806659e-13, 5.760173e-13, 5.742446e-13, 
    5.73489e-13, 5.728286e-13, 5.712195e-13, 5.723308e-13, 5.718928e-13, 
    5.729351e-13, 5.735967e-13, 5.732696e-13, 5.752881e-13, 5.745036e-13, 
    5.786309e-13, 5.768546e-13, 5.81482e-13, 5.80376e-13, 5.817471e-13, 
    5.810477e-13, 5.822456e-13, 5.811675e-13, 5.830348e-13, 5.834408e-13, 
    5.831633e-13, 5.842297e-13, 5.811077e-13, 5.823073e-13, 5.732604e-13, 
    5.733137e-13, 5.735624e-13, 5.724687e-13, 5.724019e-13, 5.713995e-13, 
    5.722917e-13, 5.726713e-13, 5.736352e-13, 5.742048e-13, 5.747461e-13, 
    5.759357e-13, 5.772628e-13, 5.79117e-13, 5.804477e-13, 5.813392e-13, 
    5.807927e-13, 5.812752e-13, 5.807358e-13, 5.80483e-13, 5.832886e-13, 
    5.817137e-13, 5.840764e-13, 5.839458e-13, 5.828768e-13, 5.839605e-13, 
    5.733512e-13, 5.730441e-13, 5.719769e-13, 5.728121e-13, 5.712903e-13, 
    5.721421e-13, 5.726316e-13, 5.745197e-13, 5.749346e-13, 5.753187e-13, 
    5.760774e-13, 5.770503e-13, 5.787554e-13, 5.802373e-13, 5.815893e-13, 
    5.814903e-13, 5.815252e-13, 5.818269e-13, 5.810792e-13, 5.819496e-13, 
    5.820954e-13, 5.817138e-13, 5.839283e-13, 5.83296e-13, 5.839431e-13, 
    5.835314e-13, 5.73144e-13, 5.736607e-13, 5.733815e-13, 5.739064e-13, 
    5.735364e-13, 5.751801e-13, 5.756726e-13, 5.779752e-13, 5.770311e-13, 
    5.785339e-13, 5.77184e-13, 5.774231e-13, 5.78582e-13, 5.77257e-13, 
    5.801556e-13, 5.781904e-13, 5.818386e-13, 5.79878e-13, 5.819613e-13, 
    5.815834e-13, 5.822092e-13, 5.827692e-13, 5.834737e-13, 5.847722e-13, 
    5.844717e-13, 5.855572e-13, 5.744308e-13, 5.751002e-13, 5.750416e-13, 
    5.757421e-13, 5.7626e-13, 5.773819e-13, 5.791793e-13, 5.785038e-13, 
    5.797441e-13, 5.799929e-13, 5.781086e-13, 5.792655e-13, 5.755483e-13, 
    5.761492e-13, 5.757917e-13, 5.744834e-13, 5.78659e-13, 5.765174e-13, 
    5.804696e-13, 5.793117e-13, 5.826893e-13, 5.8101e-13, 5.843061e-13, 
    5.85712e-13, 5.870355e-13, 5.885786e-13, 5.754658e-13, 5.750111e-13, 
    5.758255e-13, 5.76951e-13, 5.779954e-13, 5.793823e-13, 5.795243e-13, 
    5.797838e-13, 5.80456e-13, 5.81021e-13, 5.798656e-13, 5.811627e-13, 
    5.762878e-13, 5.78845e-13, 5.748388e-13, 5.760458e-13, 5.768848e-13, 
    5.765172e-13, 5.784267e-13, 5.788762e-13, 5.807012e-13, 5.797585e-13, 
    5.853649e-13, 5.828869e-13, 5.897535e-13, 5.878378e-13, 5.748521e-13, 
    5.754644e-13, 5.775931e-13, 5.765808e-13, 5.79475e-13, 5.801864e-13, 
    5.807644e-13, 5.815028e-13, 5.815828e-13, 5.820201e-13, 5.813033e-13, 
    5.81992e-13, 5.793852e-13, 5.805506e-13, 5.773504e-13, 5.781298e-13, 
    5.777714e-13, 5.773779e-13, 5.78592e-13, 5.798837e-13, 5.799118e-13, 
    5.803253e-13, 5.814899e-13, 5.794867e-13, 5.856833e-13, 5.818585e-13, 
    5.761319e-13, 5.773093e-13, 5.774781e-13, 5.77022e-13, 5.801151e-13, 
    5.78995e-13, 5.820095e-13, 5.811955e-13, 5.825292e-13, 5.818666e-13, 
    5.81769e-13, 5.809176e-13, 5.80387e-13, 5.790463e-13, 5.779544e-13, 
    5.770882e-13, 5.772897e-13, 5.78241e-13, 5.799628e-13, 5.815898e-13, 
    5.812334e-13, 5.824279e-13, 5.792653e-13, 5.805918e-13, 5.800793e-13, 
    5.814159e-13, 5.784857e-13, 5.809796e-13, 5.778473e-13, 5.781223e-13, 
    5.789728e-13, 5.806814e-13, 5.8106e-13, 5.814632e-13, 5.812145e-13, 
    5.800066e-13, 5.798088e-13, 5.789523e-13, 5.787154e-13, 5.780626e-13, 
    5.775215e-13, 5.780157e-13, 5.785343e-13, 5.800073e-13, 5.813328e-13, 
    5.82777e-13, 5.831305e-13, 5.848144e-13, 5.83443e-13, 5.857044e-13, 
    5.837809e-13, 5.871096e-13, 5.811248e-13, 5.837254e-13, 5.790117e-13, 
    5.795204e-13, 5.804392e-13, 5.825462e-13, 5.814096e-13, 5.82739e-13, 
    5.798011e-13, 5.782735e-13, 5.778788e-13, 5.771408e-13, 5.778956e-13, 
    5.778343e-13, 5.785562e-13, 5.783243e-13, 5.800562e-13, 5.791262e-13, 
    5.817664e-13, 5.827287e-13, 5.854433e-13, 5.871045e-13, 5.887944e-13, 
    5.895394e-13, 5.897662e-13, 5.898609e-13 ;

 LITR1C_vr =
  0.001751179, 0.001751172, 0.001751173, 0.001751168, 0.001751171, 
    0.001751167, 0.001751177, 0.001751172, 0.001751175, 0.001751178, 
    0.001751157, 0.001751168, 0.001751147, 0.001751153, 0.001751137, 
    0.001751148, 0.001751135, 0.001751137, 0.00175113, 0.001751132, 
    0.001751123, 0.001751129, 0.001751118, 0.001751124, 0.001751123, 
    0.001751129, 0.001751165, 0.001751159, 0.001751166, 0.001751165, 
    0.001751165, 0.001751171, 0.001751173, 0.001751179, 0.001751178, 
    0.001751174, 0.001751165, 0.001751168, 0.00175116, 0.00175116, 
    0.001751151, 0.001751155, 0.00175114, 0.001751144, 0.001751132, 
    0.001751135, 0.001751132, 0.001751133, 0.001751132, 0.001751137, 
    0.001751135, 0.001751139, 0.001751154, 0.00175115, 0.001751163, 
    0.001751172, 0.001751177, 0.001751181, 0.00175118, 0.001751179, 
    0.001751174, 0.001751169, 0.001751165, 0.001751162, 0.00175116, 
    0.001751152, 0.001751148, 0.001751139, 0.001751141, 0.001751138, 
    0.001751135, 0.001751131, 0.001751132, 0.00175113, 0.001751138, 
    0.001751133, 0.001751142, 0.001751139, 0.001751159, 0.001751167, 
    0.00175117, 0.001751173, 0.00175118, 0.001751175, 0.001751177, 
    0.001751172, 0.00175117, 0.001751171, 0.001751162, 0.001751166, 
    0.001751148, 0.001751156, 0.001751136, 0.00175114, 0.001751135, 
    0.001751138, 0.001751132, 0.001751137, 0.001751129, 0.001751127, 
    0.001751128, 0.001751124, 0.001751137, 0.001751132, 0.001751171, 
    0.001751171, 0.00175117, 0.001751174, 0.001751175, 0.001751179, 
    0.001751175, 0.001751174, 0.001751169, 0.001751167, 0.001751165, 
    0.00175116, 0.001751154, 0.001751146, 0.00175114, 0.001751136, 
    0.001751139, 0.001751137, 0.001751139, 0.00175114, 0.001751128, 
    0.001751135, 0.001751125, 0.001751125, 0.00175113, 0.001751125, 
    0.001751171, 0.001751172, 0.001751177, 0.001751173, 0.00175118, 
    0.001751176, 0.001751174, 0.001751166, 0.001751164, 0.001751162, 
    0.001751159, 0.001751155, 0.001751147, 0.001751141, 0.001751135, 
    0.001751136, 0.001751135, 0.001751134, 0.001751137, 0.001751134, 
    0.001751133, 0.001751135, 0.001751125, 0.001751128, 0.001751125, 
    0.001751127, 0.001751172, 0.001751169, 0.001751171, 0.001751168, 
    0.00175117, 0.001751163, 0.001751161, 0.001751151, 0.001751155, 
    0.001751148, 0.001751154, 0.001751153, 0.001751148, 0.001751154, 
    0.001751141, 0.00175115, 0.001751134, 0.001751143, 0.001751134, 
    0.001751135, 0.001751133, 0.00175113, 0.001751127, 0.001751121, 
    0.001751123, 0.001751118, 0.001751166, 0.001751163, 0.001751163, 
    0.00175116, 0.001751158, 0.001751153, 0.001751146, 0.001751148, 
    0.001751143, 0.001751142, 0.00175115, 0.001751145, 0.001751161, 
    0.001751159, 0.00175116, 0.001751166, 0.001751148, 0.001751157, 
    0.00175114, 0.001751145, 0.00175113, 0.001751138, 0.001751123, 
    0.001751117, 0.001751112, 0.001751105, 0.001751162, 0.001751164, 
    0.00175116, 0.001751155, 0.001751151, 0.001751145, 0.001751144, 
    0.001751143, 0.00175114, 0.001751138, 0.001751143, 0.001751137, 
    0.001751158, 0.001751147, 0.001751164, 0.001751159, 0.001751155, 
    0.001751157, 0.001751149, 0.001751147, 0.001751139, 0.001751143, 
    0.001751119, 0.00175113, 0.0017511, 0.001751108, 0.001751164, 
    0.001751162, 0.001751152, 0.001751157, 0.001751144, 0.001751141, 
    0.001751139, 0.001751136, 0.001751135, 0.001751133, 0.001751136, 
    0.001751133, 0.001751145, 0.00175114, 0.001751153, 0.00175115, 
    0.001751152, 0.001751153, 0.001751148, 0.001751143, 0.001751142, 
    0.001751141, 0.001751136, 0.001751144, 0.001751118, 0.001751134, 
    0.001751159, 0.001751154, 0.001751153, 0.001751155, 0.001751142, 
    0.001751146, 0.001751133, 0.001751137, 0.001751131, 0.001751134, 
    0.001751134, 0.001751138, 0.00175114, 0.001751146, 0.001751151, 
    0.001751155, 0.001751154, 0.00175115, 0.001751142, 0.001751135, 
    0.001751137, 0.001751132, 0.001751145, 0.00175114, 0.001751142, 
    0.001751136, 0.001751149, 0.001751138, 0.001751151, 0.00175115, 
    0.001751147, 0.001751139, 0.001751137, 0.001751136, 0.001751137, 
    0.001751142, 0.001751143, 0.001751147, 0.001751148, 0.00175115, 
    0.001751153, 0.001751151, 0.001751148, 0.001751142, 0.001751136, 
    0.00175113, 0.001751129, 0.001751121, 0.001751127, 0.001751118, 
    0.001751126, 0.001751111, 0.001751137, 0.001751126, 0.001751146, 
    0.001751144, 0.00175114, 0.001751131, 0.001751136, 0.00175113, 
    0.001751143, 0.00175115, 0.001751151, 0.001751154, 0.001751151, 
    0.001751151, 0.001751148, 0.001751149, 0.001751142, 0.001751146, 
    0.001751134, 0.00175113, 0.001751119, 0.001751111, 0.001751104, 
    0.001751101, 0.0017511, 0.0017511,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732906e-07, 9.73287e-07, 9.732877e-07, 9.732847e-07, 9.732863e-07, 
    9.732844e-07, 9.7329e-07, 9.732868e-07, 9.732888e-07, 9.732903e-07, 
    9.732789e-07, 9.732846e-07, 9.73273e-07, 9.732767e-07, 9.732676e-07, 
    9.732736e-07, 9.732664e-07, 9.732678e-07, 9.732636e-07, 9.732648e-07, 
    9.732595e-07, 9.732631e-07, 9.732568e-07, 9.732604e-07, 9.732598e-07, 
    9.732632e-07, 9.732834e-07, 9.732796e-07, 9.732836e-07, 9.732831e-07, 
    9.732834e-07, 9.732863e-07, 9.732878e-07, 9.73291e-07, 9.732904e-07, 
    9.73288e-07, 9.732829e-07, 9.732846e-07, 9.732802e-07, 9.732803e-07, 
    9.732753e-07, 9.732776e-07, 9.732693e-07, 9.732715e-07, 9.732647e-07, 
    9.732665e-07, 9.732648e-07, 9.732654e-07, 9.732648e-07, 9.732673e-07, 
    9.732663e-07, 9.732685e-07, 9.732771e-07, 9.732746e-07, 9.732822e-07, 
    9.732868e-07, 9.732897e-07, 9.732919e-07, 9.732917e-07, 9.732911e-07, 
    9.73288e-07, 9.732853e-07, 9.732831e-07, 9.732817e-07, 9.732803e-07, 
    9.73276e-07, 9.732738e-07, 9.732687e-07, 9.732696e-07, 9.732681e-07, 
    9.732667e-07, 9.732642e-07, 9.732646e-07, 9.732635e-07, 9.732681e-07, 
    9.732651e-07, 9.732702e-07, 9.732688e-07, 9.7328e-07, 9.732842e-07, 
    9.73286e-07, 9.732876e-07, 9.732914e-07, 9.732887e-07, 9.732897e-07, 
    9.732872e-07, 9.732858e-07, 9.732864e-07, 9.732817e-07, 9.732835e-07, 
    9.732737e-07, 9.732779e-07, 9.732669e-07, 9.732695e-07, 9.732662e-07, 
    9.732679e-07, 9.732649e-07, 9.732676e-07, 9.732631e-07, 9.732621e-07, 
    9.732628e-07, 9.732603e-07, 9.732677e-07, 9.732648e-07, 9.732865e-07, 
    9.732864e-07, 9.732858e-07, 9.732884e-07, 9.732886e-07, 9.73291e-07, 
    9.732888e-07, 9.732879e-07, 9.732856e-07, 9.732843e-07, 9.732829e-07, 
    9.732801e-07, 9.732769e-07, 9.732724e-07, 9.732693e-07, 9.732672e-07, 
    9.732685e-07, 9.732673e-07, 9.732686e-07, 9.732693e-07, 9.732626e-07, 
    9.732663e-07, 9.732606e-07, 9.73261e-07, 9.732635e-07, 9.732609e-07, 
    9.732863e-07, 9.73287e-07, 9.732896e-07, 9.732876e-07, 9.732912e-07, 
    9.732892e-07, 9.73288e-07, 9.732835e-07, 9.732825e-07, 9.732815e-07, 
    9.732797e-07, 9.732775e-07, 9.732734e-07, 9.732698e-07, 9.732665e-07, 
    9.732668e-07, 9.732668e-07, 9.73266e-07, 9.732678e-07, 9.732657e-07, 
    9.732654e-07, 9.732663e-07, 9.73261e-07, 9.732624e-07, 9.73261e-07, 
    9.732619e-07, 9.732868e-07, 9.732855e-07, 9.732862e-07, 9.73285e-07, 
    9.732859e-07, 9.732819e-07, 9.732807e-07, 9.732752e-07, 9.732775e-07, 
    9.732739e-07, 9.732771e-07, 9.732765e-07, 9.732738e-07, 9.732769e-07, 
    9.732699e-07, 9.732747e-07, 9.73266e-07, 9.732706e-07, 9.732656e-07, 
    9.732665e-07, 9.732651e-07, 9.732637e-07, 9.732621e-07, 9.732589e-07, 
    9.732597e-07, 9.732571e-07, 9.732837e-07, 9.732821e-07, 9.732822e-07, 
    9.732805e-07, 9.732793e-07, 9.732767e-07, 9.732723e-07, 9.732739e-07, 
    9.73271e-07, 9.732704e-07, 9.73275e-07, 9.732721e-07, 9.73281e-07, 
    9.732796e-07, 9.732804e-07, 9.732836e-07, 9.732736e-07, 9.732787e-07, 
    9.732693e-07, 9.73272e-07, 9.732639e-07, 9.732679e-07, 9.732601e-07, 
    9.732566e-07, 9.732536e-07, 9.732498e-07, 9.732812e-07, 9.732823e-07, 
    9.732804e-07, 9.732777e-07, 9.732752e-07, 9.732719e-07, 9.732715e-07, 
    9.732709e-07, 9.732693e-07, 9.732679e-07, 9.732707e-07, 9.732676e-07, 
    9.732793e-07, 9.732731e-07, 9.732827e-07, 9.732798e-07, 9.732778e-07, 
    9.732787e-07, 9.732742e-07, 9.73273e-07, 9.732687e-07, 9.73271e-07, 
    9.732576e-07, 9.732635e-07, 9.73247e-07, 9.732516e-07, 9.732827e-07, 
    9.732812e-07, 9.732761e-07, 9.732786e-07, 9.732717e-07, 9.732699e-07, 
    9.732686e-07, 9.732668e-07, 9.732665e-07, 9.732655e-07, 9.732672e-07, 
    9.732656e-07, 9.732719e-07, 9.73269e-07, 9.732768e-07, 9.732748e-07, 
    9.732757e-07, 9.732767e-07, 9.732737e-07, 9.732706e-07, 9.732706e-07, 
    9.732696e-07, 9.732668e-07, 9.732717e-07, 9.732568e-07, 9.73266e-07, 
    9.732796e-07, 9.732768e-07, 9.732764e-07, 9.732775e-07, 9.732701e-07, 
    9.732728e-07, 9.732655e-07, 9.732676e-07, 9.732643e-07, 9.732659e-07, 
    9.732661e-07, 9.732681e-07, 9.732695e-07, 9.732727e-07, 9.732753e-07, 
    9.732773e-07, 9.732769e-07, 9.732746e-07, 9.732705e-07, 9.732665e-07, 
    9.732674e-07, 9.732646e-07, 9.732721e-07, 9.732689e-07, 9.732702e-07, 
    9.73267e-07, 9.73274e-07, 9.73268e-07, 9.732755e-07, 9.732748e-07, 
    9.732728e-07, 9.732687e-07, 9.732678e-07, 9.732669e-07, 9.732674e-07, 
    9.732704e-07, 9.732709e-07, 9.732729e-07, 9.732735e-07, 9.732751e-07, 
    9.732763e-07, 9.732752e-07, 9.732739e-07, 9.732704e-07, 9.732672e-07, 
    9.732637e-07, 9.732629e-07, 9.732588e-07, 9.732621e-07, 9.732568e-07, 
    9.732613e-07, 9.732533e-07, 9.732677e-07, 9.732614e-07, 9.732728e-07, 
    9.732715e-07, 9.732693e-07, 9.732643e-07, 9.73267e-07, 9.732638e-07, 
    9.732709e-07, 9.732745e-07, 9.732754e-07, 9.732772e-07, 9.732754e-07, 
    9.732755e-07, 9.732738e-07, 9.732744e-07, 9.732703e-07, 9.732724e-07, 
    9.732662e-07, 9.732638e-07, 9.732573e-07, 9.732533e-07, 9.732494e-07, 
    9.732476e-07, 9.73247e-07, 9.732468e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  5.391992e-25, -6.764499e-25, 1.56858e-25, 2.941087e-25, 1.235256e-24, 
    -2.745014e-25, -4.117521e-25, 8.82326e-26, 1.02938e-24, 2.646978e-25, 
    2.450906e-25, -2.941087e-25, 7.25468e-25, 2.450906e-25, 6.666463e-25, 
    -7.352717e-25, 2.941087e-26, -1.078398e-25, 9.411477e-25, -9.313441e-25, 
    -3.088141e-25, 1.372507e-25, -1.764652e-25, 3.137159e-25, -3.431268e-26, 
    -4.901811e-26, 6.666463e-25, -2.450906e-25, 5.931191e-25, -2.548942e-25, 
    3.62734e-25, 4.901811e-27, 4.41163e-26, 7.842898e-26, -2.695996e-25, 
    -5.882173e-26, 1.176435e-25, 1.470543e-25, 4.215557e-25, 0, 
    -2.156797e-25, 1.176435e-25, -8.03897e-25, -7.842898e-26, -1.470543e-25, 
    5.048866e-25, 7.842898e-26, 4.803775e-25, 4.901811e-26, 9.803622e-27, 
    -2.450906e-25, 6.176282e-25, -6.862535e-26, 3.137159e-25, -2.058761e-25, 
    9.117368e-25, 4.803775e-25, 6.862535e-25, -5.98021e-25, 2.156797e-25, 
    1.323489e-25, -2.941087e-25, 3.431268e-25, 6.666463e-25, 4.117521e-25, 
    -9.901658e-25, 5.98021e-25, -1.176435e-25, 1.176435e-25, -1.81367e-25, 
    4.852793e-25, -8.725224e-25, 2.450906e-25, -6.372354e-26, 8.82326e-26, 
    -2.695996e-25, -4.901811e-25, -7.842898e-25, -2.794032e-25, 
    -3.823413e-25, -2.352869e-25, 6.862535e-26, 6.078246e-25, -2.009742e-25, 
    4.852793e-25, 4.65672e-25, 1.039184e-24, -6.862535e-26, 5.637083e-25, 
    1.176435e-25, -4.852793e-25, 5.539047e-25, -1.960724e-25, 1.176435e-25, 
    -3.921449e-25, 5.19592e-25, -1.960724e-26, -1.470543e-25, -6.568427e-25, 
    -1.02938e-24, -8.03897e-25, 5.882173e-26, 1.960724e-26, 7.352717e-26, 
    -6.274318e-25, 6.078246e-25, -1.862688e-25, 3.137159e-25, -5.048866e-25, 
    3.431268e-25, -7.842898e-25, -1.323489e-25, 2.254833e-25, 6.372354e-26, 
    -2.843051e-25, -2.156797e-25, 1.470543e-25, 3.725376e-25, 3.235195e-25, 
    -4.460648e-25, 4.65672e-25, -1.960724e-26, 9.313441e-26, 6.47039e-25, 
    3.823413e-25, 1.470543e-25, 3.088141e-25, 1.176435e-25, 9.313441e-25, 
    -2.352869e-25, 5.44101e-25, -4.362612e-25, -1.960724e-26, 4.754757e-25, 
    2.303851e-25, -9.803622e-27, -8.431115e-25, -7.107626e-25, 4.117521e-25, 
    8.725224e-25, -1.519561e-25, -5.882173e-25, 3.186177e-25, 3.431268e-25, 
    3.039123e-25, 3.039123e-25, -2.745014e-25, -3.186177e-25, 5.391992e-26, 
    3.235195e-25, 4.41163e-25, -4.215557e-25, -1.372507e-25, -2.450906e-25, 
    -6.127264e-25, 6.862535e-26, -3.921449e-25, -9.803622e-26, 1.470543e-25, 
    -5.882173e-26, -1.960724e-26, -6.617445e-25, 1.078398e-25, -4.705739e-25, 
    -4.215557e-25, 1.960724e-25, -6.323336e-25, -7.940934e-25, -7.352717e-26, 
    -2.352869e-25, -8.921296e-25, 7.058608e-25, 1.666616e-25, 4.019485e-25, 
    4.950829e-25, -2.941087e-26, 2.843051e-25, -4.264576e-25, 5.686101e-25, 
    -1.078398e-25, 3.921449e-25, -2.646978e-25, -4.41163e-25, -8.82326e-26, 
    -5.588064e-25, -3.921449e-26, 1.274471e-25, 2.254833e-25, -3.725376e-25, 
    1.666616e-25, 2.352869e-25, -4.803775e-25, 6.2253e-25, 9.313441e-26, 
    3.38225e-25, 4.999847e-25, 4.852793e-25, 1.617598e-25, -2.548942e-25, 
    8.431115e-25, 6.47039e-25, -1.274471e-25, -4.901811e-25, 3.921449e-25, 
    -9.803622e-27, 6.122413e-41, -7.842898e-26, 1.960724e-25, 7.646825e-25, 
    -2.156797e-25, -1.862688e-25, -2.941087e-26, 8.284061e-25, 1.048988e-24, 
    1.127417e-24, 3.823413e-25, -3.921449e-26, -3.921449e-25, 2.303851e-25, 
    -5.98021e-25, -1.421525e-25, 2.401887e-25, 9.803622e-26, -4.607703e-25, 
    -5.391992e-25, -2.941087e-26, 7.058608e-25, 5.686101e-25, -1.666616e-25, 
    -4.068503e-25, -4.215557e-25, -5.784137e-25, 7.842898e-26, 3.872431e-25, 
    3.039123e-25, -5.882173e-25, 4.509666e-25, 2.941087e-25, 1.715634e-25, 
    1.666616e-25, -2.548942e-25, 3.333231e-25, -4.117521e-25, -3.823413e-25, 
    -3.137159e-25, 3.235195e-25, 5.19592e-25, 7.548789e-25, 1.274471e-25, 
    6.274318e-25, -5.097883e-25, 2.843051e-25, -9.60755e-25, 1.372507e-25, 
    1.960724e-26, 5.490028e-25, 7.25468e-25, -6.176282e-25, 5.097883e-25, 
    -4.41163e-26, -2.352869e-25, -1.078398e-25, -6.274318e-25, -9.803622e-25, 
    2.450906e-25, -2.156797e-25, -2.941087e-25, 6.862535e-25, -1.078398e-25, 
    8.333079e-25, -1.039184e-24, 1.56858e-25, 5.097883e-25, -1.666616e-25, 
    -2.450906e-25, -4.852793e-25, -6.372354e-25, 2.745014e-25, -6.862535e-25, 
    2.058761e-25, -9.803622e-27, -1.372507e-25, 2.450906e-25, -3.725376e-25, 
    -6.666463e-25, -2.548942e-25, 5.686101e-25, 6.127264e-25, -7.156644e-25, 
    -4.019485e-25, -3.62734e-25, 1.470543e-25, -9.313441e-26, 4.65672e-25, 
    -2.352869e-25, -1.715634e-25, 5.882173e-26, -2.695996e-25, 4.215557e-25, 
    -1.960724e-25, -6.862535e-26, -1.56858e-25, 4.901811e-25, 4.41163e-26, 
    1.862688e-25, 5.391992e-25, 1.715634e-25, -6.323336e-25, -2.941087e-25, 
    4.509666e-25, 2.941087e-25, -7.548789e-25, 1.862688e-25, 5.686101e-25, 
    1.068595e-24, -7.352717e-25, 1.068595e-24, 9.803622e-26, -9.705585e-25, 
    -5.293956e-25, 1.911706e-25, 3.921449e-26, -1.176435e-24, 1.56858e-25, 
    -5.490028e-25, 6.862535e-25, -5.588064e-25, 1.176435e-25, 8.333079e-26, 
    3.137159e-25, 1.715634e-25, 4.41163e-25, 1.617598e-25, 5.048866e-25, 
    3.62734e-25, 5.686101e-25, 5.882173e-25, -1.960724e-26,
  9.436746e-32, 9.436709e-32, 9.436716e-32, 9.436686e-32, 9.436703e-32, 
    9.436684e-32, 9.436739e-32, 9.436708e-32, 9.436728e-32, 9.436743e-32, 
    9.436628e-32, 9.436685e-32, 9.436569e-32, 9.436606e-32, 9.436515e-32, 
    9.436575e-32, 9.436503e-32, 9.436517e-32, 9.436475e-32, 9.436487e-32, 
    9.436434e-32, 9.43647e-32, 9.436406e-32, 9.436442e-32, 9.436437e-32, 
    9.436471e-32, 9.436674e-32, 9.436635e-32, 9.436676e-32, 9.436671e-32, 
    9.436673e-32, 9.436703e-32, 9.436718e-32, 9.436749e-32, 9.436743e-32, 
    9.436721e-32, 9.436668e-32, 9.436686e-32, 9.436641e-32, 9.436642e-32, 
    9.436592e-32, 9.436615e-32, 9.436531e-32, 9.436555e-32, 9.436487e-32, 
    9.436504e-32, 9.436487e-32, 9.436492e-32, 9.436487e-32, 9.436512e-32, 
    9.436501e-32, 9.436524e-32, 9.436611e-32, 9.436585e-32, 9.436661e-32, 
    9.436707e-32, 9.436738e-32, 9.436759e-32, 9.436756e-32, 9.436751e-32, 
    9.436721e-32, 9.436692e-32, 9.436671e-32, 9.436656e-32, 9.436642e-32, 
    9.436599e-32, 9.436577e-32, 9.436527e-32, 9.436535e-32, 9.43652e-32, 
    9.436505e-32, 9.436481e-32, 9.436485e-32, 9.436474e-32, 9.436521e-32, 
    9.43649e-32, 9.436541e-32, 9.436527e-32, 9.436638e-32, 9.436681e-32, 
    9.436699e-32, 9.436715e-32, 9.436754e-32, 9.436727e-32, 9.436738e-32, 
    9.436712e-32, 9.436696e-32, 9.436705e-32, 9.436656e-32, 9.436675e-32, 
    9.436575e-32, 9.436618e-32, 9.436507e-32, 9.436534e-32, 9.436501e-32, 
    9.436518e-32, 9.436489e-32, 9.436515e-32, 9.43647e-32, 9.43646e-32, 
    9.436467e-32, 9.436441e-32, 9.436516e-32, 9.436487e-32, 9.436705e-32, 
    9.436703e-32, 9.436698e-32, 9.436724e-32, 9.436725e-32, 9.436749e-32, 
    9.436728e-32, 9.436719e-32, 9.436696e-32, 9.436682e-32, 9.436669e-32, 
    9.436641e-32, 9.436608e-32, 9.436564e-32, 9.436532e-32, 9.436511e-32, 
    9.436524e-32, 9.436512e-32, 9.436525e-32, 9.436531e-32, 9.436464e-32, 
    9.436501e-32, 9.436445e-32, 9.436448e-32, 9.436474e-32, 9.436447e-32, 
    9.436702e-32, 9.43671e-32, 9.436736e-32, 9.436715e-32, 9.436752e-32, 
    9.436732e-32, 9.43672e-32, 9.436675e-32, 9.436665e-32, 9.436655e-32, 
    9.436637e-32, 9.436614e-32, 9.436572e-32, 9.436537e-32, 9.436504e-32, 
    9.436507e-32, 9.436506e-32, 9.436499e-32, 9.436517e-32, 9.436496e-32, 
    9.436492e-32, 9.436501e-32, 9.436448e-32, 9.436464e-32, 9.436448e-32, 
    9.436458e-32, 9.436708e-32, 9.436695e-32, 9.436702e-32, 9.436689e-32, 
    9.436698e-32, 9.436659e-32, 9.436646e-32, 9.436591e-32, 9.436614e-32, 
    9.436578e-32, 9.436611e-32, 9.436605e-32, 9.436577e-32, 9.436609e-32, 
    9.436539e-32, 9.436586e-32, 9.436498e-32, 9.436545e-32, 9.436495e-32, 
    9.436505e-32, 9.43649e-32, 9.436476e-32, 9.436459e-32, 9.436428e-32, 
    9.436435e-32, 9.436409e-32, 9.436676e-32, 9.436661e-32, 9.436662e-32, 
    9.436645e-32, 9.436632e-32, 9.436606e-32, 9.436562e-32, 9.436579e-32, 
    9.436549e-32, 9.436543e-32, 9.436588e-32, 9.43656e-32, 9.43665e-32, 
    9.436635e-32, 9.436644e-32, 9.436675e-32, 9.436575e-32, 9.436626e-32, 
    9.436531e-32, 9.436559e-32, 9.436478e-32, 9.436518e-32, 9.436439e-32, 
    9.436406e-32, 9.436374e-32, 9.436337e-32, 9.436652e-32, 9.436663e-32, 
    9.436643e-32, 9.436616e-32, 9.436591e-32, 9.436558e-32, 9.436554e-32, 
    9.436548e-32, 9.436532e-32, 9.436518e-32, 9.436546e-32, 9.436515e-32, 
    9.436632e-32, 9.436571e-32, 9.436667e-32, 9.436638e-32, 9.436618e-32, 
    9.436626e-32, 9.436581e-32, 9.436569e-32, 9.436526e-32, 9.436548e-32, 
    9.436414e-32, 9.436473e-32, 9.436309e-32, 9.436354e-32, 9.436666e-32, 
    9.436652e-32, 9.436601e-32, 9.436625e-32, 9.436555e-32, 9.436538e-32, 
    9.436524e-32, 9.436507e-32, 9.436505e-32, 9.436494e-32, 9.436511e-32, 
    9.436495e-32, 9.436558e-32, 9.43653e-32, 9.436607e-32, 9.436588e-32, 
    9.436597e-32, 9.436606e-32, 9.436577e-32, 9.436545e-32, 9.436545e-32, 
    9.436535e-32, 9.436507e-32, 9.436555e-32, 9.436406e-32, 9.436498e-32, 
    9.436636e-32, 9.436607e-32, 9.436604e-32, 9.436614e-32, 9.43654e-32, 
    9.436567e-32, 9.436494e-32, 9.436514e-32, 9.436482e-32, 9.436498e-32, 
    9.4365e-32, 9.436521e-32, 9.436534e-32, 9.436565e-32, 9.436592e-32, 
    9.436613e-32, 9.436608e-32, 9.436585e-32, 9.436544e-32, 9.436504e-32, 
    9.436513e-32, 9.436484e-32, 9.43656e-32, 9.436528e-32, 9.436541e-32, 
    9.436508e-32, 9.436579e-32, 9.436519e-32, 9.436594e-32, 9.436588e-32, 
    9.436567e-32, 9.436526e-32, 9.436517e-32, 9.436508e-32, 9.436514e-32, 
    9.436542e-32, 9.436547e-32, 9.436568e-32, 9.436574e-32, 9.436589e-32, 
    9.436602e-32, 9.436591e-32, 9.436578e-32, 9.436542e-32, 9.436511e-32, 
    9.436476e-32, 9.436467e-32, 9.436427e-32, 9.43646e-32, 9.436406e-32, 
    9.436452e-32, 9.436372e-32, 9.436515e-32, 9.436453e-32, 9.436567e-32, 
    9.436554e-32, 9.436532e-32, 9.436481e-32, 9.436509e-32, 9.436477e-32, 
    9.436548e-32, 9.436584e-32, 9.436594e-32, 9.436611e-32, 9.436593e-32, 
    9.436595e-32, 9.436577e-32, 9.436583e-32, 9.436541e-32, 9.436564e-32, 
    9.4365e-32, 9.436477e-32, 9.436412e-32, 9.436372e-32, 9.436331e-32, 
    9.436313e-32, 9.436308e-32, 9.436306e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.030664e-14, 4.041577e-14, 4.039457e-14, 4.048251e-14, 4.043375e-14, 
    4.049131e-14, 4.032879e-14, 4.042009e-14, 4.036182e-14, 4.031649e-14, 
    4.065291e-14, 4.048644e-14, 4.082571e-14, 4.071972e-14, 4.098579e-14, 
    4.08092e-14, 4.102137e-14, 4.098074e-14, 4.110308e-14, 4.106805e-14, 
    4.122429e-14, 4.111924e-14, 4.130525e-14, 4.119924e-14, 4.121581e-14, 
    4.111577e-14, 4.052e-14, 4.063219e-14, 4.051334e-14, 4.052934e-14, 
    4.052217e-14, 4.043475e-14, 4.039064e-14, 4.029832e-14, 4.031509e-14, 
    4.038291e-14, 4.053654e-14, 4.048444e-14, 4.061578e-14, 4.061281e-14, 
    4.075881e-14, 4.069301e-14, 4.09381e-14, 4.086852e-14, 4.106951e-14, 
    4.101899e-14, 4.106714e-14, 4.105254e-14, 4.106733e-14, 4.099322e-14, 
    4.102497e-14, 4.095976e-14, 4.070533e-14, 4.078016e-14, 4.055679e-14, 
    4.042219e-14, 4.033279e-14, 4.026927e-14, 4.027826e-14, 4.029537e-14, 
    4.038331e-14, 4.046595e-14, 4.052888e-14, 4.057095e-14, 4.061239e-14, 
    4.073762e-14, 4.080392e-14, 4.095214e-14, 4.092544e-14, 4.09707e-14, 
    4.101397e-14, 4.108652e-14, 4.107459e-14, 4.110653e-14, 4.096953e-14, 
    4.106059e-14, 4.091024e-14, 4.095136e-14, 4.062352e-14, 4.049851e-14, 
    4.044522e-14, 4.039864e-14, 4.028516e-14, 4.036354e-14, 4.033264e-14, 
    4.040615e-14, 4.045281e-14, 4.042974e-14, 4.05721e-14, 4.051677e-14, 
    4.080785e-14, 4.068258e-14, 4.100892e-14, 4.093092e-14, 4.102761e-14, 
    4.097829e-14, 4.106277e-14, 4.098674e-14, 4.111843e-14, 4.114707e-14, 
    4.11275e-14, 4.12027e-14, 4.098252e-14, 4.106712e-14, 4.042909e-14, 
    4.043285e-14, 4.045039e-14, 4.037326e-14, 4.036855e-14, 4.029785e-14, 
    4.036077e-14, 4.038754e-14, 4.045553e-14, 4.04957e-14, 4.053387e-14, 
    4.061777e-14, 4.071136e-14, 4.084213e-14, 4.093598e-14, 4.099885e-14, 
    4.096031e-14, 4.099433e-14, 4.095629e-14, 4.093846e-14, 4.113633e-14, 
    4.102526e-14, 4.119189e-14, 4.118268e-14, 4.110729e-14, 4.118372e-14, 
    4.04355e-14, 4.041384e-14, 4.033858e-14, 4.039748e-14, 4.029015e-14, 
    4.035023e-14, 4.038475e-14, 4.05179e-14, 4.054717e-14, 4.057425e-14, 
    4.062776e-14, 4.069638e-14, 4.081663e-14, 4.092114e-14, 4.101649e-14, 
    4.100951e-14, 4.101196e-14, 4.103324e-14, 4.098051e-14, 4.104189e-14, 
    4.105218e-14, 4.102526e-14, 4.118145e-14, 4.113685e-14, 4.118248e-14, 
    4.115345e-14, 4.042088e-14, 4.045732e-14, 4.043763e-14, 4.047465e-14, 
    4.044856e-14, 4.056448e-14, 4.059921e-14, 4.07616e-14, 4.069502e-14, 
    4.0801e-14, 4.07058e-14, 4.072267e-14, 4.08044e-14, 4.071096e-14, 
    4.091537e-14, 4.077678e-14, 4.103407e-14, 4.08958e-14, 4.104272e-14, 
    4.101608e-14, 4.106021e-14, 4.10997e-14, 4.114939e-14, 4.124096e-14, 
    4.121977e-14, 4.129633e-14, 4.051164e-14, 4.055885e-14, 4.055471e-14, 
    4.060412e-14, 4.064063e-14, 4.071977e-14, 4.084653e-14, 4.079888e-14, 
    4.088636e-14, 4.09039e-14, 4.077102e-14, 4.08526e-14, 4.059045e-14, 
    4.063282e-14, 4.060762e-14, 4.051535e-14, 4.080983e-14, 4.065879e-14, 
    4.093753e-14, 4.085586e-14, 4.109406e-14, 4.097563e-14, 4.12081e-14, 
    4.130724e-14, 4.140058e-14, 4.150941e-14, 4.058463e-14, 4.055256e-14, 
    4.061e-14, 4.068937e-14, 4.076303e-14, 4.086084e-14, 4.087085e-14, 
    4.088916e-14, 4.093656e-14, 4.097641e-14, 4.089492e-14, 4.09864e-14, 
    4.06426e-14, 4.082294e-14, 4.054041e-14, 4.062554e-14, 4.068471e-14, 
    4.065878e-14, 4.079345e-14, 4.082515e-14, 4.095386e-14, 4.088737e-14, 
    4.128276e-14, 4.1108e-14, 4.159227e-14, 4.145716e-14, 4.054134e-14, 
    4.058453e-14, 4.073466e-14, 4.066326e-14, 4.086738e-14, 4.091755e-14, 
    4.095831e-14, 4.101039e-14, 4.101603e-14, 4.104687e-14, 4.099632e-14, 
    4.104489e-14, 4.086105e-14, 4.094323e-14, 4.071754e-14, 4.077251e-14, 
    4.074723e-14, 4.071948e-14, 4.08051e-14, 4.08962e-14, 4.089818e-14, 
    4.092735e-14, 4.100948e-14, 4.08682e-14, 4.130522e-14, 4.103547e-14, 
    4.06316e-14, 4.071464e-14, 4.072655e-14, 4.069438e-14, 4.091252e-14, 
    4.083353e-14, 4.104613e-14, 4.098871e-14, 4.108278e-14, 4.103604e-14, 
    4.102916e-14, 4.096911e-14, 4.09317e-14, 4.083714e-14, 4.076014e-14, 
    4.069905e-14, 4.071326e-14, 4.078035e-14, 4.090178e-14, 4.101652e-14, 
    4.099139e-14, 4.107563e-14, 4.085259e-14, 4.094614e-14, 4.090999e-14, 
    4.100426e-14, 4.079761e-14, 4.097349e-14, 4.075258e-14, 4.077198e-14, 
    4.083196e-14, 4.095246e-14, 4.097916e-14, 4.10076e-14, 4.099006e-14, 
    4.090486e-14, 4.089092e-14, 4.083051e-14, 4.081381e-14, 4.076776e-14, 
    4.072961e-14, 4.076446e-14, 4.080104e-14, 4.090492e-14, 4.09984e-14, 
    4.110025e-14, 4.112518e-14, 4.124393e-14, 4.114722e-14, 4.130671e-14, 
    4.117105e-14, 4.140581e-14, 4.098373e-14, 4.116714e-14, 4.08347e-14, 
    4.087058e-14, 4.093537e-14, 4.108397e-14, 4.100382e-14, 4.109757e-14, 
    4.089037e-14, 4.078265e-14, 4.07548e-14, 4.070276e-14, 4.075599e-14, 
    4.075167e-14, 4.080258e-14, 4.078623e-14, 4.090836e-14, 4.084278e-14, 
    4.102898e-14, 4.109684e-14, 4.128829e-14, 4.140545e-14, 4.152462e-14, 
    4.157717e-14, 4.159316e-14, 4.159984e-14 ;

 LITR1N_vr =
  5.55759e-05, 5.557569e-05, 5.557573e-05, 5.557556e-05, 5.557566e-05, 
    5.557554e-05, 5.557586e-05, 5.557568e-05, 5.557579e-05, 5.557589e-05, 
    5.557523e-05, 5.557555e-05, 5.55749e-05, 5.55751e-05, 5.557459e-05, 
    5.557493e-05, 5.557452e-05, 5.55746e-05, 5.557436e-05, 5.557443e-05, 
    5.557412e-05, 5.557433e-05, 5.557397e-05, 5.557417e-05, 5.557414e-05, 
    5.557434e-05, 5.557549e-05, 5.557527e-05, 5.55755e-05, 5.557547e-05, 
    5.557549e-05, 5.557566e-05, 5.557574e-05, 5.557592e-05, 5.557589e-05, 
    5.557575e-05, 5.557546e-05, 5.557556e-05, 5.55753e-05, 5.557531e-05, 
    5.557503e-05, 5.557515e-05, 5.557468e-05, 5.557481e-05, 5.557442e-05, 
    5.557452e-05, 5.557443e-05, 5.557446e-05, 5.557443e-05, 5.557457e-05, 
    5.557451e-05, 5.557464e-05, 5.557513e-05, 5.557498e-05, 5.557542e-05, 
    5.557568e-05, 5.557585e-05, 5.557598e-05, 5.557596e-05, 5.557593e-05, 
    5.557575e-05, 5.557559e-05, 5.557547e-05, 5.557539e-05, 5.557531e-05, 
    5.557507e-05, 5.557494e-05, 5.557465e-05, 5.55747e-05, 5.557462e-05, 
    5.557453e-05, 5.557439e-05, 5.557442e-05, 5.557435e-05, 5.557462e-05, 
    5.557444e-05, 5.557473e-05, 5.557465e-05, 5.557529e-05, 5.557553e-05, 
    5.557563e-05, 5.557573e-05, 5.557594e-05, 5.557579e-05, 5.557585e-05, 
    5.557571e-05, 5.557562e-05, 5.557566e-05, 5.557539e-05, 5.55755e-05, 
    5.557493e-05, 5.557517e-05, 5.557454e-05, 5.557469e-05, 5.557451e-05, 
    5.55746e-05, 5.557444e-05, 5.557458e-05, 5.557433e-05, 5.557427e-05, 
    5.557431e-05, 5.557416e-05, 5.557459e-05, 5.557443e-05, 5.557567e-05, 
    5.557566e-05, 5.557562e-05, 5.557577e-05, 5.557578e-05, 5.557592e-05, 
    5.55758e-05, 5.557575e-05, 5.557561e-05, 5.557554e-05, 5.557546e-05, 
    5.55753e-05, 5.557512e-05, 5.557486e-05, 5.557468e-05, 5.557456e-05, 
    5.557464e-05, 5.557457e-05, 5.557464e-05, 5.557468e-05, 5.55743e-05, 
    5.557451e-05, 5.557419e-05, 5.55742e-05, 5.557435e-05, 5.55742e-05, 
    5.557565e-05, 5.55757e-05, 5.557584e-05, 5.557573e-05, 5.557594e-05, 
    5.557582e-05, 5.557575e-05, 5.557549e-05, 5.557544e-05, 5.557538e-05, 
    5.557528e-05, 5.557515e-05, 5.557491e-05, 5.557471e-05, 5.557453e-05, 
    5.557454e-05, 5.557454e-05, 5.55745e-05, 5.55746e-05, 5.557448e-05, 
    5.557446e-05, 5.557451e-05, 5.557421e-05, 5.55743e-05, 5.55742e-05, 
    5.557426e-05, 5.557568e-05, 5.557561e-05, 5.557565e-05, 5.557558e-05, 
    5.557563e-05, 5.55754e-05, 5.557534e-05, 5.557502e-05, 5.557515e-05, 
    5.557494e-05, 5.557513e-05, 5.55751e-05, 5.557494e-05, 5.557512e-05, 
    5.557472e-05, 5.557499e-05, 5.557449e-05, 5.557476e-05, 5.557448e-05, 
    5.557453e-05, 5.557444e-05, 5.557436e-05, 5.557427e-05, 5.557409e-05, 
    5.557413e-05, 5.557399e-05, 5.557551e-05, 5.557541e-05, 5.557542e-05, 
    5.557532e-05, 5.557526e-05, 5.55751e-05, 5.557486e-05, 5.557495e-05, 
    5.557478e-05, 5.557475e-05, 5.5575e-05, 5.557484e-05, 5.557535e-05, 
    5.557527e-05, 5.557532e-05, 5.55755e-05, 5.557493e-05, 5.557522e-05, 
    5.557468e-05, 5.557484e-05, 5.557438e-05, 5.55746e-05, 5.557416e-05, 
    5.557396e-05, 5.557378e-05, 5.557357e-05, 5.557536e-05, 5.557543e-05, 
    5.557531e-05, 5.557516e-05, 5.557502e-05, 5.557483e-05, 5.557481e-05, 
    5.557477e-05, 5.557468e-05, 5.55746e-05, 5.557476e-05, 5.557459e-05, 
    5.557525e-05, 5.55749e-05, 5.557545e-05, 5.557528e-05, 5.557517e-05, 
    5.557522e-05, 5.557496e-05, 5.55749e-05, 5.557465e-05, 5.557478e-05, 
    5.557401e-05, 5.557435e-05, 5.557341e-05, 5.557367e-05, 5.557545e-05, 
    5.557536e-05, 5.557507e-05, 5.557521e-05, 5.557482e-05, 5.557472e-05, 
    5.557464e-05, 5.557454e-05, 5.557453e-05, 5.557447e-05, 5.557456e-05, 
    5.557447e-05, 5.557483e-05, 5.557467e-05, 5.557511e-05, 5.5575e-05, 
    5.557505e-05, 5.55751e-05, 5.557494e-05, 5.557476e-05, 5.557476e-05, 
    5.55747e-05, 5.557454e-05, 5.557482e-05, 5.557397e-05, 5.557449e-05, 
    5.557527e-05, 5.557511e-05, 5.557509e-05, 5.557515e-05, 5.557473e-05, 
    5.557488e-05, 5.557447e-05, 5.557458e-05, 5.55744e-05, 5.557449e-05, 
    5.55745e-05, 5.557462e-05, 5.557469e-05, 5.557487e-05, 5.557502e-05, 
    5.557514e-05, 5.557511e-05, 5.557498e-05, 5.557475e-05, 5.557453e-05, 
    5.557458e-05, 5.557441e-05, 5.557484e-05, 5.557466e-05, 5.557473e-05, 
    5.557455e-05, 5.557495e-05, 5.557461e-05, 5.557504e-05, 5.5575e-05, 
    5.557488e-05, 5.557465e-05, 5.55746e-05, 5.557454e-05, 5.557458e-05, 
    5.557474e-05, 5.557477e-05, 5.557489e-05, 5.557492e-05, 5.557501e-05, 
    5.557508e-05, 5.557502e-05, 5.557494e-05, 5.557474e-05, 5.557456e-05, 
    5.557436e-05, 5.557432e-05, 5.557408e-05, 5.557427e-05, 5.557396e-05, 
    5.557423e-05, 5.557377e-05, 5.557459e-05, 5.557423e-05, 5.557488e-05, 
    5.557481e-05, 5.557468e-05, 5.55744e-05, 5.557455e-05, 5.557437e-05, 
    5.557477e-05, 5.557498e-05, 5.557503e-05, 5.557514e-05, 5.557503e-05, 
    5.557504e-05, 5.557494e-05, 5.557497e-05, 5.557474e-05, 5.557486e-05, 
    5.55745e-05, 5.557437e-05, 5.5574e-05, 5.557377e-05, 5.557354e-05, 
    5.557344e-05, 5.557341e-05, 5.55734e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  6.985294e-13, 7.004207e-13, 7.000534e-13, 7.015774e-13, 7.007323e-13, 
    7.017299e-13, 6.989133e-13, 7.004955e-13, 6.994858e-13, 6.987002e-13, 
    7.045305e-13, 7.016454e-13, 7.075251e-13, 7.056883e-13, 7.102994e-13, 
    7.07239e-13, 7.10916e-13, 7.102118e-13, 7.12332e-13, 7.117249e-13, 
    7.144326e-13, 7.126122e-13, 7.158357e-13, 7.139984e-13, 7.142857e-13, 
    7.12552e-13, 7.02227e-13, 7.041713e-13, 7.021115e-13, 7.02389e-13, 
    7.022647e-13, 7.007496e-13, 6.999852e-13, 6.983853e-13, 6.986759e-13, 
    6.998512e-13, 7.025138e-13, 7.016108e-13, 7.038869e-13, 7.038355e-13, 
    7.063657e-13, 7.052254e-13, 7.094728e-13, 7.08267e-13, 7.117503e-13, 
    7.108748e-13, 7.117091e-13, 7.114562e-13, 7.117124e-13, 7.104281e-13, 
    7.109785e-13, 7.098482e-13, 7.054389e-13, 7.067358e-13, 7.028646e-13, 
    7.00532e-13, 6.989826e-13, 6.978819e-13, 6.980375e-13, 6.983341e-13, 
    6.998581e-13, 7.012904e-13, 7.02381e-13, 7.0311e-13, 7.038282e-13, 
    7.059985e-13, 7.071475e-13, 7.097162e-13, 7.092535e-13, 7.100378e-13, 
    7.107877e-13, 7.120451e-13, 7.118382e-13, 7.123919e-13, 7.100175e-13, 
    7.115957e-13, 7.0899e-13, 7.097028e-13, 7.040212e-13, 7.018545e-13, 
    7.00931e-13, 7.001239e-13, 6.981572e-13, 6.995154e-13, 6.9898e-13, 
    7.00254e-13, 7.010627e-13, 7.006628e-13, 7.031299e-13, 7.021711e-13, 
    7.072156e-13, 7.050445e-13, 7.107002e-13, 7.093485e-13, 7.110242e-13, 
    7.101694e-13, 7.116335e-13, 7.103159e-13, 7.125981e-13, 7.130944e-13, 
    7.127552e-13, 7.140585e-13, 7.102427e-13, 7.117088e-13, 7.006515e-13, 
    7.007167e-13, 7.010207e-13, 6.99684e-13, 6.996024e-13, 6.983772e-13, 
    6.994676e-13, 6.999315e-13, 7.011097e-13, 7.018059e-13, 7.024675e-13, 
    7.039215e-13, 7.055434e-13, 7.078097e-13, 7.094361e-13, 7.105256e-13, 
    7.098578e-13, 7.104474e-13, 7.097882e-13, 7.094792e-13, 7.129083e-13, 
    7.109835e-13, 7.138711e-13, 7.137115e-13, 7.12405e-13, 7.137295e-13, 
    7.007625e-13, 7.003872e-13, 6.990829e-13, 7.001038e-13, 6.982437e-13, 
    6.992848e-13, 6.99883e-13, 7.021907e-13, 7.026978e-13, 7.031673e-13, 
    7.040946e-13, 7.052838e-13, 7.073677e-13, 7.091789e-13, 7.108314e-13, 
    7.107104e-13, 7.10753e-13, 7.111217e-13, 7.102079e-13, 7.112717e-13, 
    7.114499e-13, 7.109835e-13, 7.136902e-13, 7.129174e-13, 7.137082e-13, 
    7.13205e-13, 7.005093e-13, 7.011408e-13, 7.007996e-13, 7.014411e-13, 
    7.00989e-13, 7.029979e-13, 7.035998e-13, 7.064141e-13, 7.052602e-13, 
    7.070969e-13, 7.05447e-13, 7.057394e-13, 7.071559e-13, 7.055364e-13, 
    7.09079e-13, 7.066771e-13, 7.11136e-13, 7.087398e-13, 7.112861e-13, 
    7.108242e-13, 7.11589e-13, 7.122734e-13, 7.131345e-13, 7.147216e-13, 
    7.143543e-13, 7.15681e-13, 7.020821e-13, 7.029003e-13, 7.028287e-13, 
    7.036849e-13, 7.043177e-13, 7.056891e-13, 7.078859e-13, 7.070602e-13, 
    7.085762e-13, 7.088802e-13, 7.065773e-13, 7.079912e-13, 7.03448e-13, 
    7.041824e-13, 7.037454e-13, 7.021464e-13, 7.0725e-13, 7.046324e-13, 
    7.094629e-13, 7.080476e-13, 7.121758e-13, 7.101234e-13, 7.14152e-13, 
    7.158702e-13, 7.174878e-13, 7.193738e-13, 7.033472e-13, 7.027913e-13, 
    7.037867e-13, 7.051623e-13, 7.064389e-13, 7.081339e-13, 7.083075e-13, 
    7.086247e-13, 7.094462e-13, 7.101368e-13, 7.087246e-13, 7.103099e-13, 
    7.043518e-13, 7.074772e-13, 7.025807e-13, 7.040561e-13, 7.050815e-13, 
    7.046322e-13, 7.06966e-13, 7.075154e-13, 7.097459e-13, 7.085937e-13, 
    7.154459e-13, 7.124174e-13, 7.208099e-13, 7.184684e-13, 7.02597e-13, 
    7.033454e-13, 7.059472e-13, 7.047098e-13, 7.082472e-13, 7.091167e-13, 
    7.098232e-13, 7.107257e-13, 7.108234e-13, 7.113579e-13, 7.104819e-13, 
    7.113235e-13, 7.081375e-13, 7.095618e-13, 7.056505e-13, 7.066031e-13, 
    7.061651e-13, 7.056842e-13, 7.071679e-13, 7.087467e-13, 7.087811e-13, 
    7.092865e-13, 7.107099e-13, 7.082616e-13, 7.158352e-13, 7.111603e-13, 
    7.041611e-13, 7.056003e-13, 7.058066e-13, 7.052491e-13, 7.090295e-13, 
    7.076606e-13, 7.11345e-13, 7.1035e-13, 7.119802e-13, 7.111702e-13, 
    7.11051e-13, 7.100103e-13, 7.093619e-13, 7.077233e-13, 7.063887e-13, 
    7.053301e-13, 7.055763e-13, 7.06739e-13, 7.088434e-13, 7.108319e-13, 
    7.103964e-13, 7.118564e-13, 7.07991e-13, 7.096122e-13, 7.089858e-13, 
    7.106195e-13, 7.070381e-13, 7.100862e-13, 7.062579e-13, 7.06594e-13, 
    7.076334e-13, 7.097217e-13, 7.101845e-13, 7.106772e-13, 7.103733e-13, 
    7.088969e-13, 7.086551e-13, 7.076083e-13, 7.073189e-13, 7.065209e-13, 
    7.058596e-13, 7.064636e-13, 7.070976e-13, 7.088978e-13, 7.105179e-13, 
    7.122831e-13, 7.12715e-13, 7.147731e-13, 7.13097e-13, 7.15861e-13, 
    7.135099e-13, 7.175784e-13, 7.102637e-13, 7.134422e-13, 7.076809e-13, 
    7.083027e-13, 7.094256e-13, 7.120009e-13, 7.106118e-13, 7.122366e-13, 
    7.086457e-13, 7.067788e-13, 7.062963e-13, 7.053943e-13, 7.063169e-13, 
    7.062419e-13, 7.071243e-13, 7.068408e-13, 7.089576e-13, 7.078209e-13, 
    7.110479e-13, 7.122239e-13, 7.155418e-13, 7.175722e-13, 7.196376e-13, 
    7.205482e-13, 7.208253e-13, 7.209411e-13 ;

 LITR2C =
  1.939601e-05, 1.939599e-05, 1.939599e-05, 1.939597e-05, 1.939598e-05, 
    1.939597e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 1.9396e-05, 
    1.939594e-05, 1.939597e-05, 1.939591e-05, 1.939593e-05, 1.939588e-05, 
    1.939592e-05, 1.939588e-05, 1.939589e-05, 1.939586e-05, 1.939587e-05, 
    1.939584e-05, 1.939586e-05, 1.939583e-05, 1.939585e-05, 1.939584e-05, 
    1.939586e-05, 1.939597e-05, 1.939595e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939598e-05, 1.939599e-05, 1.939601e-05, 1.9396e-05, 
    1.939599e-05, 1.939596e-05, 1.939597e-05, 1.939595e-05, 1.939595e-05, 
    1.939593e-05, 1.939594e-05, 1.939589e-05, 1.939591e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939588e-05, 
    1.939588e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 1.939596e-05, 
    1.939599e-05, 1.9396e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 
    1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 
    1.939593e-05, 1.939592e-05, 1.939589e-05, 1.939589e-05, 1.939589e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939586e-05, 1.939589e-05, 
    1.939587e-05, 1.93959e-05, 1.939589e-05, 1.939595e-05, 1.939597e-05, 
    1.939598e-05, 1.939599e-05, 1.939601e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 
    1.939592e-05, 1.939594e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 1.939585e-05, 
    1.939586e-05, 1.939585e-05, 1.939589e-05, 1.939587e-05, 1.939598e-05, 
    1.939598e-05, 1.939598e-05, 1.939599e-05, 1.939599e-05, 1.939601e-05, 
    1.9396e-05, 1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939597e-05, 
    1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939588e-05, 1.939589e-05, 1.939589e-05, 1.939586e-05, 
    1.939588e-05, 1.939585e-05, 1.939585e-05, 1.939586e-05, 1.939585e-05, 
    1.939598e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 1.939601e-05, 
    1.9396e-05, 1.939599e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939594e-05, 1.939591e-05, 1.93959e-05, 1.939588e-05, 
    1.939588e-05, 1.939588e-05, 1.939588e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939585e-05, 1.939586e-05, 1.939585e-05, 
    1.939585e-05, 1.939599e-05, 1.939598e-05, 1.939598e-05, 1.939597e-05, 
    1.939598e-05, 1.939596e-05, 1.939595e-05, 1.939592e-05, 1.939594e-05, 
    1.939592e-05, 1.939593e-05, 1.939593e-05, 1.939592e-05, 1.939593e-05, 
    1.93959e-05, 1.939592e-05, 1.939587e-05, 1.93959e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939586e-05, 1.939585e-05, 1.939584e-05, 
    1.939584e-05, 1.939583e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939592e-05, 
    1.93959e-05, 1.93959e-05, 1.939592e-05, 1.939591e-05, 1.939595e-05, 
    1.939595e-05, 1.939595e-05, 1.939597e-05, 1.939592e-05, 1.939594e-05, 
    1.939589e-05, 1.939591e-05, 1.939587e-05, 1.939589e-05, 1.939584e-05, 
    1.939583e-05, 1.939581e-05, 1.939579e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939594e-05, 1.939592e-05, 1.939591e-05, 1.939591e-05, 
    1.93959e-05, 1.939589e-05, 1.939589e-05, 1.93959e-05, 1.939588e-05, 
    1.939595e-05, 1.939591e-05, 1.939596e-05, 1.939595e-05, 1.939594e-05, 
    1.939594e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939583e-05, 1.939586e-05, 1.939578e-05, 1.93958e-05, 1.939596e-05, 
    1.939596e-05, 1.939593e-05, 1.939594e-05, 1.939591e-05, 1.93959e-05, 
    1.939589e-05, 1.939588e-05, 1.939588e-05, 1.939587e-05, 1.939588e-05, 
    1.939587e-05, 1.939591e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.93959e-05, 
    1.939589e-05, 1.939588e-05, 1.939591e-05, 1.939583e-05, 1.939587e-05, 
    1.939595e-05, 1.939593e-05, 1.939593e-05, 1.939594e-05, 1.93959e-05, 
    1.939591e-05, 1.939587e-05, 1.939588e-05, 1.939587e-05, 1.939587e-05, 
    1.939588e-05, 1.939589e-05, 1.939589e-05, 1.939591e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.939588e-05, 
    1.939588e-05, 1.939587e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939588e-05, 1.939592e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 
    1.939591e-05, 1.939589e-05, 1.939589e-05, 1.939588e-05, 1.939588e-05, 
    1.93959e-05, 1.93959e-05, 1.939591e-05, 1.939591e-05, 1.939592e-05, 
    1.939593e-05, 1.939592e-05, 1.939592e-05, 1.93959e-05, 1.939588e-05, 
    1.939586e-05, 1.939586e-05, 1.939584e-05, 1.939585e-05, 1.939583e-05, 
    1.939585e-05, 1.939581e-05, 1.939588e-05, 1.939585e-05, 1.939591e-05, 
    1.939591e-05, 1.939589e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 
    1.93959e-05, 1.939592e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 
    1.939593e-05, 1.939592e-05, 1.939592e-05, 1.93959e-05, 1.939591e-05, 
    1.939588e-05, 1.939586e-05, 1.939583e-05, 1.939581e-05, 1.939579e-05, 
    1.939578e-05, 1.939578e-05, 1.939577e-05 ;

 LITR2C_TO_SOIL1C =
  1.063689e-13, 1.066571e-13, 1.066011e-13, 1.068334e-13, 1.067046e-13, 
    1.068567e-13, 1.064274e-13, 1.066685e-13, 1.065146e-13, 1.063949e-13, 
    1.072836e-13, 1.068438e-13, 1.0774e-13, 1.074601e-13, 1.081629e-13, 
    1.076964e-13, 1.082569e-13, 1.081496e-13, 1.084727e-13, 1.083802e-13, 
    1.087929e-13, 1.085154e-13, 1.090068e-13, 1.087267e-13, 1.087705e-13, 
    1.085063e-13, 1.069325e-13, 1.072288e-13, 1.069149e-13, 1.069572e-13, 
    1.069382e-13, 1.067073e-13, 1.065908e-13, 1.063469e-13, 1.063912e-13, 
    1.065703e-13, 1.069762e-13, 1.068385e-13, 1.071855e-13, 1.071776e-13, 
    1.075633e-13, 1.073895e-13, 1.080369e-13, 1.078531e-13, 1.083841e-13, 
    1.082506e-13, 1.083778e-13, 1.083392e-13, 1.083783e-13, 1.081825e-13, 
    1.082664e-13, 1.080941e-13, 1.07422e-13, 1.076197e-13, 1.070297e-13, 
    1.066741e-13, 1.064379e-13, 1.062702e-13, 1.062939e-13, 1.063391e-13, 
    1.065714e-13, 1.067897e-13, 1.069559e-13, 1.070671e-13, 1.071765e-13, 
    1.075073e-13, 1.076825e-13, 1.08074e-13, 1.080035e-13, 1.08123e-13, 
    1.082373e-13, 1.08429e-13, 1.083975e-13, 1.084819e-13, 1.081199e-13, 
    1.083605e-13, 1.079633e-13, 1.08072e-13, 1.072059e-13, 1.068757e-13, 
    1.067349e-13, 1.066119e-13, 1.063121e-13, 1.065192e-13, 1.064376e-13, 
    1.066317e-13, 1.06755e-13, 1.06694e-13, 1.070701e-13, 1.069239e-13, 
    1.076929e-13, 1.073619e-13, 1.08224e-13, 1.08018e-13, 1.082734e-13, 
    1.081431e-13, 1.083663e-13, 1.081654e-13, 1.085133e-13, 1.085889e-13, 
    1.085372e-13, 1.087359e-13, 1.081543e-13, 1.083777e-13, 1.066923e-13, 
    1.067023e-13, 1.067486e-13, 1.065449e-13, 1.065324e-13, 1.063457e-13, 
    1.065119e-13, 1.065826e-13, 1.067622e-13, 1.068683e-13, 1.069691e-13, 
    1.071907e-13, 1.07438e-13, 1.077834e-13, 1.080313e-13, 1.081974e-13, 
    1.080956e-13, 1.081855e-13, 1.08085e-13, 1.080379e-13, 1.085606e-13, 
    1.082672e-13, 1.087073e-13, 1.08683e-13, 1.084839e-13, 1.086858e-13, 
    1.067092e-13, 1.06652e-13, 1.064532e-13, 1.066088e-13, 1.063253e-13, 
    1.06484e-13, 1.065752e-13, 1.069269e-13, 1.070042e-13, 1.070758e-13, 
    1.072171e-13, 1.073984e-13, 1.07716e-13, 1.079921e-13, 1.08244e-13, 
    1.082255e-13, 1.08232e-13, 1.082882e-13, 1.081489e-13, 1.083111e-13, 
    1.083383e-13, 1.082672e-13, 1.086797e-13, 1.085619e-13, 1.086825e-13, 
    1.086058e-13, 1.066706e-13, 1.067669e-13, 1.067149e-13, 1.068127e-13, 
    1.067438e-13, 1.0705e-13, 1.071417e-13, 1.075707e-13, 1.073948e-13, 
    1.076748e-13, 1.074233e-13, 1.074678e-13, 1.076837e-13, 1.074369e-13, 
    1.079769e-13, 1.076108e-13, 1.082904e-13, 1.079252e-13, 1.083133e-13, 
    1.082429e-13, 1.083595e-13, 1.084638e-13, 1.085951e-13, 1.08837e-13, 
    1.08781e-13, 1.089832e-13, 1.069104e-13, 1.070351e-13, 1.070242e-13, 
    1.071547e-13, 1.072511e-13, 1.074602e-13, 1.07795e-13, 1.076692e-13, 
    1.079002e-13, 1.079466e-13, 1.075955e-13, 1.078111e-13, 1.071186e-13, 
    1.072305e-13, 1.071639e-13, 1.069202e-13, 1.076981e-13, 1.072991e-13, 
    1.080354e-13, 1.078197e-13, 1.084489e-13, 1.081361e-13, 1.087501e-13, 
    1.090121e-13, 1.092586e-13, 1.095461e-13, 1.071032e-13, 1.070185e-13, 
    1.071702e-13, 1.073799e-13, 1.075745e-13, 1.078328e-13, 1.078593e-13, 
    1.079076e-13, 1.080329e-13, 1.081381e-13, 1.079229e-13, 1.081645e-13, 
    1.072563e-13, 1.077327e-13, 1.069864e-13, 1.072113e-13, 1.073676e-13, 
    1.072991e-13, 1.076548e-13, 1.077385e-13, 1.080785e-13, 1.079029e-13, 
    1.089474e-13, 1.084857e-13, 1.09765e-13, 1.094081e-13, 1.069889e-13, 
    1.071029e-13, 1.074995e-13, 1.073109e-13, 1.078501e-13, 1.079826e-13, 
    1.080903e-13, 1.082279e-13, 1.082428e-13, 1.083243e-13, 1.081907e-13, 
    1.08319e-13, 1.078334e-13, 1.080505e-13, 1.074543e-13, 1.075995e-13, 
    1.075327e-13, 1.074594e-13, 1.076856e-13, 1.079262e-13, 1.079315e-13, 
    1.080085e-13, 1.082255e-13, 1.078523e-13, 1.090067e-13, 1.082941e-13, 
    1.072273e-13, 1.074466e-13, 1.074781e-13, 1.073931e-13, 1.079693e-13, 
    1.077607e-13, 1.083223e-13, 1.081706e-13, 1.084191e-13, 1.082956e-13, 
    1.082775e-13, 1.081188e-13, 1.0802e-13, 1.077702e-13, 1.075668e-13, 
    1.074055e-13, 1.07443e-13, 1.076202e-13, 1.07941e-13, 1.082441e-13, 
    1.081777e-13, 1.084002e-13, 1.07811e-13, 1.080582e-13, 1.079627e-13, 
    1.082117e-13, 1.076658e-13, 1.081304e-13, 1.075469e-13, 1.075981e-13, 
    1.077565e-13, 1.080748e-13, 1.081454e-13, 1.082205e-13, 1.081742e-13, 
    1.079491e-13, 1.079123e-13, 1.077527e-13, 1.077086e-13, 1.07587e-13, 
    1.074862e-13, 1.075782e-13, 1.076749e-13, 1.079493e-13, 1.081962e-13, 
    1.084653e-13, 1.085311e-13, 1.088448e-13, 1.085893e-13, 1.090106e-13, 
    1.086523e-13, 1.092724e-13, 1.081575e-13, 1.086419e-13, 1.077638e-13, 
    1.078586e-13, 1.080297e-13, 1.084223e-13, 1.082105e-13, 1.084582e-13, 
    1.079108e-13, 1.076263e-13, 1.075527e-13, 1.074152e-13, 1.075559e-13, 
    1.075444e-13, 1.076789e-13, 1.076357e-13, 1.079584e-13, 1.077851e-13, 
    1.08277e-13, 1.084563e-13, 1.08962e-13, 1.092715e-13, 1.095863e-13, 
    1.097251e-13, 1.097674e-13, 1.09785e-13 ;

 LITR2C_vr =
  0.001107532, 0.001107531, 0.001107531, 0.00110753, 0.001107531, 0.00110753, 
    0.001107532, 0.001107531, 0.001107531, 0.001107532, 0.001107528, 
    0.00110753, 0.001107527, 0.001107528, 0.001107525, 0.001107527, 
    0.001107525, 0.001107525, 0.001107524, 0.001107524, 0.001107523, 
    0.001107524, 0.001107522, 0.001107523, 0.001107523, 0.001107524, 
    0.00110753, 0.001107529, 0.00110753, 0.00110753, 0.00110753, 0.001107531, 
    0.001107531, 0.001107532, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.001107527, 0.001107528, 
    0.001107526, 0.001107526, 0.001107524, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107525, 0.001107525, 
    0.001107528, 0.001107527, 0.001107529, 0.001107531, 0.001107532, 
    0.001107532, 0.001107532, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107527, 
    0.001107525, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107529, 0.00110753, 0.001107531, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.00110753, 
    0.001107531, 0.001107529, 0.00110753, 0.001107527, 0.001107528, 
    0.001107525, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107525, 0.001107524, 0.001107523, 0.001107524, 0.001107523, 
    0.001107525, 0.001107524, 0.001107531, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.00110753, 0.00110753, 0.00110753, 0.001107529, 0.001107528, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107525, 
    0.001107525, 0.001107526, 0.001107523, 0.001107525, 0.001107523, 
    0.001107523, 0.001107524, 0.001107523, 0.001107531, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.00110753, 0.00110753, 0.001107529, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107525, 0.001107525, 
    0.001107525, 0.001107525, 0.001107524, 0.001107524, 0.001107525, 
    0.001107523, 0.001107523, 0.001107523, 0.001107523, 0.001107531, 
    0.00110753, 0.001107531, 0.00110753, 0.001107531, 0.001107529, 
    0.001107529, 0.001107527, 0.001107528, 0.001107527, 0.001107528, 
    0.001107528, 0.001107527, 0.001107528, 0.001107526, 0.001107527, 
    0.001107524, 0.001107526, 0.001107524, 0.001107525, 0.001107524, 
    0.001107524, 0.001107523, 0.001107522, 0.001107523, 0.001107522, 
    0.00110753, 0.001107529, 0.00110753, 0.001107529, 0.001107529, 
    0.001107528, 0.001107526, 0.001107527, 0.001107526, 0.001107526, 
    0.001107527, 0.001107526, 0.001107529, 0.001107529, 0.001107529, 
    0.00110753, 0.001107527, 0.001107528, 0.001107526, 0.001107526, 
    0.001107524, 0.001107525, 0.001107523, 0.001107522, 0.001107521, 
    0.00110752, 0.001107529, 0.00110753, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107526, 
    0.001107525, 0.001107526, 0.001107525, 0.001107529, 0.001107527, 
    0.00110753, 0.001107529, 0.001107528, 0.001107528, 0.001107527, 
    0.001107527, 0.001107525, 0.001107526, 0.001107522, 0.001107524, 
    0.001107519, 0.00110752, 0.00110753, 0.001107529, 0.001107528, 
    0.001107528, 0.001107526, 0.001107526, 0.001107525, 0.001107525, 
    0.001107525, 0.001107524, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107528, 0.001107527, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107526, 0.001107522, 0.001107524, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107526, 0.001107527, 0.001107524, 
    0.001107525, 0.001107524, 0.001107524, 0.001107525, 0.001107525, 
    0.001107526, 0.001107527, 0.001107527, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107526, 0.001107525, 0.001107526, 0.001107525, 0.001107527, 
    0.001107525, 0.001107527, 0.001107527, 0.001107527, 0.001107525, 
    0.001107525, 0.001107525, 0.001107525, 0.001107526, 0.001107526, 
    0.001107527, 0.001107527, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107526, 0.001107525, 0.001107524, 0.001107524, 
    0.001107522, 0.001107523, 0.001107522, 0.001107523, 0.001107521, 
    0.001107525, 0.001107523, 0.001107527, 0.001107526, 0.001107526, 
    0.001107524, 0.001107525, 0.001107524, 0.001107526, 0.001107527, 
    0.001107527, 0.001107528, 0.001107527, 0.001107527, 0.001107527, 
    0.001107527, 0.001107526, 0.001107526, 0.001107525, 0.001107524, 
    0.001107522, 0.001107521, 0.001107519, 0.001107519, 0.001107519, 
    0.001107519,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684264e-07, 2.684262e-07, 2.684262e-07, 2.68426e-07, 2.684261e-07, 
    2.68426e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 2.684264e-07, 
    2.684256e-07, 2.68426e-07, 2.684252e-07, 2.684254e-07, 2.684248e-07, 
    2.684252e-07, 2.684247e-07, 2.684248e-07, 2.684245e-07, 2.684246e-07, 
    2.684242e-07, 2.684245e-07, 2.68424e-07, 2.684243e-07, 2.684242e-07, 
    2.684245e-07, 2.684259e-07, 2.684257e-07, 2.684259e-07, 2.684259e-07, 
    2.684259e-07, 2.684261e-07, 2.684262e-07, 2.684265e-07, 2.684264e-07, 
    2.684263e-07, 2.684259e-07, 2.68426e-07, 2.684257e-07, 2.684257e-07, 
    2.684253e-07, 2.684255e-07, 2.684249e-07, 2.684251e-07, 2.684246e-07, 
    2.684247e-07, 2.684246e-07, 2.684246e-07, 2.684246e-07, 2.684248e-07, 
    2.684247e-07, 2.684248e-07, 2.684255e-07, 2.684253e-07, 2.684259e-07, 
    2.684262e-07, 2.684264e-07, 2.684266e-07, 2.684265e-07, 2.684265e-07, 
    2.684263e-07, 2.684261e-07, 2.684259e-07, 2.684258e-07, 2.684257e-07, 
    2.684254e-07, 2.684252e-07, 2.684249e-07, 2.684249e-07, 2.684248e-07, 
    2.684247e-07, 2.684245e-07, 2.684245e-07, 2.684245e-07, 2.684248e-07, 
    2.684246e-07, 2.68425e-07, 2.684249e-07, 2.684257e-07, 2.68426e-07, 
    2.684261e-07, 2.684262e-07, 2.684265e-07, 2.684263e-07, 2.684264e-07, 
    2.684262e-07, 2.684261e-07, 2.684262e-07, 2.684258e-07, 2.684259e-07, 
    2.684252e-07, 2.684255e-07, 2.684247e-07, 2.684249e-07, 2.684247e-07, 
    2.684248e-07, 2.684246e-07, 2.684248e-07, 2.684245e-07, 2.684244e-07, 
    2.684244e-07, 2.684242e-07, 2.684248e-07, 2.684246e-07, 2.684262e-07, 
    2.684261e-07, 2.684261e-07, 2.684263e-07, 2.684263e-07, 2.684265e-07, 
    2.684263e-07, 2.684262e-07, 2.684261e-07, 2.68426e-07, 2.684259e-07, 
    2.684257e-07, 2.684255e-07, 2.684251e-07, 2.684249e-07, 2.684247e-07, 
    2.684248e-07, 2.684247e-07, 2.684249e-07, 2.684249e-07, 2.684244e-07, 
    2.684247e-07, 2.684243e-07, 2.684243e-07, 2.684245e-07, 2.684243e-07, 
    2.684261e-07, 2.684262e-07, 2.684264e-07, 2.684262e-07, 2.684265e-07, 
    2.684264e-07, 2.684263e-07, 2.684259e-07, 2.684259e-07, 2.684258e-07, 
    2.684257e-07, 2.684255e-07, 2.684252e-07, 2.684249e-07, 2.684247e-07, 
    2.684247e-07, 2.684247e-07, 2.684247e-07, 2.684248e-07, 2.684246e-07, 
    2.684246e-07, 2.684247e-07, 2.684243e-07, 2.684244e-07, 2.684243e-07, 
    2.684244e-07, 2.684262e-07, 2.684261e-07, 2.684261e-07, 2.68426e-07, 
    2.684261e-07, 2.684258e-07, 2.684257e-07, 2.684253e-07, 2.684255e-07, 
    2.684252e-07, 2.684255e-07, 2.684254e-07, 2.684252e-07, 2.684255e-07, 
    2.684249e-07, 2.684253e-07, 2.684247e-07, 2.68425e-07, 2.684246e-07, 
    2.684247e-07, 2.684246e-07, 2.684245e-07, 2.684244e-07, 2.684241e-07, 
    2.684242e-07, 2.68424e-07, 2.68426e-07, 2.684258e-07, 2.684259e-07, 
    2.684257e-07, 2.684256e-07, 2.684254e-07, 2.684251e-07, 2.684253e-07, 
    2.68425e-07, 2.68425e-07, 2.684253e-07, 2.684251e-07, 2.684258e-07, 
    2.684257e-07, 2.684257e-07, 2.684259e-07, 2.684252e-07, 2.684256e-07, 
    2.684249e-07, 2.684251e-07, 2.684245e-07, 2.684248e-07, 2.684242e-07, 
    2.68424e-07, 2.684237e-07, 2.684235e-07, 2.684258e-07, 2.684259e-07, 
    2.684257e-07, 2.684255e-07, 2.684253e-07, 2.684251e-07, 2.684251e-07, 
    2.68425e-07, 2.684249e-07, 2.684248e-07, 2.68425e-07, 2.684248e-07, 
    2.684256e-07, 2.684252e-07, 2.684259e-07, 2.684257e-07, 2.684255e-07, 
    2.684256e-07, 2.684253e-07, 2.684252e-07, 2.684249e-07, 2.68425e-07, 
    2.68424e-07, 2.684245e-07, 2.684233e-07, 2.684236e-07, 2.684259e-07, 
    2.684258e-07, 2.684254e-07, 2.684256e-07, 2.684251e-07, 2.684249e-07, 
    2.684249e-07, 2.684247e-07, 2.684247e-07, 2.684246e-07, 2.684247e-07, 
    2.684246e-07, 2.684251e-07, 2.684249e-07, 2.684255e-07, 2.684253e-07, 
    2.684254e-07, 2.684254e-07, 2.684252e-07, 2.68425e-07, 2.68425e-07, 
    2.684249e-07, 2.684247e-07, 2.684251e-07, 2.68424e-07, 2.684247e-07, 
    2.684257e-07, 2.684255e-07, 2.684254e-07, 2.684255e-07, 2.68425e-07, 
    2.684251e-07, 2.684246e-07, 2.684248e-07, 2.684245e-07, 2.684247e-07, 
    2.684247e-07, 2.684248e-07, 2.684249e-07, 2.684251e-07, 2.684253e-07, 
    2.684255e-07, 2.684255e-07, 2.684253e-07, 2.68425e-07, 2.684247e-07, 
    2.684248e-07, 2.684245e-07, 2.684251e-07, 2.684249e-07, 2.68425e-07, 
    2.684247e-07, 2.684253e-07, 2.684248e-07, 2.684254e-07, 2.684253e-07, 
    2.684252e-07, 2.684249e-07, 2.684248e-07, 2.684247e-07, 2.684248e-07, 
    2.68425e-07, 2.68425e-07, 2.684252e-07, 2.684252e-07, 2.684253e-07, 
    2.684254e-07, 2.684253e-07, 2.684252e-07, 2.68425e-07, 2.684247e-07, 
    2.684245e-07, 2.684244e-07, 2.684241e-07, 2.684244e-07, 2.68424e-07, 
    2.684243e-07, 2.684237e-07, 2.684248e-07, 2.684243e-07, 2.684251e-07, 
    2.684251e-07, 2.684249e-07, 2.684245e-07, 2.684247e-07, 2.684245e-07, 
    2.68425e-07, 2.684253e-07, 2.684253e-07, 2.684255e-07, 2.684253e-07, 
    2.684254e-07, 2.684252e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684247e-07, 2.684245e-07, 2.68424e-07, 2.684237e-07, 2.684234e-07, 
    2.684233e-07, 2.684233e-07, 2.684233e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  5.637083e-26, 1.593089e-25, 8.578169e-26, -3.186177e-26, -1.642107e-25, 
    -3.676358e-26, 1.127417e-25, 1.936215e-25, -6.862535e-26, -1.151926e-25, 
    -1.225453e-26, -6.617445e-26, 1.249962e-25, -5.391992e-26, 6.372354e-26, 
    8.578169e-26, 7.107626e-26, -6.127264e-26, 1.470543e-25, -1.862688e-25, 
    7.842898e-26, -1.764652e-25, 6.617445e-26, -7.352717e-27, 1.249962e-25, 
    -2.377378e-25, -9.803622e-26, -1.519561e-25, -4.41163e-26, -3.431268e-26, 
    5.637083e-26, 2.156797e-25, -4.41163e-26, -5.882173e-26, 7.352717e-27, 
    1.593089e-25, -2.205815e-26, 9.558531e-26, -1.102908e-25, -8.82326e-26, 
    1.323489e-25, -2.695996e-26, -6.862535e-26, 1.249962e-25, -2.009742e-25, 
    2.59796e-25, -5.391992e-26, 6.372354e-26, 3.308722e-25, 1.004871e-25, 
    -1.936215e-25, 8.087988e-26, -8.82326e-26, -5.637083e-26, 8.333079e-26, 
    1.446034e-25, 1.102908e-25, 1.02938e-25, 8.087988e-26, -1.225453e-26, 
    -7.652491e-42, 8.333079e-26, -1.127417e-25, 1.960724e-26, 1.715634e-25, 
    -1.274471e-25, 9.068351e-26, -3.676358e-26, -2.941087e-26, 1.347998e-25, 
    -2.450906e-27, -1.200944e-25, -2.450905e-26, 1.200944e-25, -1.053889e-25, 
    1.838179e-25, -2.254833e-25, -1.960724e-26, 5.146902e-26, -3.921449e-26, 
    -1.249962e-25, 1.530638e-41, -1.225453e-26, 1.053889e-25, -4.901811e-26, 
    7.842898e-26, 1.176435e-25, -2.352869e-25, 1.078398e-25, 4.901811e-27, 
    -6.372354e-26, -1.446034e-25, 1.764652e-25, -1.764652e-25, 2.181306e-25, 
    -1.446034e-25, 4.65672e-26, 8.087988e-26, 1.102908e-25, 1.004871e-25, 
    3.921449e-26, -9.313441e-26, -9.313441e-26, 1.053889e-25, 7.352717e-27, 
    2.254833e-25, 3.431268e-26, 7.352717e-27, -1.372507e-25, -1.176435e-25, 
    -2.107779e-25, -7.107626e-26, -1.225453e-25, -1.397016e-25, 2.450905e-26, 
    -1.519561e-25, 1.54407e-25, 1.176435e-25, -5.391992e-26, 5.146902e-26, 
    1.715634e-25, 5.391992e-26, 2.450906e-27, -1.960724e-26, 1.053889e-25, 
    1.56858e-25, 1.911706e-25, 3.014614e-25, -8.333079e-26, -1.176435e-25, 
    -4.901811e-27, 7.842898e-26, -1.789161e-25, -2.990105e-25, -3.431268e-26, 
    2.695996e-26, -3.676358e-26, -1.225453e-26, 1.102908e-25, 9.803622e-27, 
    -9.068351e-26, 1.519561e-25, 7.597807e-26, -2.303851e-25, 2.303851e-25, 
    -4.166539e-26, 3.676358e-26, -8.087988e-26, 2.941087e-26, -1.421525e-25, 
    9.803622e-27, -2.941087e-25, 6.372354e-26, -1.838179e-25, 2.941087e-26, 
    4.41163e-26, 1.29898e-25, 1.911706e-25, 1.936215e-25, -4.901811e-27, 
    -1.470543e-25, 7.107626e-26, -7.842898e-26, -7.842898e-26, -1.56858e-25, 
    1.960724e-26, 1.642107e-25, -6.127264e-26, 4.901811e-26, 1.715634e-26, 
    2.205815e-26, -1.789161e-25, -1.274471e-25, -5.146902e-26, 2.941087e-26, 
    9.558531e-26, 8.82326e-26, -3.676358e-26, -4.901811e-26, 1.225453e-26, 
    -2.034252e-25, -6.862535e-26, 1.470543e-26, 1.02938e-25, -3.431268e-26, 
    2.450905e-26, -1.372507e-25, 6.617445e-26, 6.617445e-26, -4.166539e-26, 
    2.205815e-25, -1.470543e-25, -6.617445e-26, -1.691125e-25, -7.352717e-27, 
    -9.068351e-26, -1.470543e-25, -8.333079e-26, -2.254833e-25, 
    -1.642107e-25, 8.333079e-26, -7.107626e-26, 3.186177e-26, 3.186177e-26, 
    2.450905e-26, -4.901811e-27, -1.960724e-26, 1.29898e-25, -1.887197e-25, 
    1.004871e-25, -8.578169e-26, 1.127417e-25, -1.495052e-25, -4.901811e-27, 
    -2.254833e-25, -3.676358e-26, -1.151926e-25, 8.578169e-26, -3.921449e-26, 
    -3.431268e-26, 2.941087e-26, 4.901811e-27, 1.911706e-25, -1.960724e-26, 
    -1.470543e-25, 1.691125e-25, 1.642107e-25, -8.333079e-26, 7.597807e-26, 
    -1.200944e-25, 4.65672e-26, -7.352717e-26, -1.249962e-25, -2.205815e-26, 
    9.803622e-27, 1.617598e-25, -9.313441e-26, -2.230324e-25, -3.431268e-26, 
    -1.715634e-26, -7.107626e-26, -7.597807e-26, -2.303851e-25, 
    -2.009742e-25, -3.259704e-25, -1.176435e-25, -5.637083e-26, 1.078398e-25, 
    3.11265e-25, 2.058761e-25, 3.872431e-25, 1.004871e-25, 1.715634e-26, 
    2.303851e-25, 8.578169e-26, 2.08327e-25, 1.960724e-26, -1.225453e-25, 
    9.803622e-26, 2.794032e-25, 1.495052e-25, 1.911706e-25, 1.274471e-25, 
    1.249962e-25, 9.558531e-26, 2.475414e-25, -4.166539e-26, 2.303851e-25, 
    2.818541e-25, -3.161668e-25, 1.519561e-25, -1.372507e-25, 2.941087e-26, 
    1.789161e-25, 3.186177e-26, 6.127264e-26, 2.695996e-26, 6.372354e-26, 
    1.249962e-25, -8.578169e-26, 1.56858e-25, -3.039123e-25, -2.107779e-25, 
    -2.671487e-25, 3.186177e-26, -1.470543e-26, -3.431268e-26, -1.470543e-25, 
    5.391992e-26, -4.41163e-26, 4.901811e-26, -7.352717e-27, 1.446034e-25, 
    2.450906e-27, -1.225453e-25, 3.872431e-25, 2.034252e-25, 1.397016e-25, 
    -7.352717e-26, -1.960724e-26, -9.068351e-26, 2.695996e-26, -2.622469e-25, 
    -1.519561e-25, 1.960724e-25, 3.676358e-25, -5.146902e-26, -1.446034e-25, 
    2.695996e-26, -6.127264e-26, -4.166539e-26, 1.740143e-25, -2.524433e-25, 
    -2.695996e-26, -9.803622e-27, 9.068351e-26, -1.789161e-25, 6.372354e-26, 
    -2.181306e-25, -6.862535e-26, -1.200944e-25, 8.578169e-26, -1.053889e-25, 
    1.200944e-25, -1.960724e-26, -1.740143e-25, 2.941087e-26, 3.431268e-25, 
    -7.842898e-26, 1.200944e-25, -1.960724e-26, 6.127264e-26, -7.842898e-26, 
    1.715634e-26, -2.32836e-25, -1.495052e-25, 1.470543e-26, -2.794032e-25,
  2.676251e-32, 2.676248e-32, 2.676249e-32, 2.676247e-32, 2.676248e-32, 
    2.676246e-32, 2.67625e-32, 2.676248e-32, 2.676249e-32, 2.676251e-32, 
    2.676242e-32, 2.676246e-32, 2.676238e-32, 2.676241e-32, 2.676234e-32, 
    2.676238e-32, 2.676233e-32, 2.676234e-32, 2.676231e-32, 2.676232e-32, 
    2.676228e-32, 2.676231e-32, 2.676226e-32, 2.676229e-32, 2.676228e-32, 
    2.676231e-32, 2.676246e-32, 2.676243e-32, 2.676246e-32, 2.676245e-32, 
    2.676245e-32, 2.676248e-32, 2.676249e-32, 2.676251e-32, 2.676251e-32, 
    2.676249e-32, 2.676245e-32, 2.676247e-32, 2.676243e-32, 2.676243e-32, 
    2.676239e-32, 2.676241e-32, 2.676235e-32, 2.676237e-32, 2.676232e-32, 
    2.676233e-32, 2.676232e-32, 2.676232e-32, 2.676232e-32, 2.676234e-32, 
    2.676233e-32, 2.676234e-32, 2.676241e-32, 2.676239e-32, 2.676244e-32, 
    2.676248e-32, 2.67625e-32, 2.676252e-32, 2.676252e-32, 2.676251e-32, 
    2.676249e-32, 2.676247e-32, 2.676245e-32, 2.676244e-32, 2.676243e-32, 
    2.67624e-32, 2.676238e-32, 2.676235e-32, 2.676235e-32, 2.676234e-32, 
    2.676233e-32, 2.676232e-32, 2.676232e-32, 2.676231e-32, 2.676234e-32, 
    2.676232e-32, 2.676236e-32, 2.676235e-32, 2.676243e-32, 2.676246e-32, 
    2.676247e-32, 2.676249e-32, 2.676251e-32, 2.676249e-32, 2.67625e-32, 
    2.676248e-32, 2.676247e-32, 2.676248e-32, 2.676244e-32, 2.676246e-32, 
    2.676238e-32, 2.676242e-32, 2.676233e-32, 2.676235e-32, 2.676233e-32, 
    2.676234e-32, 2.676232e-32, 2.676234e-32, 2.676231e-32, 2.67623e-32, 
    2.67623e-32, 2.676229e-32, 2.676234e-32, 2.676232e-32, 2.676248e-32, 
    2.676248e-32, 2.676247e-32, 2.676249e-32, 2.676249e-32, 2.676251e-32, 
    2.676249e-32, 2.676249e-32, 2.676247e-32, 2.676246e-32, 2.676245e-32, 
    2.676243e-32, 2.676241e-32, 2.676237e-32, 2.676235e-32, 2.676234e-32, 
    2.676234e-32, 2.676234e-32, 2.676235e-32, 2.676235e-32, 2.67623e-32, 
    2.676233e-32, 2.676229e-32, 2.676229e-32, 2.676231e-32, 2.676229e-32, 
    2.676248e-32, 2.676248e-32, 2.67625e-32, 2.676249e-32, 2.676251e-32, 
    2.67625e-32, 2.676249e-32, 2.676246e-32, 2.676245e-32, 2.676244e-32, 
    2.676243e-32, 2.676241e-32, 2.676238e-32, 2.676236e-32, 2.676233e-32, 
    2.676233e-32, 2.676233e-32, 2.676233e-32, 2.676234e-32, 2.676232e-32, 
    2.676232e-32, 2.676233e-32, 2.676229e-32, 2.67623e-32, 2.676229e-32, 
    2.67623e-32, 2.676248e-32, 2.676247e-32, 2.676248e-32, 2.676247e-32, 
    2.676247e-32, 2.676244e-32, 2.676244e-32, 2.676239e-32, 2.676241e-32, 
    2.676239e-32, 2.676241e-32, 2.67624e-32, 2.676238e-32, 2.676241e-32, 
    2.676236e-32, 2.676239e-32, 2.676233e-32, 2.676236e-32, 2.676232e-32, 
    2.676233e-32, 2.676232e-32, 2.676231e-32, 2.67623e-32, 2.676227e-32, 
    2.676228e-32, 2.676226e-32, 2.676246e-32, 2.676244e-32, 2.676245e-32, 
    2.676243e-32, 2.676242e-32, 2.676241e-32, 2.676237e-32, 2.676239e-32, 
    2.676236e-32, 2.676236e-32, 2.676239e-32, 2.676237e-32, 2.676244e-32, 
    2.676243e-32, 2.676243e-32, 2.676246e-32, 2.676238e-32, 2.676242e-32, 
    2.676235e-32, 2.676237e-32, 2.676231e-32, 2.676234e-32, 2.676228e-32, 
    2.676226e-32, 2.676224e-32, 2.676221e-32, 2.676244e-32, 2.676245e-32, 
    2.676243e-32, 2.676241e-32, 2.676239e-32, 2.676237e-32, 2.676237e-32, 
    2.676236e-32, 2.676235e-32, 2.676234e-32, 2.676236e-32, 2.676234e-32, 
    2.676242e-32, 2.676238e-32, 2.676245e-32, 2.676243e-32, 2.676242e-32, 
    2.676242e-32, 2.676239e-32, 2.676238e-32, 2.676235e-32, 2.676236e-32, 
    2.676227e-32, 2.676231e-32, 2.676219e-32, 2.676222e-32, 2.676245e-32, 
    2.676244e-32, 2.67624e-32, 2.676242e-32, 2.676237e-32, 2.676236e-32, 
    2.676234e-32, 2.676233e-32, 2.676233e-32, 2.676232e-32, 2.676234e-32, 
    2.676232e-32, 2.676237e-32, 2.676235e-32, 2.676241e-32, 2.676239e-32, 
    2.67624e-32, 2.676241e-32, 2.676238e-32, 2.676236e-32, 2.676236e-32, 
    2.676235e-32, 2.676233e-32, 2.676237e-32, 2.676226e-32, 2.676233e-32, 
    2.676243e-32, 2.676241e-32, 2.67624e-32, 2.676241e-32, 2.676236e-32, 
    2.676238e-32, 2.676232e-32, 2.676234e-32, 2.676232e-32, 2.676233e-32, 
    2.676233e-32, 2.676234e-32, 2.676235e-32, 2.676238e-32, 2.676239e-32, 
    2.676241e-32, 2.676241e-32, 2.676239e-32, 2.676236e-32, 2.676233e-32, 
    2.676234e-32, 2.676232e-32, 2.676237e-32, 2.676235e-32, 2.676236e-32, 
    2.676233e-32, 2.676239e-32, 2.676234e-32, 2.67624e-32, 2.676239e-32, 
    2.676238e-32, 2.676235e-32, 2.676234e-32, 2.676233e-32, 2.676234e-32, 
    2.676236e-32, 2.676236e-32, 2.676238e-32, 2.676238e-32, 2.676239e-32, 
    2.67624e-32, 2.676239e-32, 2.676239e-32, 2.676236e-32, 2.676234e-32, 
    2.676231e-32, 2.67623e-32, 2.676227e-32, 2.67623e-32, 2.676226e-32, 
    2.676229e-32, 2.676223e-32, 2.676234e-32, 2.676229e-32, 2.676238e-32, 
    2.676237e-32, 2.676235e-32, 2.676232e-32, 2.676234e-32, 2.676231e-32, 
    2.676236e-32, 2.676239e-32, 2.67624e-32, 2.676241e-32, 2.67624e-32, 
    2.67624e-32, 2.676239e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676233e-32, 2.676231e-32, 2.676226e-32, 2.676223e-32, 2.67622e-32, 
    2.676219e-32, 2.676219e-32, 2.676219e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  2.944134e-15, 2.952113e-15, 2.950563e-15, 2.956993e-15, 2.953428e-15, 
    2.957636e-15, 2.945754e-15, 2.952429e-15, 2.948169e-15, 2.944854e-15, 
    2.969452e-15, 2.95728e-15, 2.982086e-15, 2.974336e-15, 2.99379e-15, 
    2.980879e-15, 2.996392e-15, 2.993421e-15, 3.002366e-15, 2.999805e-15, 
    3.011228e-15, 3.003548e-15, 3.017148e-15, 3.009396e-15, 3.010609e-15, 
    3.003294e-15, 2.959733e-15, 2.967936e-15, 2.959246e-15, 2.960417e-15, 
    2.959892e-15, 2.9535e-15, 2.950275e-15, 2.943526e-15, 2.944752e-15, 
    2.949711e-15, 2.960943e-15, 2.957134e-15, 2.966736e-15, 2.96652e-15, 
    2.977194e-15, 2.972383e-15, 2.990303e-15, 2.985216e-15, 2.999912e-15, 
    2.996218e-15, 2.999738e-15, 2.998671e-15, 2.999752e-15, 2.994333e-15, 
    2.996655e-15, 2.991887e-15, 2.973284e-15, 2.978755e-15, 2.962424e-15, 
    2.952582e-15, 2.946046e-15, 2.941402e-15, 2.942059e-15, 2.94331e-15, 
    2.949739e-15, 2.955782e-15, 2.960383e-15, 2.963459e-15, 2.966489e-15, 
    2.975645e-15, 2.980493e-15, 2.99133e-15, 2.989377e-15, 2.992687e-15, 
    2.99585e-15, 3.001155e-15, 3.000283e-15, 3.002619e-15, 2.992601e-15, 
    2.999259e-15, 2.988266e-15, 2.991273e-15, 2.967303e-15, 2.958162e-15, 
    2.954266e-15, 2.950861e-15, 2.942563e-15, 2.948294e-15, 2.946035e-15, 
    2.95141e-15, 2.954821e-15, 2.953134e-15, 2.963543e-15, 2.959498e-15, 
    2.98078e-15, 2.97162e-15, 2.995481e-15, 2.989778e-15, 2.996848e-15, 
    2.993242e-15, 2.999419e-15, 2.99386e-15, 3.003488e-15, 3.005582e-15, 
    3.004151e-15, 3.00965e-15, 2.993551e-15, 2.999737e-15, 2.953087e-15, 
    2.953362e-15, 2.954644e-15, 2.949005e-15, 2.94866e-15, 2.943492e-15, 
    2.948092e-15, 2.950049e-15, 2.95502e-15, 2.957957e-15, 2.960748e-15, 
    2.966882e-15, 2.973725e-15, 2.983286e-15, 2.990148e-15, 2.994745e-15, 
    2.991927e-15, 2.994415e-15, 2.991633e-15, 2.99033e-15, 3.004797e-15, 
    2.996676e-15, 3.008859e-15, 3.008186e-15, 3.002674e-15, 3.008262e-15, 
    2.953555e-15, 2.951972e-15, 2.946469e-15, 2.950776e-15, 2.942929e-15, 
    2.947321e-15, 2.949845e-15, 2.95958e-15, 2.96172e-15, 2.9637e-15, 
    2.967613e-15, 2.97263e-15, 2.981422e-15, 2.989063e-15, 2.996035e-15, 
    2.995524e-15, 2.995704e-15, 2.997259e-15, 2.993404e-15, 2.997892e-15, 
    2.998644e-15, 2.996676e-15, 3.008096e-15, 3.004835e-15, 3.008172e-15, 
    3.006049e-15, 2.952487e-15, 2.955151e-15, 2.953711e-15, 2.956418e-15, 
    2.95451e-15, 2.962986e-15, 2.965525e-15, 2.977399e-15, 2.97253e-15, 
    2.980279e-15, 2.973319e-15, 2.974552e-15, 2.980528e-15, 2.973696e-15, 
    2.988641e-15, 2.978508e-15, 2.99732e-15, 2.98721e-15, 2.997953e-15, 
    2.996004e-15, 2.999231e-15, 3.002119e-15, 3.005751e-15, 3.012447e-15, 
    3.010898e-15, 3.016495e-15, 2.959122e-15, 2.962574e-15, 2.962272e-15, 
    2.965884e-15, 2.968554e-15, 2.974339e-15, 2.983608e-15, 2.980124e-15, 
    2.98652e-15, 2.987803e-15, 2.978087e-15, 2.984052e-15, 2.964885e-15, 
    2.967983e-15, 2.96614e-15, 2.959394e-15, 2.980925e-15, 2.969882e-15, 
    2.990261e-15, 2.98429e-15, 3.001707e-15, 2.993047e-15, 3.010044e-15, 
    3.017293e-15, 3.024118e-15, 3.032075e-15, 2.964459e-15, 2.962114e-15, 
    2.966314e-15, 2.972117e-15, 2.977503e-15, 2.984654e-15, 2.985386e-15, 
    2.986725e-15, 2.990191e-15, 2.993104e-15, 2.987146e-15, 2.993835e-15, 
    2.968698e-15, 2.981883e-15, 2.961226e-15, 2.96745e-15, 2.971776e-15, 
    2.96988e-15, 2.979727e-15, 2.982045e-15, 2.991455e-15, 2.986594e-15, 
    3.015503e-15, 3.002726e-15, 3.038134e-15, 3.028255e-15, 2.961294e-15, 
    2.964452e-15, 2.975428e-15, 2.970208e-15, 2.985132e-15, 2.9888e-15, 
    2.991781e-15, 2.995589e-15, 2.996001e-15, 2.998256e-15, 2.99456e-15, 
    2.998111e-15, 2.984669e-15, 2.990678e-15, 2.974177e-15, 2.978196e-15, 
    2.976348e-15, 2.974319e-15, 2.980579e-15, 2.98724e-15, 2.987385e-15, 
    2.989517e-15, 2.995522e-15, 2.985193e-15, 3.017146e-15, 2.997422e-15, 
    2.967893e-15, 2.973965e-15, 2.974835e-15, 2.972484e-15, 2.988433e-15, 
    2.982657e-15, 2.998202e-15, 2.994004e-15, 3.000881e-15, 2.997464e-15, 
    2.996961e-15, 2.992571e-15, 2.989835e-15, 2.982922e-15, 2.977291e-15, 
    2.972825e-15, 2.973864e-15, 2.978769e-15, 2.987647e-15, 2.996037e-15, 
    2.994199e-15, 3.000359e-15, 2.984051e-15, 2.990891e-15, 2.988248e-15, 
    2.995141e-15, 2.980031e-15, 2.992891e-15, 2.976739e-15, 2.978157e-15, 
    2.982543e-15, 2.991353e-15, 2.993305e-15, 2.995384e-15, 2.994102e-15, 
    2.987873e-15, 2.986853e-15, 2.982437e-15, 2.981215e-15, 2.977849e-15, 
    2.975059e-15, 2.977607e-15, 2.980282e-15, 2.987877e-15, 2.994712e-15, 
    3.002159e-15, 3.003982e-15, 3.012665e-15, 3.005593e-15, 3.017255e-15, 
    3.007335e-15, 3.024501e-15, 2.99364e-15, 3.007049e-15, 2.982743e-15, 
    2.985366e-15, 2.990104e-15, 3.000969e-15, 2.995108e-15, 3.001963e-15, 
    2.986814e-15, 2.978937e-15, 2.976901e-15, 2.973096e-15, 2.976988e-15, 
    2.976672e-15, 2.980395e-15, 2.979199e-15, 2.988129e-15, 2.983333e-15, 
    2.996948e-15, 3.00191e-15, 3.015908e-15, 3.024474e-15, 3.033188e-15, 
    3.03703e-15, 3.038199e-15, 3.038688e-15 ;

 LITR2N_vr =
  1.532743e-05, 1.532741e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 
    1.53274e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 1.532743e-05, 
    1.532738e-05, 1.53274e-05, 1.532735e-05, 1.532737e-05, 1.532733e-05, 
    1.532736e-05, 1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532732e-05, 
    1.53273e-05, 1.532731e-05, 1.532729e-05, 1.53273e-05, 1.53273e-05, 
    1.532731e-05, 1.53274e-05, 1.532738e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532737e-05, 1.532734e-05, 1.532735e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532733e-05, 
    1.532733e-05, 1.532734e-05, 1.532737e-05, 1.532736e-05, 1.532739e-05, 
    1.532741e-05, 1.532742e-05, 1.532743e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 
    1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532733e-05, 
    1.532732e-05, 1.532734e-05, 1.532734e-05, 1.532738e-05, 1.53274e-05, 
    1.532741e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 
    1.532736e-05, 1.532738e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532731e-05, 1.532731e-05, 
    1.532731e-05, 1.53273e-05, 1.532733e-05, 1.532732e-05, 1.532741e-05, 
    1.532741e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532734e-05, 1.532733e-05, 
    1.532734e-05, 1.532733e-05, 1.532734e-05, 1.532734e-05, 1.532731e-05, 
    1.532733e-05, 1.53273e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.532741e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 
    1.532742e-05, 1.532742e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.532731e-05, 1.532741e-05, 1.532741e-05, 1.532741e-05, 1.53274e-05, 
    1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532736e-05, 1.532737e-05, 
    1.532736e-05, 1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532737e-05, 
    1.532734e-05, 1.532736e-05, 1.532732e-05, 1.532734e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 
    1.53273e-05, 1.532729e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532736e-05, 
    1.532735e-05, 1.532734e-05, 1.532736e-05, 1.532735e-05, 1.532739e-05, 
    1.532738e-05, 1.532738e-05, 1.53274e-05, 1.532736e-05, 1.532738e-05, 
    1.532734e-05, 1.532735e-05, 1.532732e-05, 1.532733e-05, 1.53273e-05, 
    1.532729e-05, 1.532727e-05, 1.532726e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532735e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532738e-05, 1.532736e-05, 1.53274e-05, 1.532738e-05, 1.532737e-05, 
    1.532738e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532735e-05, 
    1.532729e-05, 1.532731e-05, 1.532725e-05, 1.532726e-05, 1.53274e-05, 
    1.532739e-05, 1.532737e-05, 1.532738e-05, 1.532735e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532733e-05, 
    1.532732e-05, 1.532735e-05, 1.532734e-05, 1.532737e-05, 1.532736e-05, 
    1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532735e-05, 1.532729e-05, 1.532732e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 1.532732e-05, 
    1.532733e-05, 1.532733e-05, 1.532734e-05, 1.532735e-05, 1.532736e-05, 
    1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532736e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532733e-05, 
    1.532734e-05, 1.532734e-05, 1.532735e-05, 1.532736e-05, 1.532736e-05, 
    1.532737e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532732e-05, 1.532731e-05, 1.53273e-05, 1.532731e-05, 1.532729e-05, 
    1.532731e-05, 1.532727e-05, 1.532733e-05, 1.532731e-05, 1.532735e-05, 
    1.532735e-05, 1.532734e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532734e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532733e-05, 1.532732e-05, 1.532729e-05, 1.532727e-05, 1.532726e-05, 
    1.532725e-05, 1.532725e-05, 1.532724e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.063689e-13, 1.066571e-13, 1.066011e-13, 1.068334e-13, 1.067046e-13, 
    1.068567e-13, 1.064274e-13, 1.066685e-13, 1.065146e-13, 1.063949e-13, 
    1.072836e-13, 1.068438e-13, 1.0774e-13, 1.074601e-13, 1.081629e-13, 
    1.076964e-13, 1.082569e-13, 1.081496e-13, 1.084727e-13, 1.083802e-13, 
    1.087929e-13, 1.085154e-13, 1.090068e-13, 1.087267e-13, 1.087705e-13, 
    1.085063e-13, 1.069325e-13, 1.072288e-13, 1.069149e-13, 1.069572e-13, 
    1.069382e-13, 1.067073e-13, 1.065908e-13, 1.063469e-13, 1.063912e-13, 
    1.065703e-13, 1.069762e-13, 1.068385e-13, 1.071855e-13, 1.071776e-13, 
    1.075633e-13, 1.073895e-13, 1.080369e-13, 1.078531e-13, 1.083841e-13, 
    1.082506e-13, 1.083778e-13, 1.083392e-13, 1.083783e-13, 1.081825e-13, 
    1.082664e-13, 1.080941e-13, 1.07422e-13, 1.076197e-13, 1.070297e-13, 
    1.066741e-13, 1.064379e-13, 1.062702e-13, 1.062939e-13, 1.063391e-13, 
    1.065714e-13, 1.067897e-13, 1.069559e-13, 1.070671e-13, 1.071765e-13, 
    1.075073e-13, 1.076825e-13, 1.08074e-13, 1.080035e-13, 1.08123e-13, 
    1.082373e-13, 1.08429e-13, 1.083975e-13, 1.084819e-13, 1.081199e-13, 
    1.083605e-13, 1.079633e-13, 1.08072e-13, 1.072059e-13, 1.068757e-13, 
    1.067349e-13, 1.066119e-13, 1.063121e-13, 1.065192e-13, 1.064376e-13, 
    1.066317e-13, 1.06755e-13, 1.06694e-13, 1.070701e-13, 1.069239e-13, 
    1.076929e-13, 1.073619e-13, 1.08224e-13, 1.08018e-13, 1.082734e-13, 
    1.081431e-13, 1.083663e-13, 1.081654e-13, 1.085133e-13, 1.085889e-13, 
    1.085372e-13, 1.087359e-13, 1.081543e-13, 1.083777e-13, 1.066923e-13, 
    1.067023e-13, 1.067486e-13, 1.065449e-13, 1.065324e-13, 1.063457e-13, 
    1.065119e-13, 1.065826e-13, 1.067622e-13, 1.068683e-13, 1.069691e-13, 
    1.071907e-13, 1.07438e-13, 1.077834e-13, 1.080313e-13, 1.081974e-13, 
    1.080956e-13, 1.081855e-13, 1.08085e-13, 1.080379e-13, 1.085606e-13, 
    1.082672e-13, 1.087073e-13, 1.08683e-13, 1.084839e-13, 1.086858e-13, 
    1.067092e-13, 1.06652e-13, 1.064532e-13, 1.066088e-13, 1.063253e-13, 
    1.06484e-13, 1.065752e-13, 1.069269e-13, 1.070042e-13, 1.070758e-13, 
    1.072171e-13, 1.073984e-13, 1.07716e-13, 1.079921e-13, 1.08244e-13, 
    1.082255e-13, 1.08232e-13, 1.082882e-13, 1.081489e-13, 1.083111e-13, 
    1.083383e-13, 1.082672e-13, 1.086797e-13, 1.085619e-13, 1.086825e-13, 
    1.086058e-13, 1.066706e-13, 1.067669e-13, 1.067149e-13, 1.068127e-13, 
    1.067438e-13, 1.0705e-13, 1.071417e-13, 1.075707e-13, 1.073948e-13, 
    1.076748e-13, 1.074233e-13, 1.074678e-13, 1.076837e-13, 1.074369e-13, 
    1.079769e-13, 1.076108e-13, 1.082904e-13, 1.079252e-13, 1.083133e-13, 
    1.082429e-13, 1.083595e-13, 1.084638e-13, 1.085951e-13, 1.08837e-13, 
    1.08781e-13, 1.089832e-13, 1.069104e-13, 1.070351e-13, 1.070242e-13, 
    1.071547e-13, 1.072511e-13, 1.074602e-13, 1.07795e-13, 1.076692e-13, 
    1.079002e-13, 1.079466e-13, 1.075955e-13, 1.078111e-13, 1.071186e-13, 
    1.072305e-13, 1.071639e-13, 1.069202e-13, 1.076981e-13, 1.072991e-13, 
    1.080354e-13, 1.078197e-13, 1.084489e-13, 1.081361e-13, 1.087501e-13, 
    1.090121e-13, 1.092586e-13, 1.095461e-13, 1.071032e-13, 1.070185e-13, 
    1.071702e-13, 1.073799e-13, 1.075745e-13, 1.078328e-13, 1.078593e-13, 
    1.079076e-13, 1.080329e-13, 1.081381e-13, 1.079229e-13, 1.081645e-13, 
    1.072563e-13, 1.077327e-13, 1.069864e-13, 1.072113e-13, 1.073676e-13, 
    1.072991e-13, 1.076548e-13, 1.077385e-13, 1.080785e-13, 1.079029e-13, 
    1.089474e-13, 1.084857e-13, 1.09765e-13, 1.094081e-13, 1.069889e-13, 
    1.071029e-13, 1.074995e-13, 1.073109e-13, 1.078501e-13, 1.079826e-13, 
    1.080903e-13, 1.082279e-13, 1.082428e-13, 1.083243e-13, 1.081907e-13, 
    1.08319e-13, 1.078334e-13, 1.080505e-13, 1.074543e-13, 1.075995e-13, 
    1.075327e-13, 1.074594e-13, 1.076856e-13, 1.079262e-13, 1.079315e-13, 
    1.080085e-13, 1.082255e-13, 1.078523e-13, 1.090067e-13, 1.082941e-13, 
    1.072273e-13, 1.074466e-13, 1.074781e-13, 1.073931e-13, 1.079693e-13, 
    1.077607e-13, 1.083223e-13, 1.081706e-13, 1.084191e-13, 1.082956e-13, 
    1.082775e-13, 1.081188e-13, 1.0802e-13, 1.077702e-13, 1.075668e-13, 
    1.074055e-13, 1.07443e-13, 1.076202e-13, 1.07941e-13, 1.082441e-13, 
    1.081777e-13, 1.084002e-13, 1.07811e-13, 1.080582e-13, 1.079627e-13, 
    1.082117e-13, 1.076658e-13, 1.081304e-13, 1.075469e-13, 1.075981e-13, 
    1.077565e-13, 1.080748e-13, 1.081454e-13, 1.082205e-13, 1.081742e-13, 
    1.079491e-13, 1.079123e-13, 1.077527e-13, 1.077086e-13, 1.07587e-13, 
    1.074862e-13, 1.075782e-13, 1.076749e-13, 1.079493e-13, 1.081962e-13, 
    1.084653e-13, 1.085311e-13, 1.088448e-13, 1.085893e-13, 1.090106e-13, 
    1.086523e-13, 1.092724e-13, 1.081575e-13, 1.086419e-13, 1.077638e-13, 
    1.078586e-13, 1.080297e-13, 1.084223e-13, 1.082105e-13, 1.084582e-13, 
    1.079108e-13, 1.076263e-13, 1.075527e-13, 1.074152e-13, 1.075559e-13, 
    1.075444e-13, 1.076789e-13, 1.076357e-13, 1.079584e-13, 1.077851e-13, 
    1.08277e-13, 1.084563e-13, 1.08962e-13, 1.092715e-13, 1.095863e-13, 
    1.097251e-13, 1.097674e-13, 1.09785e-13 ;

 LITR3C =
  9.698e-06, 9.69799e-06, 9.697992e-06, 9.697985e-06, 9.697988e-06, 
    9.697984e-06, 9.697998e-06, 9.69799e-06, 9.697995e-06, 9.697999e-06, 
    9.697969e-06, 9.697984e-06, 9.697954e-06, 9.697963e-06, 9.697939e-06, 
    9.697955e-06, 9.697936e-06, 9.697939e-06, 9.697928e-06, 9.697932e-06, 
    9.697918e-06, 9.697927e-06, 9.697911e-06, 9.69792e-06, 9.697918e-06, 
    9.697927e-06, 9.697981e-06, 9.697971e-06, 9.697981e-06, 9.69798e-06, 
    9.697981e-06, 9.697988e-06, 9.697993e-06, 9.698001e-06, 9.697999e-06, 
    9.697993e-06, 9.697979e-06, 9.697984e-06, 9.697972e-06, 9.697973e-06, 
    9.697959e-06, 9.697966e-06, 9.697944e-06, 9.69795e-06, 9.697932e-06, 
    9.697937e-06, 9.697932e-06, 9.697933e-06, 9.697932e-06, 9.697938e-06, 
    9.697936e-06, 9.697942e-06, 9.697965e-06, 9.697957e-06, 9.697977e-06, 
    9.697989e-06, 9.697997e-06, 9.698004e-06, 9.698003e-06, 9.698001e-06, 
    9.697993e-06, 9.697986e-06, 9.69798e-06, 9.697977e-06, 9.697973e-06, 
    9.697961e-06, 9.697956e-06, 9.697942e-06, 9.697945e-06, 9.69794e-06, 
    9.697937e-06, 9.69793e-06, 9.697931e-06, 9.697928e-06, 9.697941e-06, 
    9.697933e-06, 9.697946e-06, 9.697942e-06, 9.697972e-06, 9.697983e-06, 
    9.697987e-06, 9.697992e-06, 9.698002e-06, 9.697995e-06, 9.697997e-06, 
    9.697991e-06, 9.697987e-06, 9.697989e-06, 9.697977e-06, 9.697981e-06, 
    9.697955e-06, 9.697967e-06, 9.697937e-06, 9.697944e-06, 9.697936e-06, 
    9.69794e-06, 9.697932e-06, 9.697939e-06, 9.697927e-06, 9.697925e-06, 
    9.697927e-06, 9.69792e-06, 9.697939e-06, 9.697932e-06, 9.697989e-06, 
    9.697988e-06, 9.697987e-06, 9.697994e-06, 9.697995e-06, 9.698001e-06, 
    9.697996e-06, 9.697993e-06, 9.697987e-06, 9.697983e-06, 9.697979e-06, 
    9.697972e-06, 9.697964e-06, 9.697952e-06, 9.697944e-06, 9.697938e-06, 
    9.697941e-06, 9.697938e-06, 9.697942e-06, 9.697944e-06, 9.697926e-06, 
    9.697936e-06, 9.697921e-06, 9.697922e-06, 9.697928e-06, 9.697922e-06, 
    9.697988e-06, 9.69799e-06, 9.697997e-06, 9.697992e-06, 9.698001e-06, 
    9.697997e-06, 9.697993e-06, 9.697981e-06, 9.697978e-06, 9.697976e-06, 
    9.697971e-06, 9.697965e-06, 9.697955e-06, 9.697945e-06, 9.697937e-06, 
    9.697937e-06, 9.697937e-06, 9.697935e-06, 9.69794e-06, 9.697934e-06, 
    9.697933e-06, 9.697936e-06, 9.697922e-06, 9.697926e-06, 9.697922e-06, 
    9.697924e-06, 9.69799e-06, 9.697987e-06, 9.697988e-06, 9.697985e-06, 
    9.697987e-06, 9.697977e-06, 9.697974e-06, 9.697959e-06, 9.697966e-06, 
    9.697956e-06, 9.697965e-06, 9.697963e-06, 9.697956e-06, 9.697964e-06, 
    9.697946e-06, 9.697958e-06, 9.697935e-06, 9.697947e-06, 9.697934e-06, 
    9.697937e-06, 9.697933e-06, 9.697929e-06, 9.697925e-06, 9.697917e-06, 
    9.697918e-06, 9.697911e-06, 9.697982e-06, 9.697977e-06, 9.697977e-06, 
    9.697974e-06, 9.69797e-06, 9.697963e-06, 9.697952e-06, 9.697956e-06, 
    9.697948e-06, 9.697947e-06, 9.697958e-06, 9.697951e-06, 9.697975e-06, 
    9.697971e-06, 9.697973e-06, 9.697981e-06, 9.697955e-06, 9.697968e-06, 
    9.697944e-06, 9.697951e-06, 9.697929e-06, 9.69794e-06, 9.697919e-06, 
    9.69791e-06, 9.697902e-06, 9.697892e-06, 9.697975e-06, 9.697978e-06, 
    9.697973e-06, 9.697966e-06, 9.697959e-06, 9.69795e-06, 9.697949e-06, 
    9.697947e-06, 9.697944e-06, 9.69794e-06, 9.697947e-06, 9.697939e-06, 
    9.69797e-06, 9.697954e-06, 9.697979e-06, 9.697971e-06, 9.697967e-06, 
    9.697968e-06, 9.697957e-06, 9.697954e-06, 9.697942e-06, 9.697948e-06, 
    9.697913e-06, 9.697928e-06, 9.697885e-06, 9.697897e-06, 9.697979e-06, 
    9.697975e-06, 9.697962e-06, 9.697968e-06, 9.69795e-06, 9.697946e-06, 
    9.697942e-06, 9.697937e-06, 9.697937e-06, 9.697934e-06, 9.697938e-06, 
    9.697934e-06, 9.69795e-06, 9.697943e-06, 9.697963e-06, 9.697958e-06, 
    9.69796e-06, 9.697963e-06, 9.697956e-06, 9.697947e-06, 9.697947e-06, 
    9.697945e-06, 9.697937e-06, 9.69795e-06, 9.697911e-06, 9.697935e-06, 
    9.697971e-06, 9.697964e-06, 9.697962e-06, 9.697966e-06, 9.697946e-06, 
    9.697953e-06, 9.697934e-06, 9.697939e-06, 9.69793e-06, 9.697935e-06, 
    9.697936e-06, 9.697941e-06, 9.697944e-06, 9.697953e-06, 9.697959e-06, 
    9.697965e-06, 9.697964e-06, 9.697957e-06, 9.697947e-06, 9.697937e-06, 
    9.697938e-06, 9.697931e-06, 9.697951e-06, 9.697943e-06, 9.697946e-06, 
    9.697937e-06, 9.697957e-06, 9.69794e-06, 9.69796e-06, 9.697958e-06, 
    9.697953e-06, 9.697942e-06, 9.69794e-06, 9.697937e-06, 9.697939e-06, 
    9.697947e-06, 9.697947e-06, 9.697953e-06, 9.697955e-06, 9.697958e-06, 
    9.697962e-06, 9.697959e-06, 9.697956e-06, 9.697947e-06, 9.697938e-06, 
    9.697929e-06, 9.697927e-06, 9.697917e-06, 9.697925e-06, 9.69791e-06, 
    9.697923e-06, 9.697902e-06, 9.697939e-06, 9.697923e-06, 9.697953e-06, 
    9.697949e-06, 9.697944e-06, 9.69793e-06, 9.697937e-06, 9.697929e-06, 
    9.697947e-06, 9.697957e-06, 9.69796e-06, 9.697965e-06, 9.69796e-06, 
    9.69796e-06, 9.697956e-06, 9.697957e-06, 9.697947e-06, 9.697952e-06, 
    9.697936e-06, 9.697929e-06, 9.697912e-06, 9.697902e-06, 9.697891e-06, 
    9.697887e-06, 9.697885e-06, 9.697885e-06 ;

 LITR3C_TO_SOIL2C =
  5.318442e-14, 5.332856e-14, 5.330056e-14, 5.341671e-14, 5.33523e-14, 
    5.342833e-14, 5.321368e-14, 5.333426e-14, 5.32573e-14, 5.319743e-14, 
    5.364177e-14, 5.342189e-14, 5.387e-14, 5.373001e-14, 5.408143e-14, 
    5.38482e-14, 5.412843e-14, 5.407476e-14, 5.423635e-14, 5.419008e-14, 
    5.439645e-14, 5.425771e-14, 5.450338e-14, 5.436335e-14, 5.438525e-14, 
    5.425311e-14, 5.346621e-14, 5.36144e-14, 5.345742e-14, 5.347856e-14, 
    5.346909e-14, 5.335362e-14, 5.329536e-14, 5.317343e-14, 5.319558e-14, 
    5.328516e-14, 5.348807e-14, 5.341925e-14, 5.359272e-14, 5.358881e-14, 
    5.378164e-14, 5.369473e-14, 5.401844e-14, 5.392654e-14, 5.419202e-14, 
    5.412529e-14, 5.418887e-14, 5.41696e-14, 5.418913e-14, 5.409125e-14, 
    5.413319e-14, 5.404705e-14, 5.3711e-14, 5.380984e-14, 5.351481e-14, 
    5.333703e-14, 5.321896e-14, 5.313507e-14, 5.314693e-14, 5.316953e-14, 
    5.328568e-14, 5.339484e-14, 5.347795e-14, 5.353351e-14, 5.358824e-14, 
    5.375365e-14, 5.384122e-14, 5.403699e-14, 5.400172e-14, 5.40615e-14, 
    5.411865e-14, 5.421448e-14, 5.419872e-14, 5.424091e-14, 5.405995e-14, 
    5.418023e-14, 5.398164e-14, 5.403596e-14, 5.360295e-14, 5.343783e-14, 
    5.336745e-14, 5.330593e-14, 5.315605e-14, 5.325956e-14, 5.321876e-14, 
    5.331585e-14, 5.337748e-14, 5.334701e-14, 5.353503e-14, 5.346195e-14, 
    5.384641e-14, 5.368095e-14, 5.411198e-14, 5.400896e-14, 5.413667e-14, 
    5.407153e-14, 5.418312e-14, 5.408269e-14, 5.425663e-14, 5.429445e-14, 
    5.42686e-14, 5.436793e-14, 5.407712e-14, 5.418886e-14, 5.334615e-14, 
    5.335112e-14, 5.337428e-14, 5.327241e-14, 5.326619e-14, 5.317282e-14, 
    5.325592e-14, 5.329127e-14, 5.338107e-14, 5.343412e-14, 5.348454e-14, 
    5.359535e-14, 5.371897e-14, 5.389169e-14, 5.401564e-14, 5.409868e-14, 
    5.404778e-14, 5.409272e-14, 5.404247e-14, 5.401893e-14, 5.428027e-14, 
    5.413357e-14, 5.435365e-14, 5.434149e-14, 5.424191e-14, 5.434286e-14, 
    5.335461e-14, 5.332601e-14, 5.32266e-14, 5.33044e-14, 5.316264e-14, 
    5.324199e-14, 5.328758e-14, 5.346345e-14, 5.35021e-14, 5.353788e-14, 
    5.360855e-14, 5.369918e-14, 5.3858e-14, 5.399604e-14, 5.412198e-14, 
    5.411276e-14, 5.4116e-14, 5.41441e-14, 5.407446e-14, 5.415554e-14, 
    5.416912e-14, 5.413357e-14, 5.433986e-14, 5.428096e-14, 5.434123e-14, 
    5.430289e-14, 5.333531e-14, 5.338344e-14, 5.335743e-14, 5.340633e-14, 
    5.337186e-14, 5.352497e-14, 5.357084e-14, 5.378532e-14, 5.369739e-14, 
    5.383736e-14, 5.371162e-14, 5.37339e-14, 5.384186e-14, 5.371843e-14, 
    5.398843e-14, 5.380537e-14, 5.41452e-14, 5.396257e-14, 5.415663e-14, 
    5.412143e-14, 5.417972e-14, 5.423188e-14, 5.429751e-14, 5.441847e-14, 
    5.439048e-14, 5.449159e-14, 5.345518e-14, 5.351753e-14, 5.351207e-14, 
    5.357732e-14, 5.362555e-14, 5.373007e-14, 5.389749e-14, 5.383457e-14, 
    5.39501e-14, 5.397327e-14, 5.379776e-14, 5.390552e-14, 5.355927e-14, 
    5.361524e-14, 5.358194e-14, 5.346007e-14, 5.384903e-14, 5.364954e-14, 
    5.401768e-14, 5.390982e-14, 5.422444e-14, 5.406802e-14, 5.437506e-14, 
    5.450601e-14, 5.462929e-14, 5.477304e-14, 5.355158e-14, 5.350922e-14, 
    5.358509e-14, 5.368993e-14, 5.378721e-14, 5.39164e-14, 5.392963e-14, 
    5.39538e-14, 5.401641e-14, 5.406904e-14, 5.396141e-14, 5.408224e-14, 
    5.362815e-14, 5.386635e-14, 5.349318e-14, 5.360561e-14, 5.368376e-14, 
    5.364952e-14, 5.382738e-14, 5.386926e-14, 5.403925e-14, 5.395143e-14, 
    5.447367e-14, 5.424285e-14, 5.488249e-14, 5.470403e-14, 5.349441e-14, 
    5.355145e-14, 5.374974e-14, 5.365544e-14, 5.392503e-14, 5.39913e-14, 
    5.404514e-14, 5.411392e-14, 5.412137e-14, 5.416211e-14, 5.409534e-14, 
    5.415949e-14, 5.391667e-14, 5.402522e-14, 5.372713e-14, 5.379973e-14, 
    5.376634e-14, 5.372969e-14, 5.384278e-14, 5.39631e-14, 5.396572e-14, 
    5.400424e-14, 5.411272e-14, 5.392613e-14, 5.450334e-14, 5.414705e-14, 
    5.361362e-14, 5.37233e-14, 5.373902e-14, 5.369654e-14, 5.398466e-14, 
    5.388032e-14, 5.416113e-14, 5.408529e-14, 5.420953e-14, 5.414781e-14, 
    5.413872e-14, 5.405941e-14, 5.400999e-14, 5.38851e-14, 5.378339e-14, 
    5.370271e-14, 5.372148e-14, 5.381009e-14, 5.397047e-14, 5.412202e-14, 
    5.408882e-14, 5.42001e-14, 5.39055e-14, 5.402906e-14, 5.398132e-14, 
    5.410583e-14, 5.383288e-14, 5.406519e-14, 5.377342e-14, 5.379904e-14, 
    5.387825e-14, 5.403741e-14, 5.407268e-14, 5.411023e-14, 5.408707e-14, 
    5.397455e-14, 5.395612e-14, 5.387634e-14, 5.385428e-14, 5.379346e-14, 
    5.374307e-14, 5.37891e-14, 5.383741e-14, 5.397462e-14, 5.409808e-14, 
    5.423262e-14, 5.426554e-14, 5.44224e-14, 5.429465e-14, 5.450531e-14, 
    5.432612e-14, 5.46362e-14, 5.407871e-14, 5.432096e-14, 5.388187e-14, 
    5.392926e-14, 5.401484e-14, 5.421111e-14, 5.410525e-14, 5.422908e-14, 
    5.395541e-14, 5.381312e-14, 5.377635e-14, 5.37076e-14, 5.377792e-14, 
    5.37722e-14, 5.383945e-14, 5.381785e-14, 5.397917e-14, 5.389254e-14, 
    5.413848e-14, 5.422811e-14, 5.448098e-14, 5.463573e-14, 5.479314e-14, 
    5.486254e-14, 5.488367e-14, 5.489249e-14 ;

 LITR3C_vr =
  0.0005537658, 0.0005537653, 0.0005537654, 0.0005537649, 0.0005537652, 
    0.0005537649, 0.0005537657, 0.0005537652, 0.0005537656, 0.0005537658, 
    0.0005537641, 0.0005537649, 0.0005537632, 0.0005537637, 0.0005537624, 
    0.0005537632, 0.0005537622, 0.0005537624, 0.0005537617, 0.000553762, 
    0.0005537611, 0.0005537617, 0.0005537607, 0.0005537613, 0.0005537612, 
    0.0005537617, 0.0005537648, 0.0005537642, 0.0005537648, 0.0005537647, 
    0.0005537647, 0.0005537652, 0.0005537654, 0.0005537659, 0.0005537658, 
    0.0005537655, 0.0005537646, 0.0005537649, 0.0005537642, 0.0005537643, 
    0.0005537635, 0.0005537638, 0.0005537626, 0.0005537629, 0.0005537619, 
    0.0005537622, 0.000553762, 0.000553762, 0.000553762, 0.0005537623, 
    0.0005537621, 0.0005537625, 0.0005537638, 0.0005537634, 0.0005537645, 
    0.0005537652, 0.0005537657, 0.000553766, 0.000553766, 0.0005537659, 
    0.0005537655, 0.000553765, 0.0005537647, 0.0005537645, 0.0005537643, 
    0.0005537636, 0.0005537633, 0.0005537625, 0.0005537627, 0.0005537624, 
    0.0005537622, 0.0005537618, 0.0005537619, 0.0005537617, 0.0005537624, 
    0.000553762, 0.0005537627, 0.0005537625, 0.0005537642, 0.0005537649, 
    0.0005537651, 0.0005537653, 0.0005537659, 0.0005537655, 0.0005537657, 
    0.0005537653, 0.0005537651, 0.0005537652, 0.0005537645, 0.0005537648, 
    0.0005537632, 0.0005537639, 0.0005537622, 0.0005537627, 0.0005537621, 
    0.0005537624, 0.000553762, 0.0005537624, 0.0005537617, 0.0005537616, 
    0.0005537616, 0.0005537613, 0.0005537624, 0.000553762, 0.0005537652, 
    0.0005537652, 0.0005537651, 0.0005537655, 0.0005537655, 0.0005537659, 
    0.0005537656, 0.0005537654, 0.000553765, 0.0005537649, 0.0005537646, 
    0.0005537642, 0.0005537638, 0.0005537631, 0.0005537626, 0.0005537623, 
    0.0005537625, 0.0005537623, 0.0005537625, 0.0005537626, 0.0005537616, 
    0.0005537621, 0.0005537613, 0.0005537614, 0.0005537617, 0.0005537613, 
    0.0005537652, 0.0005537653, 0.0005537657, 0.0005537653, 0.0005537659, 
    0.0005537656, 0.0005537655, 0.0005537648, 0.0005537646, 0.0005537645, 
    0.0005537642, 0.0005537638, 0.0005537632, 0.0005537627, 0.0005537622, 
    0.0005537622, 0.0005537622, 0.0005537621, 0.0005537624, 0.0005537621, 
    0.000553762, 0.0005537621, 0.0005537614, 0.0005537616, 0.0005537614, 
    0.0005537615, 0.0005537652, 0.000553765, 0.0005537652, 0.000553765, 
    0.0005537651, 0.0005537645, 0.0005537643, 0.0005537635, 0.0005537638, 
    0.0005537633, 0.0005537638, 0.0005537637, 0.0005537633, 0.0005537638, 
    0.0005537627, 0.0005537634, 0.0005537621, 0.0005537628, 0.0005537621, 
    0.0005537622, 0.000553762, 0.0005537618, 0.0005537615, 0.000553761, 
    0.0005537611, 0.0005537608, 0.0005537648, 0.0005537645, 0.0005537646, 
    0.0005537643, 0.0005537641, 0.0005537637, 0.0005537631, 0.0005537633, 
    0.0005537629, 0.0005537628, 0.0005537635, 0.000553763, 0.0005537644, 
    0.0005537642, 0.0005537643, 0.0005537648, 0.0005537632, 0.000553764, 
    0.0005537626, 0.000553763, 0.0005537618, 0.0005537624, 0.0005537612, 
    0.0005537607, 0.0005537602, 0.0005537597, 0.0005537644, 0.0005537646, 
    0.0005537643, 0.0005537639, 0.0005537635, 0.000553763, 0.0005537629, 
    0.0005537628, 0.0005537626, 0.0005537624, 0.0005537628, 0.0005537624, 
    0.0005537641, 0.0005537632, 0.0005537646, 0.0005537642, 0.0005537639, 
    0.0005537641, 0.0005537634, 0.0005537632, 0.0005537625, 0.0005537628, 
    0.0005537609, 0.0005537617, 0.0005537593, 0.0005537599, 0.0005537646, 
    0.0005537644, 0.0005537636, 0.000553764, 0.0005537629, 0.0005537627, 
    0.0005537625, 0.0005537622, 0.0005537622, 0.000553762, 0.0005537623, 
    0.0005537621, 0.000553763, 0.0005537626, 0.0005537637, 0.0005537635, 
    0.0005537636, 0.0005537637, 0.0005537633, 0.0005537628, 0.0005537628, 
    0.0005537627, 0.0005537622, 0.0005537629, 0.0005537607, 0.0005537621, 
    0.0005537642, 0.0005537638, 0.0005537637, 0.0005537638, 0.0005537627, 
    0.0005537631, 0.000553762, 0.0005537624, 0.0005537618, 0.0005537621, 
    0.0005537621, 0.0005537624, 0.0005537627, 0.0005537631, 0.0005537635, 
    0.0005537638, 0.0005537638, 0.0005537634, 0.0005537628, 0.0005537622, 
    0.0005537623, 0.0005537619, 0.000553763, 0.0005537625, 0.0005537627, 
    0.0005537622, 0.0005537633, 0.0005537624, 0.0005537635, 0.0005537635, 
    0.0005537631, 0.0005537625, 0.0005537624, 0.0005537622, 0.0005537623, 
    0.0005537628, 0.0005537628, 0.0005537631, 0.0005537632, 0.0005537635, 
    0.0005537636, 0.0005537635, 0.0005537633, 0.0005537628, 0.0005537623, 
    0.0005537618, 0.0005537617, 0.000553761, 0.0005537616, 0.0005537607, 
    0.0005537614, 0.0005537602, 0.0005537624, 0.0005537614, 0.0005537631, 
    0.0005537629, 0.0005537626, 0.0005537618, 0.0005537622, 0.0005537618, 
    0.0005537628, 0.0005537634, 0.0005537635, 0.0005537638, 0.0005537635, 
    0.0005537635, 0.0005537633, 0.0005537634, 0.0005537628, 0.0005537631, 
    0.0005537621, 0.0005537618, 0.0005537608, 0.0005537602, 0.0005537596, 
    0.0005537593, 0.0005537592, 0.0005537592,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342132e-07, 1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 
    1.34213e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342128e-07, 1.34213e-07, 1.342126e-07, 1.342127e-07, 1.342124e-07, 
    1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 1.342123e-07, 
    1.342121e-07, 1.342122e-07, 1.34212e-07, 1.342121e-07, 1.342121e-07, 
    1.342122e-07, 1.34213e-07, 1.342128e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342127e-07, 1.342124e-07, 1.342125e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 
    1.342123e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 1.342129e-07, 
    1.342131e-07, 1.342132e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 
    1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 1.342124e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342124e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342128e-07, 1.34213e-07, 
    1.342131e-07, 1.342131e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342131e-07, 1.342129e-07, 1.34213e-07, 
    1.342126e-07, 1.342128e-07, 1.342124e-07, 1.342125e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 1.342122e-07, 
    1.342122e-07, 1.342121e-07, 1.342124e-07, 1.342123e-07, 1.342131e-07, 
    1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342124e-07, 1.342124e-07, 1.342124e-07, 1.342122e-07, 
    1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342123e-07, 
    1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.342122e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 
    1.342131e-07, 1.342129e-07, 1.342129e-07, 1.342127e-07, 1.342127e-07, 
    1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 
    1.342125e-07, 1.342126e-07, 1.342123e-07, 1.342125e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342121e-07, 
    1.342121e-07, 1.34212e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342126e-07, 
    1.342125e-07, 1.342125e-07, 1.342127e-07, 1.342125e-07, 1.342129e-07, 
    1.342128e-07, 1.342129e-07, 1.34213e-07, 1.342126e-07, 1.342128e-07, 
    1.342124e-07, 1.342125e-07, 1.342122e-07, 1.342124e-07, 1.342121e-07, 
    1.34212e-07, 1.342119e-07, 1.342117e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342124e-07, 1.342125e-07, 1.342124e-07, 
    1.342128e-07, 1.342126e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 
    1.34212e-07, 1.342122e-07, 1.342116e-07, 1.342118e-07, 1.342129e-07, 
    1.342129e-07, 1.342127e-07, 1.342128e-07, 1.342125e-07, 1.342125e-07, 
    1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342125e-07, 1.34212e-07, 1.342123e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342125e-07, 
    1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 1.342123e-07, 
    1.342123e-07, 1.342124e-07, 1.342125e-07, 1.342126e-07, 1.342127e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342125e-07, 
    1.342124e-07, 1.342126e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342124e-07, 1.342124e-07, 
    1.342125e-07, 1.342125e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342124e-07, 
    1.342122e-07, 1.342122e-07, 1.342121e-07, 1.342122e-07, 1.34212e-07, 
    1.342122e-07, 1.342119e-07, 1.342124e-07, 1.342122e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 
    1.342125e-07, 1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 
    1.342123e-07, 1.342122e-07, 1.34212e-07, 1.342119e-07, 1.342117e-07, 
    1.342116e-07, 1.342116e-07, 1.342116e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -6.4949e-26, 3.676358e-26, -4.166539e-26, 1.347998e-26, -5.146902e-26, 
    -6.73999e-26, -5.637083e-26, -1.274471e-25, 1.960724e-26, -2.818541e-26, 
    -1.02938e-25, -9.926167e-26, 1.225453e-25, -9.558531e-26, -3.063632e-26, 
    0, 6.617445e-26, -1.213198e-25, -3.798904e-26, 6.004719e-26, 
    1.225453e-26, 8.700715e-26, 3.308722e-26, -1.360253e-25, -4.043994e-26, 
    6.73999e-26, 6.127264e-27, -1.102908e-26, -9.068351e-26, 1.960724e-26, 
    -6.73999e-26, 4.41163e-26, 1.041635e-25, -1.053889e-25, 2.818541e-26, 
    9.068351e-26, -1.960724e-26, 7.475262e-26, -1.176435e-25, 4.289085e-26, 
    4.41163e-26, 3.676358e-27, 1.225453e-27, -3.431268e-26, -8.578169e-27, 
    -1.066144e-25, 1.225453e-27, 2.32836e-26, 8.82326e-26, -5.269447e-26, 
    2.205815e-26, 9.558531e-26, -6.127264e-26, 1.838179e-26, -1.629852e-25, 
    -6.127264e-27, 9.313441e-26, 7.842898e-26, 3.186177e-26, 5.882173e-26, 
    -4.779266e-26, 1.066144e-25, 3.431268e-26, 4.41163e-26, -6.73999e-26, 
    -7.352717e-27, 1.838179e-26, 2.450906e-27, 1.593089e-26, 2.573451e-26, 
    8.333079e-26, 4.901811e-26, -1.225453e-27, -5.269447e-26, -2.695996e-26, 
    1.262216e-25, 8.578169e-27, -2.450906e-27, 3.186177e-26, -1.02938e-25, 
    6.4949e-26, 3.186177e-26, -7.597807e-26, 2.450906e-27, 3.798904e-26, 
    1.470543e-26, -7.230172e-26, -2.205815e-26, 1.102908e-26, -1.225453e-26, 
    -1.102908e-26, -7.352717e-27, -3.186177e-26, -6.004719e-26, 6.862535e-26, 
    -2.941087e-26, -3.063632e-26, 6.617445e-26, 6.372354e-26, -5.024356e-26, 
    7.352717e-27, 8.578169e-26, 0, 4.901811e-27, -1.838179e-26, 
    -1.617598e-25, 7.597807e-26, 4.534175e-26, 4.65672e-26, 1.188689e-25, 
    2.573451e-26, 3.798904e-26, -6.004719e-26, 3.308722e-26, -4.901811e-27, 
    8.333079e-26, -9.803622e-27, 9.926167e-26, 7.352717e-27, -6.127264e-26, 
    -9.681077e-26, 1.960724e-26, 3.676358e-26, 4.901811e-27, 5.024356e-26, 
    1.078398e-25, 6.249809e-26, -2.941087e-26, 1.593089e-26, -7.230172e-26, 
    6.004719e-26, -7.597807e-26, -2.32836e-26, -1.017126e-25, -8.210533e-26, 
    -4.289085e-26, 1.090653e-25, 4.779266e-26, -1.715634e-26, -1.617598e-25, 
    -7.352717e-27, 1.960724e-26, -3.063632e-26, 7.352717e-27, -5.269447e-26, 
    -3.308722e-26, 6.004719e-26, -2.818541e-26, -5.514538e-26, -1.421525e-25, 
    7.652491e-42, 2.573451e-26, -9.803622e-27, -7.230172e-26, -1.017126e-25, 
    -1.041635e-25, 1.323489e-25, 1.225453e-26, -8.578169e-27, 3.308722e-26, 
    -5.024356e-26, -8.087988e-26, 4.534175e-26, -7.475262e-26, 2.573451e-26, 
    1.29898e-25, 3.553813e-26, -1.151926e-25, 2.08327e-26, -6.127264e-27, 
    1.16418e-25, -1.225453e-27, -9.803622e-27, 5.146902e-26, -8.087988e-26, 
    4.166539e-26, -4.534175e-26, -2.695996e-26, 6.98508e-26, 8.578169e-26, 
    -1.225453e-27, 4.779266e-26, 1.102908e-25, -8.945805e-26, 6.862535e-26, 
    1.960724e-26, 1.470543e-26, 5.269447e-26, 2.08327e-26, -5.269447e-26, 
    -1.960724e-26, -2.573451e-26, 3.553813e-26, 5.024356e-26, 7.107626e-26, 
    1.102908e-25, 9.803622e-26, -2.32836e-26, -3.431268e-26, 4.779266e-26, 
    6.73999e-26, -1.066144e-25, -3.063632e-26, 5.391992e-26, 4.65672e-26, 
    -4.41163e-26, -2.450906e-27, -2.450905e-26, -6.4949e-26, 1.715634e-26, 
    7.965443e-26, -1.262216e-25, -5.269447e-26, 2.08327e-26, 1.225453e-26, 
    1.078398e-25, 2.08327e-26, -9.803622e-27, -2.818541e-26, -9.803622e-27, 
    -8.087988e-26, 4.779266e-26, 8.333079e-26, 4.901811e-27, -3.676358e-27, 
    -5.269447e-26, 7.842898e-26, 3.431268e-26, 1.727888e-25, -1.151926e-25, 
    9.803622e-26, -6.73999e-26, -1.838179e-26, -3.921449e-26, 9.803622e-27, 
    4.901811e-26, -4.65672e-26, -2.941087e-26, -5.637083e-26, 4.534175e-26, 
    -4.043994e-26, -6.73999e-26, -2.08327e-26, 4.166539e-26, 8.578169e-27, 
    1.838179e-26, 1.960724e-26, 4.901811e-27, 7.352717e-26, 5.024356e-26, 
    3.676358e-26, -4.779266e-26, -1.372507e-25, -7.720352e-26, -2.818541e-26, 
    1.102908e-25, -8.700715e-26, -3.063632e-26, -3.553813e-26, -2.450906e-27, 
    8.578169e-27, -1.16418e-25, 4.534175e-26, 1.470543e-26, 4.534175e-26, 
    3.676358e-27, -1.29898e-25, -8.82326e-26, 9.313441e-26, 1.960724e-26, 
    4.779266e-26, -9.926167e-26, -6.862535e-26, 1.262216e-25, 1.225453e-27, 
    -9.803622e-26, 1.02938e-25, 3.063632e-26, 1.960724e-26, -2.941087e-26, 
    9.681077e-26, -9.803622e-27, 6.127264e-27, -5.024356e-26, 1.115162e-25, 
    1.225453e-27, 8.210533e-26, -1.421525e-25, -2.32836e-26, 7.107626e-26, 0, 
    2.450906e-27, -4.289085e-26, 3.308722e-26, 1.960724e-26, -1.225453e-27, 
    -4.41163e-26, 8.578169e-27, -1.066144e-25, 7.965443e-26, -1.102908e-25, 
    8.700715e-26, -2.450905e-26, -1.078398e-25, -1.225453e-27, 2.450906e-27, 
    -8.333079e-26, 6.617445e-26, -2.450905e-26, 4.901811e-26, 8.578169e-27, 
    4.779266e-26, -1.017126e-25, -6.127264e-27, -2.08327e-26, -6.98508e-26, 
    6.249809e-26, 2.695996e-26, -1.470543e-26, 2.450906e-27, 5.882173e-26, 
    5.391992e-26, 8.82326e-26, -3.431268e-26, -2.695996e-26, -2.573451e-26, 
    -1.715634e-26, 7.597807e-26, 2.450906e-27, 1.347998e-25, -3.431268e-26, 
    -7.597807e-26, -3.063632e-26, 3.676358e-27, -7.842898e-26, -4.043994e-26, 
    1.090653e-25, 5.759628e-26,
  1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 
    1.338123e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338121e-32, 1.338123e-32, 1.338119e-32, 1.33812e-32, 1.338117e-32, 
    1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338115e-32, 1.338116e-32, 
    1.338114e-32, 1.338115e-32, 1.338113e-32, 1.338114e-32, 1.338114e-32, 
    1.338115e-32, 1.338123e-32, 1.338121e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338118e-32, 1.338118e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338117e-32, 
    1.338116e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 
    1.338124e-32, 1.338125e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338117e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.338121e-32, 1.338123e-32, 
    1.338124e-32, 1.338124e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338119e-32, 1.338121e-32, 1.338117e-32, 1.338118e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 1.338115e-32, 
    1.338115e-32, 1.338114e-32, 1.338117e-32, 1.338116e-32, 1.338124e-32, 
    1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338115e-32, 
    1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338126e-32, 
    1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338116e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338115e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 
    1.338124e-32, 1.338122e-32, 1.338122e-32, 1.33812e-32, 1.33812e-32, 
    1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.33812e-32, 
    1.338118e-32, 1.338119e-32, 1.338116e-32, 1.338118e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338114e-32, 
    1.338114e-32, 1.338113e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338119e-32, 
    1.338118e-32, 1.338118e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 
    1.338121e-32, 1.338122e-32, 1.338123e-32, 1.338119e-32, 1.338121e-32, 
    1.338118e-32, 1.338119e-32, 1.338115e-32, 1.338117e-32, 1.338114e-32, 
    1.338113e-32, 1.338112e-32, 1.33811e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338117e-32, 1.338118e-32, 1.338117e-32, 
    1.338121e-32, 1.338119e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338113e-32, 1.338115e-32, 1.338109e-32, 1.338111e-32, 1.338122e-32, 
    1.338122e-32, 1.33812e-32, 1.338121e-32, 1.338118e-32, 1.338118e-32, 
    1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338116e-32, 1.338117e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338118e-32, 1.338113e-32, 1.338116e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338118e-32, 
    1.338119e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.338118e-32, 1.338119e-32, 1.33812e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338117e-32, 1.338119e-32, 1.338117e-32, 1.33812e-32, 1.33812e-32, 
    1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 
    1.338118e-32, 1.338118e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338115e-32, 1.338115e-32, 1.338114e-32, 1.338115e-32, 1.338113e-32, 
    1.338115e-32, 1.338112e-32, 1.338117e-32, 1.338115e-32, 1.338119e-32, 
    1.338118e-32, 1.338118e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 
    1.338118e-32, 1.338119e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 
    1.338116e-32, 1.338115e-32, 1.338113e-32, 1.338112e-32, 1.33811e-32, 
    1.33811e-32, 1.338109e-32, 1.338109e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.472067e-15, 1.476056e-15, 1.475282e-15, 1.478496e-15, 1.476714e-15, 
    1.478818e-15, 1.472877e-15, 1.476214e-15, 1.474084e-15, 1.472427e-15, 
    1.484726e-15, 1.47864e-15, 1.491043e-15, 1.487168e-15, 1.496895e-15, 
    1.490439e-15, 1.498196e-15, 1.49671e-15, 1.501183e-15, 1.499902e-15, 
    1.505614e-15, 1.501774e-15, 1.508574e-15, 1.504698e-15, 1.505304e-15, 
    1.501647e-15, 1.479867e-15, 1.483968e-15, 1.479623e-15, 1.480208e-15, 
    1.479946e-15, 1.47675e-15, 1.475138e-15, 1.471763e-15, 1.472376e-15, 
    1.474855e-15, 1.480472e-15, 1.478567e-15, 1.483368e-15, 1.48326e-15, 
    1.488597e-15, 1.486192e-15, 1.495151e-15, 1.492608e-15, 1.499956e-15, 
    1.498109e-15, 1.499869e-15, 1.499335e-15, 1.499876e-15, 1.497167e-15, 
    1.498327e-15, 1.495943e-15, 1.486642e-15, 1.489378e-15, 1.481212e-15, 
    1.476291e-15, 1.473023e-15, 1.470701e-15, 1.471029e-15, 1.471655e-15, 
    1.47487e-15, 1.477891e-15, 1.480191e-15, 1.481729e-15, 1.483244e-15, 
    1.487822e-15, 1.490246e-15, 1.495665e-15, 1.494689e-15, 1.496343e-15, 
    1.497925e-15, 1.500578e-15, 1.500141e-15, 1.501309e-15, 1.4963e-15, 
    1.49963e-15, 1.494133e-15, 1.495636e-15, 1.483651e-15, 1.479081e-15, 
    1.477133e-15, 1.47543e-15, 1.471282e-15, 1.474147e-15, 1.473018e-15, 
    1.475705e-15, 1.477411e-15, 1.476567e-15, 1.481771e-15, 1.479749e-15, 
    1.49039e-15, 1.48581e-15, 1.497741e-15, 1.494889e-15, 1.498424e-15, 
    1.496621e-15, 1.499709e-15, 1.49693e-15, 1.501744e-15, 1.502791e-15, 
    1.502076e-15, 1.504825e-15, 1.496776e-15, 1.499868e-15, 1.476543e-15, 
    1.476681e-15, 1.477322e-15, 1.474502e-15, 1.47433e-15, 1.471746e-15, 
    1.474046e-15, 1.475025e-15, 1.47751e-15, 1.478978e-15, 1.480374e-15, 
    1.483441e-15, 1.486863e-15, 1.491643e-15, 1.495074e-15, 1.497372e-15, 
    1.495963e-15, 1.497207e-15, 1.495817e-15, 1.495165e-15, 1.502398e-15, 
    1.498338e-15, 1.50443e-15, 1.504093e-15, 1.501337e-15, 1.504131e-15, 
    1.476777e-15, 1.475986e-15, 1.473234e-15, 1.475388e-15, 1.471464e-15, 
    1.47366e-15, 1.474922e-15, 1.47979e-15, 1.48086e-15, 1.48185e-15, 
    1.483806e-15, 1.486315e-15, 1.490711e-15, 1.494531e-15, 1.498017e-15, 
    1.497762e-15, 1.497852e-15, 1.49863e-15, 1.496702e-15, 1.498946e-15, 
    1.499322e-15, 1.498338e-15, 1.504048e-15, 1.502417e-15, 1.504086e-15, 
    1.503024e-15, 1.476243e-15, 1.477575e-15, 1.476856e-15, 1.478209e-15, 
    1.477255e-15, 1.481493e-15, 1.482763e-15, 1.488699e-15, 1.486265e-15, 
    1.49014e-15, 1.486659e-15, 1.487276e-15, 1.490264e-15, 1.486848e-15, 
    1.494321e-15, 1.489254e-15, 1.49866e-15, 1.493605e-15, 1.498976e-15, 
    1.498002e-15, 1.499616e-15, 1.501059e-15, 1.502876e-15, 1.506224e-15, 
    1.505449e-15, 1.508248e-15, 1.479561e-15, 1.481287e-15, 1.481136e-15, 
    1.482942e-15, 1.484277e-15, 1.48717e-15, 1.491804e-15, 1.490062e-15, 
    1.49326e-15, 1.493901e-15, 1.489043e-15, 1.492026e-15, 1.482442e-15, 
    1.483991e-15, 1.48307e-15, 1.479697e-15, 1.490462e-15, 1.484941e-15, 
    1.49513e-15, 1.492145e-15, 1.500853e-15, 1.496524e-15, 1.505022e-15, 
    1.508647e-15, 1.512059e-15, 1.516038e-15, 1.48223e-15, 1.481057e-15, 
    1.483157e-15, 1.486059e-15, 1.488751e-15, 1.492327e-15, 1.492693e-15, 
    1.493362e-15, 1.495095e-15, 1.496552e-15, 1.493573e-15, 1.496917e-15, 
    1.484349e-15, 1.490942e-15, 1.480613e-15, 1.483725e-15, 1.485888e-15, 
    1.48494e-15, 1.489863e-15, 1.491022e-15, 1.495728e-15, 1.493297e-15, 
    1.507752e-15, 1.501363e-15, 1.519067e-15, 1.514128e-15, 1.480647e-15, 
    1.482226e-15, 1.487714e-15, 1.485104e-15, 1.492566e-15, 1.4944e-15, 
    1.49589e-15, 1.497794e-15, 1.498e-15, 1.499128e-15, 1.49728e-15, 
    1.499055e-15, 1.492335e-15, 1.495339e-15, 1.487088e-15, 1.489098e-15, 
    1.488174e-15, 1.487159e-15, 1.490289e-15, 1.49362e-15, 1.493692e-15, 
    1.494758e-15, 1.497761e-15, 1.492596e-15, 1.508573e-15, 1.498711e-15, 
    1.483947e-15, 1.486982e-15, 1.487417e-15, 1.486242e-15, 1.494216e-15, 
    1.491329e-15, 1.499101e-15, 1.497002e-15, 1.500441e-15, 1.498732e-15, 
    1.498481e-15, 1.496285e-15, 1.494918e-15, 1.491461e-15, 1.488646e-15, 
    1.486412e-15, 1.486932e-15, 1.489385e-15, 1.493824e-15, 1.498018e-15, 
    1.4971e-15, 1.500179e-15, 1.492025e-15, 1.495445e-15, 1.494124e-15, 
    1.49757e-15, 1.490015e-15, 1.496445e-15, 1.488369e-15, 1.489079e-15, 
    1.491271e-15, 1.495676e-15, 1.496653e-15, 1.497692e-15, 1.497051e-15, 
    1.493936e-15, 1.493427e-15, 1.491218e-15, 1.490608e-15, 1.488924e-15, 
    1.48753e-15, 1.488804e-15, 1.490141e-15, 1.493938e-15, 1.497356e-15, 
    1.50108e-15, 1.501991e-15, 1.506332e-15, 1.502797e-15, 1.508627e-15, 
    1.503668e-15, 1.51225e-15, 1.49682e-15, 1.503525e-15, 1.491371e-15, 
    1.492683e-15, 1.495052e-15, 1.500484e-15, 1.497554e-15, 1.500981e-15, 
    1.493407e-15, 1.489468e-15, 1.488451e-15, 1.486548e-15, 1.488494e-15, 
    1.488336e-15, 1.490197e-15, 1.489599e-15, 1.494064e-15, 1.491667e-15, 
    1.498474e-15, 1.500955e-15, 1.507954e-15, 1.512237e-15, 1.516594e-15, 
    1.518515e-15, 1.5191e-15, 1.519344e-15 ;

 LITR3N_vr =
  7.663713e-06, 7.663706e-06, 7.663708e-06, 7.663702e-06, 7.663705e-06, 
    7.663701e-06, 7.663712e-06, 7.663706e-06, 7.66371e-06, 7.663713e-06, 
    7.663689e-06, 7.663701e-06, 7.663677e-06, 7.663684e-06, 7.663666e-06, 
    7.663678e-06, 7.663663e-06, 7.663666e-06, 7.663657e-06, 7.66366e-06, 
    7.663649e-06, 7.663656e-06, 7.663643e-06, 7.663651e-06, 7.66365e-06, 
    7.663656e-06, 7.663699e-06, 7.663691e-06, 7.663699e-06, 7.663698e-06, 
    7.663699e-06, 7.663704e-06, 7.663708e-06, 7.663714e-06, 7.663713e-06, 
    7.663709e-06, 7.663698e-06, 7.663702e-06, 7.663692e-06, 7.663692e-06, 
    7.663682e-06, 7.663686e-06, 7.663669e-06, 7.663674e-06, 7.66366e-06, 
    7.663663e-06, 7.66366e-06, 7.663661e-06, 7.66366e-06, 7.663665e-06, 
    7.663663e-06, 7.663668e-06, 7.663685e-06, 7.663681e-06, 7.663696e-06, 
    7.663705e-06, 7.663712e-06, 7.663716e-06, 7.663716e-06, 7.663714e-06, 
    7.663708e-06, 7.663702e-06, 7.663698e-06, 7.663695e-06, 7.663692e-06, 
    7.663683e-06, 7.663679e-06, 7.663668e-06, 7.66367e-06, 7.663667e-06, 
    7.663663e-06, 7.663659e-06, 7.66366e-06, 7.663657e-06, 7.663667e-06, 
    7.663661e-06, 7.663671e-06, 7.663668e-06, 7.663692e-06, 7.663701e-06, 
    7.663704e-06, 7.663707e-06, 7.663715e-06, 7.66371e-06, 7.663712e-06, 
    7.663707e-06, 7.663703e-06, 7.663705e-06, 7.663695e-06, 7.663699e-06, 
    7.663678e-06, 7.663687e-06, 7.663664e-06, 7.66367e-06, 7.663662e-06, 
    7.663666e-06, 7.663661e-06, 7.663665e-06, 7.663656e-06, 7.663654e-06, 
    7.663656e-06, 7.663651e-06, 7.663666e-06, 7.66366e-06, 7.663705e-06, 
    7.663705e-06, 7.663703e-06, 7.663709e-06, 7.66371e-06, 7.663714e-06, 
    7.66371e-06, 7.663708e-06, 7.663703e-06, 7.663701e-06, 7.663698e-06, 
    7.663692e-06, 7.663685e-06, 7.663676e-06, 7.663669e-06, 7.663665e-06, 
    7.663668e-06, 7.663665e-06, 7.663668e-06, 7.663669e-06, 7.663655e-06, 
    7.663662e-06, 7.663652e-06, 7.663652e-06, 7.663657e-06, 7.663652e-06, 
    7.663704e-06, 7.663706e-06, 7.663712e-06, 7.663707e-06, 7.663715e-06, 
    7.663711e-06, 7.663708e-06, 7.663699e-06, 7.663697e-06, 7.663695e-06, 
    7.663691e-06, 7.663686e-06, 7.663678e-06, 7.663671e-06, 7.663663e-06, 
    7.663664e-06, 7.663664e-06, 7.663662e-06, 7.663666e-06, 7.663662e-06, 
    7.663661e-06, 7.663662e-06, 7.663652e-06, 7.663655e-06, 7.663652e-06, 
    7.663654e-06, 7.663706e-06, 7.663703e-06, 7.663704e-06, 7.663702e-06, 
    7.663703e-06, 7.663695e-06, 7.663693e-06, 7.663682e-06, 7.663686e-06, 
    7.663679e-06, 7.663685e-06, 7.663684e-06, 7.663679e-06, 7.663685e-06, 
    7.663671e-06, 7.663681e-06, 7.663662e-06, 7.663672e-06, 7.663662e-06, 
    7.663663e-06, 7.663661e-06, 7.663658e-06, 7.663654e-06, 7.663648e-06, 
    7.663649e-06, 7.663643e-06, 7.663699e-06, 7.663696e-06, 7.663696e-06, 
    7.663692e-06, 7.66369e-06, 7.663684e-06, 7.663675e-06, 7.663679e-06, 
    7.663672e-06, 7.663672e-06, 7.663681e-06, 7.663675e-06, 7.663693e-06, 
    7.663691e-06, 7.663692e-06, 7.663699e-06, 7.663678e-06, 7.663689e-06, 
    7.663669e-06, 7.663675e-06, 7.663658e-06, 7.663666e-06, 7.66365e-06, 
    7.663643e-06, 7.663636e-06, 7.663629e-06, 7.663694e-06, 7.663696e-06, 
    7.663692e-06, 7.663687e-06, 7.663682e-06, 7.663674e-06, 7.663674e-06, 
    7.663672e-06, 7.663669e-06, 7.663666e-06, 7.663672e-06, 7.663666e-06, 
    7.66369e-06, 7.663677e-06, 7.663697e-06, 7.663692e-06, 7.663687e-06, 
    7.663689e-06, 7.66368e-06, 7.663677e-06, 7.663668e-06, 7.663672e-06, 
    7.663644e-06, 7.663657e-06, 7.663622e-06, 7.663632e-06, 7.663697e-06, 
    7.663694e-06, 7.663683e-06, 7.663689e-06, 7.663674e-06, 7.663671e-06, 
    7.663668e-06, 7.663664e-06, 7.663663e-06, 7.663662e-06, 7.663665e-06, 
    7.663662e-06, 7.663674e-06, 7.663669e-06, 7.663684e-06, 7.663681e-06, 
    7.663682e-06, 7.663684e-06, 7.663679e-06, 7.663672e-06, 7.663672e-06, 
    7.66367e-06, 7.663664e-06, 7.663674e-06, 7.663643e-06, 7.663662e-06, 
    7.663691e-06, 7.663685e-06, 7.663684e-06, 7.663686e-06, 7.663671e-06, 
    7.663676e-06, 7.663662e-06, 7.663665e-06, 7.663659e-06, 7.663662e-06, 
    7.663662e-06, 7.663667e-06, 7.66367e-06, 7.663676e-06, 7.663682e-06, 
    7.663686e-06, 7.663685e-06, 7.663681e-06, 7.663672e-06, 7.663663e-06, 
    7.663665e-06, 7.66366e-06, 7.663675e-06, 7.663669e-06, 7.663671e-06, 
    7.663664e-06, 7.663679e-06, 7.663667e-06, 7.663682e-06, 7.663681e-06, 
    7.663677e-06, 7.663668e-06, 7.663666e-06, 7.663664e-06, 7.663665e-06, 
    7.663672e-06, 7.663672e-06, 7.663677e-06, 7.663678e-06, 7.663682e-06, 
    7.663684e-06, 7.663682e-06, 7.663679e-06, 7.663672e-06, 7.663665e-06, 
    7.663658e-06, 7.663656e-06, 7.663647e-06, 7.663654e-06, 7.663643e-06, 
    7.663652e-06, 7.663636e-06, 7.663666e-06, 7.663652e-06, 7.663676e-06, 
    7.663674e-06, 7.663669e-06, 7.663659e-06, 7.663664e-06, 7.663658e-06, 
    7.663672e-06, 7.66368e-06, 7.663682e-06, 7.663686e-06, 7.663682e-06, 
    7.663682e-06, 7.663679e-06, 7.66368e-06, 7.663672e-06, 7.663676e-06, 
    7.663662e-06, 7.663658e-06, 7.663644e-06, 7.663636e-06, 7.663628e-06, 
    7.663624e-06, 7.663622e-06, 7.663622e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.318442e-14, 5.332856e-14, 5.330056e-14, 5.341671e-14, 5.33523e-14, 
    5.342833e-14, 5.321368e-14, 5.333426e-14, 5.32573e-14, 5.319743e-14, 
    5.364177e-14, 5.342189e-14, 5.387e-14, 5.373001e-14, 5.408143e-14, 
    5.38482e-14, 5.412843e-14, 5.407476e-14, 5.423635e-14, 5.419008e-14, 
    5.439645e-14, 5.425771e-14, 5.450338e-14, 5.436335e-14, 5.438525e-14, 
    5.425311e-14, 5.346621e-14, 5.36144e-14, 5.345742e-14, 5.347856e-14, 
    5.346909e-14, 5.335362e-14, 5.329536e-14, 5.317343e-14, 5.319558e-14, 
    5.328516e-14, 5.348807e-14, 5.341925e-14, 5.359272e-14, 5.358881e-14, 
    5.378164e-14, 5.369473e-14, 5.401844e-14, 5.392654e-14, 5.419202e-14, 
    5.412529e-14, 5.418887e-14, 5.41696e-14, 5.418913e-14, 5.409125e-14, 
    5.413319e-14, 5.404705e-14, 5.3711e-14, 5.380984e-14, 5.351481e-14, 
    5.333703e-14, 5.321896e-14, 5.313507e-14, 5.314693e-14, 5.316953e-14, 
    5.328568e-14, 5.339484e-14, 5.347795e-14, 5.353351e-14, 5.358824e-14, 
    5.375365e-14, 5.384122e-14, 5.403699e-14, 5.400172e-14, 5.40615e-14, 
    5.411865e-14, 5.421448e-14, 5.419872e-14, 5.424091e-14, 5.405995e-14, 
    5.418023e-14, 5.398164e-14, 5.403596e-14, 5.360295e-14, 5.343783e-14, 
    5.336745e-14, 5.330593e-14, 5.315605e-14, 5.325956e-14, 5.321876e-14, 
    5.331585e-14, 5.337748e-14, 5.334701e-14, 5.353503e-14, 5.346195e-14, 
    5.384641e-14, 5.368095e-14, 5.411198e-14, 5.400896e-14, 5.413667e-14, 
    5.407153e-14, 5.418312e-14, 5.408269e-14, 5.425663e-14, 5.429445e-14, 
    5.42686e-14, 5.436793e-14, 5.407712e-14, 5.418886e-14, 5.334615e-14, 
    5.335112e-14, 5.337428e-14, 5.327241e-14, 5.326619e-14, 5.317282e-14, 
    5.325592e-14, 5.329127e-14, 5.338107e-14, 5.343412e-14, 5.348454e-14, 
    5.359535e-14, 5.371897e-14, 5.389169e-14, 5.401564e-14, 5.409868e-14, 
    5.404778e-14, 5.409272e-14, 5.404247e-14, 5.401893e-14, 5.428027e-14, 
    5.413357e-14, 5.435365e-14, 5.434149e-14, 5.424191e-14, 5.434286e-14, 
    5.335461e-14, 5.332601e-14, 5.32266e-14, 5.33044e-14, 5.316264e-14, 
    5.324199e-14, 5.328758e-14, 5.346345e-14, 5.35021e-14, 5.353788e-14, 
    5.360855e-14, 5.369918e-14, 5.3858e-14, 5.399604e-14, 5.412198e-14, 
    5.411276e-14, 5.4116e-14, 5.41441e-14, 5.407446e-14, 5.415554e-14, 
    5.416912e-14, 5.413357e-14, 5.433986e-14, 5.428096e-14, 5.434123e-14, 
    5.430289e-14, 5.333531e-14, 5.338344e-14, 5.335743e-14, 5.340633e-14, 
    5.337186e-14, 5.352497e-14, 5.357084e-14, 5.378532e-14, 5.369739e-14, 
    5.383736e-14, 5.371162e-14, 5.37339e-14, 5.384186e-14, 5.371843e-14, 
    5.398843e-14, 5.380537e-14, 5.41452e-14, 5.396257e-14, 5.415663e-14, 
    5.412143e-14, 5.417972e-14, 5.423188e-14, 5.429751e-14, 5.441847e-14, 
    5.439048e-14, 5.449159e-14, 5.345518e-14, 5.351753e-14, 5.351207e-14, 
    5.357732e-14, 5.362555e-14, 5.373007e-14, 5.389749e-14, 5.383457e-14, 
    5.39501e-14, 5.397327e-14, 5.379776e-14, 5.390552e-14, 5.355927e-14, 
    5.361524e-14, 5.358194e-14, 5.346007e-14, 5.384903e-14, 5.364954e-14, 
    5.401768e-14, 5.390982e-14, 5.422444e-14, 5.406802e-14, 5.437506e-14, 
    5.450601e-14, 5.462929e-14, 5.477304e-14, 5.355158e-14, 5.350922e-14, 
    5.358509e-14, 5.368993e-14, 5.378721e-14, 5.39164e-14, 5.392963e-14, 
    5.39538e-14, 5.401641e-14, 5.406904e-14, 5.396141e-14, 5.408224e-14, 
    5.362815e-14, 5.386635e-14, 5.349318e-14, 5.360561e-14, 5.368376e-14, 
    5.364952e-14, 5.382738e-14, 5.386926e-14, 5.403925e-14, 5.395143e-14, 
    5.447367e-14, 5.424285e-14, 5.488249e-14, 5.470403e-14, 5.349441e-14, 
    5.355145e-14, 5.374974e-14, 5.365544e-14, 5.392503e-14, 5.39913e-14, 
    5.404514e-14, 5.411392e-14, 5.412137e-14, 5.416211e-14, 5.409534e-14, 
    5.415949e-14, 5.391667e-14, 5.402522e-14, 5.372713e-14, 5.379973e-14, 
    5.376634e-14, 5.372969e-14, 5.384278e-14, 5.39631e-14, 5.396572e-14, 
    5.400424e-14, 5.411272e-14, 5.392613e-14, 5.450334e-14, 5.414705e-14, 
    5.361362e-14, 5.37233e-14, 5.373902e-14, 5.369654e-14, 5.398466e-14, 
    5.388032e-14, 5.416113e-14, 5.408529e-14, 5.420953e-14, 5.414781e-14, 
    5.413872e-14, 5.405941e-14, 5.400999e-14, 5.38851e-14, 5.378339e-14, 
    5.370271e-14, 5.372148e-14, 5.381009e-14, 5.397047e-14, 5.412202e-14, 
    5.408882e-14, 5.42001e-14, 5.39055e-14, 5.402906e-14, 5.398132e-14, 
    5.410583e-14, 5.383288e-14, 5.406519e-14, 5.377342e-14, 5.379904e-14, 
    5.387825e-14, 5.403741e-14, 5.407268e-14, 5.411023e-14, 5.408707e-14, 
    5.397455e-14, 5.395612e-14, 5.387634e-14, 5.385428e-14, 5.379346e-14, 
    5.374307e-14, 5.37891e-14, 5.383741e-14, 5.397462e-14, 5.409808e-14, 
    5.423262e-14, 5.426554e-14, 5.44224e-14, 5.429465e-14, 5.450531e-14, 
    5.432612e-14, 5.46362e-14, 5.407871e-14, 5.432096e-14, 5.388187e-14, 
    5.392926e-14, 5.401484e-14, 5.421111e-14, 5.410525e-14, 5.422908e-14, 
    5.395541e-14, 5.381312e-14, 5.377635e-14, 5.37076e-14, 5.377792e-14, 
    5.37722e-14, 5.383945e-14, 5.381785e-14, 5.397917e-14, 5.389254e-14, 
    5.413848e-14, 5.422811e-14, 5.448098e-14, 5.463573e-14, 5.479314e-14, 
    5.486254e-14, 5.488367e-14, 5.489249e-14 ;

 LITTERC =
  5.976208e-05, 5.976193e-05, 5.976196e-05, 5.976184e-05, 5.976191e-05, 
    5.976183e-05, 5.976205e-05, 5.976193e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976184e-05, 5.976138e-05, 5.976153e-05, 5.976117e-05, 
    5.976141e-05, 5.976112e-05, 5.976118e-05, 5.976101e-05, 5.976106e-05, 
    5.976085e-05, 5.976099e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976179e-05, 5.976164e-05, 5.97618e-05, 5.976178e-05, 
    5.976179e-05, 5.976191e-05, 5.976197e-05, 5.976209e-05, 5.976207e-05, 
    5.976198e-05, 5.976177e-05, 5.976184e-05, 5.976166e-05, 5.976167e-05, 
    5.976147e-05, 5.976156e-05, 5.976123e-05, 5.976133e-05, 5.976106e-05, 
    5.976113e-05, 5.976106e-05, 5.976108e-05, 5.976106e-05, 5.976116e-05, 
    5.976112e-05, 5.976121e-05, 5.976154e-05, 5.976145e-05, 5.976174e-05, 
    5.976192e-05, 5.976204e-05, 5.976213e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976178e-05, 5.976172e-05, 5.976167e-05, 
    5.97615e-05, 5.976141e-05, 5.976121e-05, 5.976125e-05, 5.976119e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.976101e-05, 5.976119e-05, 
    5.976107e-05, 5.976127e-05, 5.976122e-05, 5.976165e-05, 5.976182e-05, 
    5.976189e-05, 5.976195e-05, 5.976211e-05, 5.9762e-05, 5.976204e-05, 
    5.976194e-05, 5.976188e-05, 5.976191e-05, 5.976172e-05, 5.976179e-05, 
    5.976141e-05, 5.976157e-05, 5.976114e-05, 5.976124e-05, 5.976111e-05, 
    5.976118e-05, 5.976107e-05, 5.976117e-05, 5.976099e-05, 5.976095e-05, 
    5.976098e-05, 5.976088e-05, 5.976117e-05, 5.976106e-05, 5.976191e-05, 
    5.976191e-05, 5.976189e-05, 5.976199e-05, 5.976199e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976188e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976154e-05, 5.976136e-05, 5.976123e-05, 5.976115e-05, 
    5.97612e-05, 5.976116e-05, 5.976121e-05, 5.976123e-05, 5.976097e-05, 
    5.976111e-05, 5.976089e-05, 5.976091e-05, 5.976101e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.97621e-05, 
    5.976202e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976172e-05, 
    5.976165e-05, 5.976155e-05, 5.976139e-05, 5.976126e-05, 5.976113e-05, 
    5.976114e-05, 5.976113e-05, 5.97611e-05, 5.976118e-05, 5.976109e-05, 
    5.976108e-05, 5.976111e-05, 5.976091e-05, 5.976097e-05, 5.976091e-05, 
    5.976094e-05, 5.976193e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976189e-05, 5.976173e-05, 5.976169e-05, 5.976147e-05, 5.976156e-05, 
    5.976142e-05, 5.976154e-05, 5.976152e-05, 5.976141e-05, 5.976154e-05, 
    5.976126e-05, 5.976145e-05, 5.97611e-05, 5.976129e-05, 5.976109e-05, 
    5.976113e-05, 5.976107e-05, 5.976102e-05, 5.976095e-05, 5.976083e-05, 
    5.976086e-05, 5.976075e-05, 5.97618e-05, 5.976174e-05, 5.976174e-05, 
    5.976168e-05, 5.976163e-05, 5.976153e-05, 5.976135e-05, 5.976142e-05, 
    5.97613e-05, 5.976128e-05, 5.976146e-05, 5.976135e-05, 5.97617e-05, 
    5.976164e-05, 5.976167e-05, 5.97618e-05, 5.976141e-05, 5.976161e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976074e-05, 5.976061e-05, 5.976047e-05, 5.97617e-05, 5.976175e-05, 
    5.976167e-05, 5.976157e-05, 5.976147e-05, 5.976134e-05, 5.976132e-05, 
    5.97613e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976117e-05, 
    5.976163e-05, 5.976139e-05, 5.976177e-05, 5.976165e-05, 5.976157e-05, 
    5.976161e-05, 5.976143e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976077e-05, 5.976101e-05, 5.976036e-05, 5.976054e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.97616e-05, 5.976133e-05, 5.976126e-05, 
    5.976121e-05, 5.976114e-05, 5.976113e-05, 5.976109e-05, 5.976115e-05, 
    5.976109e-05, 5.976134e-05, 5.976123e-05, 5.976153e-05, 5.976145e-05, 
    5.976149e-05, 5.976153e-05, 5.976141e-05, 5.976129e-05, 5.976129e-05, 
    5.976125e-05, 5.976114e-05, 5.976133e-05, 5.976074e-05, 5.97611e-05, 
    5.976164e-05, 5.976153e-05, 5.976151e-05, 5.976156e-05, 5.976127e-05, 
    5.976137e-05, 5.976109e-05, 5.976117e-05, 5.976104e-05, 5.97611e-05, 
    5.976111e-05, 5.976119e-05, 5.976124e-05, 5.976137e-05, 5.976147e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976128e-05, 5.976113e-05, 
    5.976116e-05, 5.976105e-05, 5.976135e-05, 5.976122e-05, 5.976127e-05, 
    5.976114e-05, 5.976142e-05, 5.976118e-05, 5.976148e-05, 5.976146e-05, 
    5.976137e-05, 5.976121e-05, 5.976118e-05, 5.976114e-05, 5.976116e-05, 
    5.976128e-05, 5.97613e-05, 5.976138e-05, 5.97614e-05, 5.976146e-05, 
    5.976151e-05, 5.976146e-05, 5.976142e-05, 5.976128e-05, 5.976115e-05, 
    5.976102e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976074e-05, 
    5.976092e-05, 5.976061e-05, 5.976117e-05, 5.976093e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976104e-05, 5.976114e-05, 5.976102e-05, 
    5.97613e-05, 5.976144e-05, 5.976148e-05, 5.976155e-05, 5.976147e-05, 
    5.976148e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976136e-05, 
    5.976111e-05, 5.976102e-05, 5.976076e-05, 5.976061e-05, 5.976045e-05, 
    5.976038e-05, 5.976036e-05, 5.976035e-05 ;

 LITTERC_HR =
  8.580827e-13, 8.604064e-13, 8.599551e-13, 8.618275e-13, 8.607893e-13, 
    8.620149e-13, 8.585544e-13, 8.604983e-13, 8.592577e-13, 8.582925e-13, 
    8.654558e-13, 8.619111e-13, 8.691352e-13, 8.668784e-13, 8.725437e-13, 
    8.687836e-13, 8.733013e-13, 8.724361e-13, 8.750411e-13, 8.742953e-13, 
    8.77622e-13, 8.753853e-13, 8.793459e-13, 8.770885e-13, 8.774415e-13, 
    8.753114e-13, 8.626257e-13, 8.650145e-13, 8.624839e-13, 8.628247e-13, 
    8.62672e-13, 8.608104e-13, 8.598713e-13, 8.579055e-13, 8.582627e-13, 
    8.597067e-13, 8.62978e-13, 8.618686e-13, 8.646651e-13, 8.64602e-13, 
    8.677107e-13, 8.663096e-13, 8.715281e-13, 8.700467e-13, 8.743264e-13, 
    8.732506e-13, 8.742757e-13, 8.739651e-13, 8.742798e-13, 8.727019e-13, 
    8.73378e-13, 8.719893e-13, 8.665719e-13, 8.681653e-13, 8.634091e-13, 
    8.605431e-13, 8.586395e-13, 8.572872e-13, 8.574784e-13, 8.578427e-13, 
    8.597151e-13, 8.614749e-13, 8.628148e-13, 8.637106e-13, 8.645929e-13, 
    8.672594e-13, 8.686712e-13, 8.718272e-13, 8.712586e-13, 8.722224e-13, 
    8.731436e-13, 8.746886e-13, 8.744345e-13, 8.751147e-13, 8.721974e-13, 
    8.741364e-13, 8.70935e-13, 8.718107e-13, 8.6483e-13, 8.621681e-13, 
    8.610334e-13, 8.600417e-13, 8.576253e-13, 8.592942e-13, 8.586364e-13, 
    8.602016e-13, 8.611951e-13, 8.607039e-13, 8.637351e-13, 8.62557e-13, 
    8.687549e-13, 8.660874e-13, 8.730362e-13, 8.713754e-13, 8.734342e-13, 
    8.72384e-13, 8.741829e-13, 8.72564e-13, 8.75368e-13, 8.759778e-13, 
    8.75561e-13, 8.771624e-13, 8.724741e-13, 8.742755e-13, 8.6069e-13, 
    8.607701e-13, 8.611436e-13, 8.595013e-13, 8.594009e-13, 8.578956e-13, 
    8.592354e-13, 8.598054e-13, 8.61253e-13, 8.621082e-13, 8.629211e-13, 
    8.647075e-13, 8.667004e-13, 8.694849e-13, 8.714831e-13, 8.728217e-13, 
    8.720011e-13, 8.727256e-13, 8.719156e-13, 8.71536e-13, 8.757491e-13, 
    8.733842e-13, 8.769321e-13, 8.76736e-13, 8.751308e-13, 8.767581e-13, 
    8.608264e-13, 8.603653e-13, 8.587627e-13, 8.60017e-13, 8.577317e-13, 
    8.590108e-13, 8.597458e-13, 8.625811e-13, 8.632041e-13, 8.637809e-13, 
    8.649203e-13, 8.663813e-13, 8.689417e-13, 8.711671e-13, 8.731973e-13, 
    8.730487e-13, 8.73101e-13, 8.735541e-13, 8.724313e-13, 8.737383e-13, 
    8.739573e-13, 8.733842e-13, 8.767098e-13, 8.757602e-13, 8.767318e-13, 
    8.761137e-13, 8.605153e-13, 8.612912e-13, 8.608719e-13, 8.616601e-13, 
    8.611046e-13, 8.635729e-13, 8.643124e-13, 8.677701e-13, 8.663524e-13, 
    8.686091e-13, 8.66582e-13, 8.669411e-13, 8.686814e-13, 8.666917e-13, 
    8.710443e-13, 8.680933e-13, 8.735717e-13, 8.706275e-13, 8.73756e-13, 
    8.731886e-13, 8.741282e-13, 8.749692e-13, 8.760271e-13, 8.77977e-13, 
    8.775258e-13, 8.791559e-13, 8.624476e-13, 8.634529e-13, 8.633649e-13, 
    8.644169e-13, 8.651944e-13, 8.668793e-13, 8.695784e-13, 8.68564e-13, 
    8.704265e-13, 8.708e-13, 8.679706e-13, 8.697077e-13, 8.641258e-13, 
    8.650281e-13, 8.644913e-13, 8.625267e-13, 8.687971e-13, 8.65581e-13, 
    8.71516e-13, 8.697771e-13, 8.748492e-13, 8.723274e-13, 8.772771e-13, 
    8.793883e-13, 8.813757e-13, 8.836929e-13, 8.640019e-13, 8.63319e-13, 
    8.645421e-13, 8.662322e-13, 8.678005e-13, 8.698832e-13, 8.700964e-13, 
    8.704861e-13, 8.714955e-13, 8.72344e-13, 8.706088e-13, 8.725566e-13, 
    8.652363e-13, 8.690762e-13, 8.630603e-13, 8.648729e-13, 8.661328e-13, 
    8.655807e-13, 8.684481e-13, 8.691232e-13, 8.718637e-13, 8.70448e-13, 
    8.78867e-13, 8.751459e-13, 8.854573e-13, 8.825805e-13, 8.630802e-13, 
    8.639998e-13, 8.671964e-13, 8.656761e-13, 8.700224e-13, 8.710906e-13, 
    8.719586e-13, 8.730675e-13, 8.731875e-13, 8.738443e-13, 8.727679e-13, 
    8.73802e-13, 8.698875e-13, 8.716375e-13, 8.668319e-13, 8.680023e-13, 
    8.674641e-13, 8.668733e-13, 8.686963e-13, 8.70636e-13, 8.706783e-13, 
    8.712993e-13, 8.730481e-13, 8.700399e-13, 8.793452e-13, 8.736015e-13, 
    8.65002e-13, 8.667702e-13, 8.670236e-13, 8.663388e-13, 8.709835e-13, 
    8.693016e-13, 8.738284e-13, 8.726059e-13, 8.746088e-13, 8.736137e-13, 
    8.734672e-13, 8.721886e-13, 8.713919e-13, 8.693786e-13, 8.677389e-13, 
    8.664382e-13, 8.667408e-13, 8.681694e-13, 8.707548e-13, 8.731981e-13, 
    8.726628e-13, 8.744566e-13, 8.697075e-13, 8.716995e-13, 8.709298e-13, 
    8.72937e-13, 8.685368e-13, 8.722818e-13, 8.675781e-13, 8.679911e-13, 
    8.692682e-13, 8.71834e-13, 8.724025e-13, 8.73008e-13, 8.726346e-13, 
    8.708206e-13, 8.705235e-13, 8.692374e-13, 8.688817e-13, 8.679013e-13, 
    8.670888e-13, 8.678309e-13, 8.686098e-13, 8.708217e-13, 8.728121e-13, 
    8.74981e-13, 8.755117e-13, 8.780403e-13, 8.75981e-13, 8.79377e-13, 
    8.764883e-13, 8.814871e-13, 8.724998e-13, 8.764051e-13, 8.693266e-13, 
    8.700905e-13, 8.714702e-13, 8.746343e-13, 8.729275e-13, 8.749238e-13, 
    8.70512e-13, 8.682182e-13, 8.676254e-13, 8.665172e-13, 8.676507e-13, 
    8.675586e-13, 8.686427e-13, 8.682944e-13, 8.708951e-13, 8.694985e-13, 
    8.734633e-13, 8.749083e-13, 8.789848e-13, 8.814794e-13, 8.84017e-13, 
    8.851359e-13, 8.854764e-13, 8.856186e-13 ;

 LITTERC_LOSS =
  1.58916e-12, 1.593464e-12, 1.592628e-12, 1.596096e-12, 1.594173e-12, 
    1.596442e-12, 1.590034e-12, 1.593634e-12, 1.591336e-12, 1.589549e-12, 
    1.602815e-12, 1.59625e-12, 1.609629e-12, 1.60545e-12, 1.615942e-12, 
    1.608978e-12, 1.617345e-12, 1.615743e-12, 1.620567e-12, 1.619186e-12, 
    1.625347e-12, 1.621205e-12, 1.62854e-12, 1.624359e-12, 1.625013e-12, 
    1.621068e-12, 1.597574e-12, 1.601998e-12, 1.597311e-12, 1.597942e-12, 
    1.59766e-12, 1.594212e-12, 1.592473e-12, 1.588832e-12, 1.589493e-12, 
    1.592168e-12, 1.598226e-12, 1.596172e-12, 1.601351e-12, 1.601234e-12, 
    1.606991e-12, 1.604396e-12, 1.614061e-12, 1.611318e-12, 1.619244e-12, 
    1.617251e-12, 1.61915e-12, 1.618574e-12, 1.619157e-12, 1.616235e-12, 
    1.617487e-12, 1.614915e-12, 1.604882e-12, 1.607833e-12, 1.599025e-12, 
    1.593717e-12, 1.590191e-12, 1.587687e-12, 1.588041e-12, 1.588716e-12, 
    1.592183e-12, 1.595443e-12, 1.597924e-12, 1.599583e-12, 1.601217e-12, 
    1.606156e-12, 1.60877e-12, 1.614615e-12, 1.613562e-12, 1.615347e-12, 
    1.617053e-12, 1.619914e-12, 1.619444e-12, 1.620704e-12, 1.615301e-12, 
    1.618892e-12, 1.612963e-12, 1.614584e-12, 1.601656e-12, 1.596726e-12, 
    1.594625e-12, 1.592788e-12, 1.588313e-12, 1.591404e-12, 1.590185e-12, 
    1.593084e-12, 1.594924e-12, 1.594015e-12, 1.599628e-12, 1.597447e-12, 
    1.608925e-12, 1.603985e-12, 1.616854e-12, 1.613778e-12, 1.617591e-12, 
    1.615646e-12, 1.618978e-12, 1.61598e-12, 1.621173e-12, 1.622302e-12, 
    1.62153e-12, 1.624496e-12, 1.615813e-12, 1.619149e-12, 1.593989e-12, 
    1.594137e-12, 1.594829e-12, 1.591787e-12, 1.591602e-12, 1.588814e-12, 
    1.591295e-12, 1.59235e-12, 1.595031e-12, 1.596615e-12, 1.598121e-12, 
    1.601429e-12, 1.60512e-12, 1.610277e-12, 1.613978e-12, 1.616457e-12, 
    1.614937e-12, 1.616279e-12, 1.614779e-12, 1.614076e-12, 1.621879e-12, 
    1.617499e-12, 1.624069e-12, 1.623706e-12, 1.620733e-12, 1.623747e-12, 
    1.594241e-12, 1.593387e-12, 1.59042e-12, 1.592742e-12, 1.58851e-12, 
    1.590879e-12, 1.59224e-12, 1.597491e-12, 1.598645e-12, 1.599713e-12, 
    1.601823e-12, 1.604529e-12, 1.609271e-12, 1.613392e-12, 1.617153e-12, 
    1.616877e-12, 1.616974e-12, 1.617813e-12, 1.615734e-12, 1.618155e-12, 
    1.61856e-12, 1.617499e-12, 1.623658e-12, 1.621899e-12, 1.623699e-12, 
    1.622554e-12, 1.593665e-12, 1.595102e-12, 1.594326e-12, 1.595785e-12, 
    1.594757e-12, 1.599328e-12, 1.600697e-12, 1.607101e-12, 1.604476e-12, 
    1.608655e-12, 1.604901e-12, 1.605566e-12, 1.608789e-12, 1.605104e-12, 
    1.613165e-12, 1.6077e-12, 1.617846e-12, 1.612393e-12, 1.618187e-12, 
    1.617136e-12, 1.618877e-12, 1.620434e-12, 1.622393e-12, 1.626005e-12, 
    1.625169e-12, 1.628188e-12, 1.597244e-12, 1.599106e-12, 1.598943e-12, 
    1.600891e-12, 1.602331e-12, 1.605451e-12, 1.61045e-12, 1.608571e-12, 
    1.612021e-12, 1.612713e-12, 1.607473e-12, 1.61069e-12, 1.600352e-12, 
    1.602023e-12, 1.601029e-12, 1.59739e-12, 1.609003e-12, 1.603047e-12, 
    1.614039e-12, 1.610818e-12, 1.620212e-12, 1.615541e-12, 1.624709e-12, 
    1.628618e-12, 1.632299e-12, 1.636591e-12, 1.600122e-12, 1.598858e-12, 
    1.601123e-12, 1.604253e-12, 1.607158e-12, 1.611015e-12, 1.61141e-12, 
    1.612131e-12, 1.614001e-12, 1.615572e-12, 1.612359e-12, 1.615966e-12, 
    1.602409e-12, 1.60952e-12, 1.598379e-12, 1.601736e-12, 1.604069e-12, 
    1.603047e-12, 1.608357e-12, 1.609607e-12, 1.614683e-12, 1.612061e-12, 
    1.627653e-12, 1.620761e-12, 1.639858e-12, 1.634531e-12, 1.598416e-12, 
    1.600119e-12, 1.606039e-12, 1.603223e-12, 1.611273e-12, 1.613251e-12, 
    1.614859e-12, 1.616912e-12, 1.617134e-12, 1.618351e-12, 1.616357e-12, 
    1.618272e-12, 1.611023e-12, 1.614264e-12, 1.605364e-12, 1.607531e-12, 
    1.606535e-12, 1.60544e-12, 1.608817e-12, 1.612409e-12, 1.612487e-12, 
    1.613637e-12, 1.616876e-12, 1.611305e-12, 1.628539e-12, 1.617901e-12, 
    1.601975e-12, 1.605249e-12, 1.605719e-12, 1.604451e-12, 1.613053e-12, 
    1.609938e-12, 1.618321e-12, 1.616057e-12, 1.619767e-12, 1.617924e-12, 
    1.617652e-12, 1.615284e-12, 1.613809e-12, 1.61008e-12, 1.607043e-12, 
    1.604635e-12, 1.605195e-12, 1.607841e-12, 1.612629e-12, 1.617154e-12, 
    1.616163e-12, 1.619485e-12, 1.610689e-12, 1.614378e-12, 1.612953e-12, 
    1.61667e-12, 1.608521e-12, 1.615457e-12, 1.606746e-12, 1.607511e-12, 
    1.609876e-12, 1.614628e-12, 1.615681e-12, 1.616802e-12, 1.61611e-12, 
    1.612751e-12, 1.612201e-12, 1.609819e-12, 1.60916e-12, 1.607344e-12, 
    1.60584e-12, 1.607214e-12, 1.608656e-12, 1.612753e-12, 1.616439e-12, 
    1.620456e-12, 1.621439e-12, 1.626122e-12, 1.622308e-12, 1.628597e-12, 
    1.623248e-12, 1.632505e-12, 1.615861e-12, 1.623093e-12, 1.609984e-12, 
    1.611399e-12, 1.613954e-12, 1.619814e-12, 1.616653e-12, 1.62035e-12, 
    1.612179e-12, 1.607931e-12, 1.606833e-12, 1.604781e-12, 1.60688e-12, 
    1.606709e-12, 1.608717e-12, 1.608072e-12, 1.612889e-12, 1.610302e-12, 
    1.617645e-12, 1.620321e-12, 1.627871e-12, 1.632491e-12, 1.637191e-12, 
    1.639263e-12, 1.639894e-12, 1.640157e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  3.916364e-18, 3.91493e-18, 3.915202e-18, 3.914062e-18, 3.914684e-18, 
    3.913945e-18, 3.916061e-18, 3.914884e-18, 3.915628e-18, 3.916218e-18, 
    3.911888e-18, 3.914007e-18, 3.909577e-18, 3.910943e-18, 3.907479e-18, 
    3.909805e-18, 3.907005e-18, 3.907518e-18, 3.905909e-18, 3.906368e-18, 
    3.90437e-18, 3.905697e-18, 3.903292e-18, 3.904672e-18, 3.904467e-18, 
    3.905745e-18, 3.913554e-18, 3.91216e-18, 3.913643e-18, 3.913443e-18, 
    3.913527e-18, 3.914681e-18, 3.915281e-18, 3.916455e-18, 3.916237e-18, 
    3.915364e-18, 3.913352e-18, 3.914016e-18, 3.91229e-18, 3.912328e-18, 
    3.910429e-18, 3.911285e-18, 3.908077e-18, 3.908982e-18, 3.906348e-18, 
    3.907014e-18, 3.906384e-18, 3.906572e-18, 3.906382e-18, 3.907356e-18, 
    3.90694e-18, 3.90779e-18, 3.91113e-18, 3.910156e-18, 3.913079e-18, 
    3.914882e-18, 3.916014e-18, 3.916839e-18, 3.916723e-18, 3.916506e-18, 
    3.915359e-18, 3.91426e-18, 3.91343e-18, 3.91288e-18, 3.912334e-18, 
    3.910756e-18, 3.909861e-18, 3.907908e-18, 3.908237e-18, 3.907662e-18, 
    3.907079e-18, 3.906133e-18, 3.906286e-18, 3.905874e-18, 3.90766e-18, 
    3.906481e-18, 3.90843e-18, 3.9079e-18, 3.912278e-18, 3.913833e-18, 
    3.914574e-18, 3.915153e-18, 3.916635e-18, 3.915617e-18, 3.91602e-18, 
    3.915041e-18, 3.914432e-18, 3.914729e-18, 3.912865e-18, 3.913593e-18, 
    3.909809e-18, 3.911436e-18, 3.907147e-18, 3.908167e-18, 3.906899e-18, 
    3.907542e-18, 3.906449e-18, 3.907432e-18, 3.905714e-18, 3.905351e-18, 
    3.905601e-18, 3.90461e-18, 3.907489e-18, 3.906393e-18, 3.914742e-18, 
    3.914694e-18, 3.914461e-18, 3.915491e-18, 3.915549e-18, 3.916466e-18, 
    3.915641e-18, 3.915298e-18, 3.91439e-18, 3.913871e-18, 3.913371e-18, 
    3.912273e-18, 3.911063e-18, 3.909348e-18, 3.908102e-18, 3.907273e-18, 
    3.907775e-18, 3.907333e-18, 3.907831e-18, 3.908061e-18, 3.905493e-18, 
    3.906942e-18, 3.904753e-18, 3.90487e-18, 3.905868e-18, 3.904857e-18, 
    3.91466e-18, 3.914938e-18, 3.915935e-18, 3.915155e-18, 3.916565e-18, 
    3.915787e-18, 3.915346e-18, 3.913598e-18, 3.913192e-18, 3.912844e-18, 
    3.912137e-18, 3.911242e-18, 3.909679e-18, 3.908306e-18, 3.907042e-18, 
    3.907132e-18, 3.907101e-18, 3.906828e-18, 3.907517e-18, 3.906714e-18, 
    3.906589e-18, 3.906931e-18, 3.904887e-18, 3.905469e-18, 3.904873e-18, 
    3.90525e-18, 3.914845e-18, 3.914372e-18, 3.914629e-18, 3.914151e-18, 
    3.914495e-18, 3.912993e-18, 3.912543e-18, 3.910415e-18, 3.911264e-18, 
    3.909888e-18, 3.911118e-18, 3.910905e-18, 3.909881e-18, 3.911045e-18, 
    3.908399e-18, 3.910226e-18, 3.906818e-18, 3.908676e-18, 3.906703e-18, 
    3.907047e-18, 3.906469e-18, 3.905962e-18, 3.905307e-18, 3.904127e-18, 
    3.904396e-18, 3.903395e-18, 3.913659e-18, 3.913055e-18, 3.913091e-18, 
    3.912447e-18, 3.911975e-18, 3.910931e-18, 3.90928e-18, 3.909895e-18, 
    3.908747e-18, 3.908522e-18, 3.910256e-18, 3.909208e-18, 3.912638e-18, 
    3.912101e-18, 3.912408e-18, 3.913621e-18, 3.909777e-18, 3.911758e-18, 
    3.908085e-18, 3.909153e-18, 3.906037e-18, 3.907602e-18, 3.904548e-18, 
    3.90329e-18, 3.902028e-18, 3.900648e-18, 3.912707e-18, 3.913119e-18, 
    3.912365e-18, 3.911356e-18, 3.910371e-18, 3.909091e-18, 3.908951e-18, 
    3.908716e-18, 3.908087e-18, 3.907568e-18, 3.908659e-18, 3.907436e-18, 
    3.91201e-18, 3.909597e-18, 3.913291e-18, 3.9122e-18, 3.911408e-18, 
    3.911738e-18, 3.909961e-18, 3.909548e-18, 3.90788e-18, 3.908732e-18, 
    3.903616e-18, 3.905879e-18, 3.899542e-18, 3.90132e-18, 3.913267e-18, 
    3.9127e-18, 3.910754e-18, 3.911677e-18, 3.908997e-18, 3.908346e-18, 
    3.907801e-18, 3.907135e-18, 3.90705e-18, 3.906654e-18, 3.907306e-18, 
    3.906673e-18, 3.909088e-18, 3.908005e-18, 3.910955e-18, 3.910247e-18, 
    3.910567e-18, 3.910931e-18, 3.90981e-18, 3.908646e-18, 3.908593e-18, 
    3.908225e-18, 3.907237e-18, 3.908985e-18, 3.903375e-18, 3.906883e-18, 
    3.912084e-18, 3.911031e-18, 3.910847e-18, 3.911261e-18, 3.908412e-18, 
    3.909447e-18, 3.906659e-18, 3.907406e-18, 3.906176e-18, 3.906789e-18, 
    3.906881e-18, 3.907663e-18, 3.908158e-18, 3.909404e-18, 3.910412e-18, 
    3.911197e-18, 3.911012e-18, 3.910149e-18, 3.908568e-18, 3.907055e-18, 
    3.90739e-18, 3.906269e-18, 3.909191e-18, 3.907979e-18, 3.908457e-18, 
    3.907207e-18, 3.909917e-18, 3.907693e-18, 3.910496e-18, 3.910244e-18, 
    3.909467e-18, 3.907916e-18, 3.907531e-18, 3.907172e-18, 3.907388e-18, 
    3.908523e-18, 3.908697e-18, 3.909479e-18, 3.909709e-18, 3.910297e-18, 
    3.910797e-18, 3.910347e-18, 3.90988e-18, 3.908511e-18, 3.907294e-18, 
    3.905959e-18, 3.905621e-18, 3.904134e-18, 3.905382e-18, 3.903361e-18, 
    3.905136e-18, 3.902036e-18, 3.907523e-18, 3.905133e-18, 3.909422e-18, 
    3.908952e-18, 3.908133e-18, 3.906197e-18, 3.907212e-18, 3.906012e-18, 
    3.908701e-18, 3.910133e-18, 3.910469e-18, 3.911154e-18, 3.910454e-18, 
    3.91051e-18, 3.909842e-18, 3.910055e-18, 3.908465e-18, 3.909317e-18, 
    3.906891e-18, 3.906014e-18, 3.90351e-18, 3.901995e-18, 3.900411e-18, 
    3.899728e-18, 3.899517e-18, 3.899431e-18 ;

 MEG_acetic_acid =
  5.874546e-19, 5.872395e-19, 5.872803e-19, 5.871092e-19, 5.872026e-19, 
    5.870917e-19, 5.874091e-19, 5.872326e-19, 5.873442e-19, 5.874328e-19, 
    5.867831e-19, 5.871011e-19, 5.864365e-19, 5.866415e-19, 5.861218e-19, 
    5.864707e-19, 5.860508e-19, 5.861277e-19, 5.858863e-19, 5.859552e-19, 
    5.856555e-19, 5.858545e-19, 5.854938e-19, 5.857007e-19, 5.856699e-19, 
    5.858617e-19, 5.870331e-19, 5.86824e-19, 5.870465e-19, 5.870164e-19, 
    5.87029e-19, 5.872021e-19, 5.872921e-19, 5.874683e-19, 5.874355e-19, 
    5.873046e-19, 5.870028e-19, 5.871025e-19, 5.868435e-19, 5.868492e-19, 
    5.865643e-19, 5.866927e-19, 5.862116e-19, 5.863472e-19, 5.859523e-19, 
    5.860521e-19, 5.859576e-19, 5.859858e-19, 5.859573e-19, 5.861035e-19, 
    5.86041e-19, 5.861685e-19, 5.866695e-19, 5.865234e-19, 5.869618e-19, 
    5.872323e-19, 5.874021e-19, 5.875259e-19, 5.875084e-19, 5.874759e-19, 
    5.873039e-19, 5.871389e-19, 5.870145e-19, 5.869319e-19, 5.868501e-19, 
    5.866133e-19, 5.864792e-19, 5.861862e-19, 5.862355e-19, 5.861492e-19, 
    5.860619e-19, 5.8592e-19, 5.859428e-19, 5.858812e-19, 5.861489e-19, 
    5.859722e-19, 5.862646e-19, 5.86185e-19, 5.868417e-19, 5.870749e-19, 
    5.871861e-19, 5.87273e-19, 5.874952e-19, 5.873425e-19, 5.87403e-19, 
    5.872562e-19, 5.871649e-19, 5.872094e-19, 5.869297e-19, 5.870389e-19, 
    5.864714e-19, 5.867154e-19, 5.86072e-19, 5.862251e-19, 5.860349e-19, 
    5.861312e-19, 5.859672e-19, 5.861147e-19, 5.858571e-19, 5.858026e-19, 
    5.858402e-19, 5.856915e-19, 5.861233e-19, 5.85959e-19, 5.872113e-19, 
    5.872041e-19, 5.871691e-19, 5.873236e-19, 5.873323e-19, 5.874698e-19, 
    5.873462e-19, 5.872947e-19, 5.871585e-19, 5.870806e-19, 5.870057e-19, 
    5.86841e-19, 5.866594e-19, 5.864022e-19, 5.862154e-19, 5.86091e-19, 
    5.861663e-19, 5.860999e-19, 5.861747e-19, 5.862091e-19, 5.85824e-19, 
    5.860412e-19, 5.857129e-19, 5.857306e-19, 5.858802e-19, 5.857286e-19, 
    5.871989e-19, 5.872406e-19, 5.873903e-19, 5.872732e-19, 5.874847e-19, 
    5.87368e-19, 5.873019e-19, 5.870396e-19, 5.869787e-19, 5.869267e-19, 
    5.868206e-19, 5.866863e-19, 5.864518e-19, 5.862459e-19, 5.860562e-19, 
    5.860698e-19, 5.860651e-19, 5.860242e-19, 5.861275e-19, 5.860072e-19, 
    5.859883e-19, 5.860397e-19, 5.85733e-19, 5.858204e-19, 5.857309e-19, 
    5.857874e-19, 5.872267e-19, 5.871558e-19, 5.871943e-19, 5.871226e-19, 
    5.871742e-19, 5.869489e-19, 5.868814e-19, 5.865623e-19, 5.866896e-19, 
    5.864831e-19, 5.866676e-19, 5.866357e-19, 5.864822e-19, 5.866567e-19, 
    5.862599e-19, 5.86534e-19, 5.860227e-19, 5.863014e-19, 5.860055e-19, 
    5.860571e-19, 5.859704e-19, 5.858943e-19, 5.85796e-19, 5.85619e-19, 
    5.856594e-19, 5.855093e-19, 5.870488e-19, 5.869583e-19, 5.869636e-19, 
    5.868671e-19, 5.867962e-19, 5.866396e-19, 5.863919e-19, 5.864842e-19, 
    5.86312e-19, 5.862783e-19, 5.865384e-19, 5.863812e-19, 5.868957e-19, 
    5.868151e-19, 5.868611e-19, 5.870432e-19, 5.864665e-19, 5.867637e-19, 
    5.862128e-19, 5.863729e-19, 5.859055e-19, 5.861403e-19, 5.856822e-19, 
    5.854935e-19, 5.853042e-19, 5.850972e-19, 5.86906e-19, 5.869678e-19, 
    5.868548e-19, 5.867034e-19, 5.865557e-19, 5.863637e-19, 5.863426e-19, 
    5.863074e-19, 5.862131e-19, 5.861351e-19, 5.862988e-19, 5.861154e-19, 
    5.868016e-19, 5.864396e-19, 5.869936e-19, 5.868301e-19, 5.867112e-19, 
    5.867607e-19, 5.864941e-19, 5.864322e-19, 5.861821e-19, 5.863099e-19, 
    5.855423e-19, 5.858817e-19, 5.849313e-19, 5.851979e-19, 5.869901e-19, 
    5.86905e-19, 5.866131e-19, 5.867515e-19, 5.863495e-19, 5.862519e-19, 
    5.861702e-19, 5.860702e-19, 5.860575e-19, 5.85998e-19, 5.860959e-19, 
    5.860009e-19, 5.863633e-19, 5.862008e-19, 5.866433e-19, 5.86537e-19, 
    5.865851e-19, 5.866396e-19, 5.864715e-19, 5.862969e-19, 5.86289e-19, 
    5.862337e-19, 5.860855e-19, 5.863477e-19, 5.855062e-19, 5.860324e-19, 
    5.868125e-19, 5.866547e-19, 5.86627e-19, 5.866891e-19, 5.862618e-19, 
    5.86417e-19, 5.859989e-19, 5.861109e-19, 5.859264e-19, 5.860184e-19, 
    5.860321e-19, 5.861494e-19, 5.862237e-19, 5.864106e-19, 5.865617e-19, 
    5.866795e-19, 5.866518e-19, 5.865223e-19, 5.862852e-19, 5.860583e-19, 
    5.861085e-19, 5.859403e-19, 5.863787e-19, 5.861968e-19, 5.862685e-19, 
    5.86081e-19, 5.864875e-19, 5.861539e-19, 5.865744e-19, 5.865367e-19, 
    5.8642e-19, 5.861873e-19, 5.861297e-19, 5.860758e-19, 5.861082e-19, 
    5.862784e-19, 5.863045e-19, 5.864218e-19, 5.864563e-19, 5.865446e-19, 
    5.866196e-19, 5.865521e-19, 5.86482e-19, 5.862767e-19, 5.86094e-19, 
    5.858938e-19, 5.858432e-19, 5.8562e-19, 5.858073e-19, 5.855041e-19, 
    5.857704e-19, 5.853054e-19, 5.861284e-19, 5.8577e-19, 5.864133e-19, 
    5.863428e-19, 5.862199e-19, 5.859296e-19, 5.860819e-19, 5.859017e-19, 
    5.863052e-19, 5.8652e-19, 5.865704e-19, 5.866731e-19, 5.86568e-19, 
    5.865764e-19, 5.864762e-19, 5.865082e-19, 5.862698e-19, 5.863976e-19, 
    5.860336e-19, 5.859021e-19, 5.855264e-19, 5.852992e-19, 5.850617e-19, 
    5.849591e-19, 5.849276e-19, 5.849146e-19 ;

 MEG_acetone =
  1.220793e-16, 1.220561e-16, 1.220605e-16, 1.220421e-16, 1.220521e-16, 
    1.220402e-16, 1.220744e-16, 1.220554e-16, 1.220674e-16, 1.22077e-16, 
    1.220069e-16, 1.220412e-16, 1.219695e-16, 1.219916e-16, 1.219356e-16, 
    1.219732e-16, 1.21928e-16, 1.219362e-16, 1.219102e-16, 1.219177e-16, 
    1.218854e-16, 1.219068e-16, 1.21868e-16, 1.218903e-16, 1.21887e-16, 
    1.219076e-16, 1.220338e-16, 1.220113e-16, 1.220353e-16, 1.22032e-16, 
    1.220334e-16, 1.220521e-16, 1.220618e-16, 1.220808e-16, 1.220772e-16, 
    1.220631e-16, 1.220306e-16, 1.220413e-16, 1.220134e-16, 1.22014e-16, 
    1.219833e-16, 1.219971e-16, 1.219453e-16, 1.219599e-16, 1.219173e-16, 
    1.219281e-16, 1.219179e-16, 1.21921e-16, 1.219179e-16, 1.219336e-16, 
    1.219269e-16, 1.219406e-16, 1.219946e-16, 1.219789e-16, 1.220262e-16, 
    1.220553e-16, 1.220736e-16, 1.22087e-16, 1.220851e-16, 1.220816e-16, 
    1.22063e-16, 1.220453e-16, 1.220318e-16, 1.220229e-16, 1.220141e-16, 
    1.219886e-16, 1.219741e-16, 1.219425e-16, 1.219478e-16, 1.219386e-16, 
    1.219291e-16, 1.219139e-16, 1.219163e-16, 1.219097e-16, 1.219385e-16, 
    1.219195e-16, 1.21951e-16, 1.219424e-16, 1.220132e-16, 1.220383e-16, 
    1.220503e-16, 1.220597e-16, 1.220837e-16, 1.220672e-16, 1.220737e-16, 
    1.220579e-16, 1.220481e-16, 1.220529e-16, 1.220227e-16, 1.220345e-16, 
    1.219733e-16, 1.219996e-16, 1.219302e-16, 1.219467e-16, 1.219262e-16, 
    1.219366e-16, 1.21919e-16, 1.219348e-16, 1.219071e-16, 1.219012e-16, 
    1.219053e-16, 1.218893e-16, 1.219358e-16, 1.219181e-16, 1.220531e-16, 
    1.220523e-16, 1.220485e-16, 1.220652e-16, 1.220661e-16, 1.22081e-16, 
    1.220676e-16, 1.220621e-16, 1.220474e-16, 1.22039e-16, 1.220309e-16, 
    1.220131e-16, 1.219936e-16, 1.219658e-16, 1.219457e-16, 1.219323e-16, 
    1.219404e-16, 1.219332e-16, 1.219413e-16, 1.21945e-16, 1.219035e-16, 
    1.219269e-16, 1.218916e-16, 1.218935e-16, 1.219096e-16, 1.218933e-16, 
    1.220517e-16, 1.220562e-16, 1.220724e-16, 1.220597e-16, 1.220826e-16, 
    1.2207e-16, 1.220628e-16, 1.220346e-16, 1.22028e-16, 1.220224e-16, 
    1.220109e-16, 1.219965e-16, 1.219712e-16, 1.21949e-16, 1.219285e-16, 
    1.2193e-16, 1.219295e-16, 1.219251e-16, 1.219362e-16, 1.219233e-16, 
    1.219212e-16, 1.219268e-16, 1.218937e-16, 1.219032e-16, 1.218935e-16, 
    1.218996e-16, 1.220547e-16, 1.220471e-16, 1.220512e-16, 1.220435e-16, 
    1.220491e-16, 1.220248e-16, 1.220175e-16, 1.219831e-16, 1.219968e-16, 
    1.219745e-16, 1.219944e-16, 1.21991e-16, 1.219744e-16, 1.219933e-16, 
    1.219505e-16, 1.2198e-16, 1.219249e-16, 1.21955e-16, 1.219231e-16, 
    1.219286e-16, 1.219193e-16, 1.219111e-16, 1.219005e-16, 1.218815e-16, 
    1.218858e-16, 1.218697e-16, 1.220355e-16, 1.220258e-16, 1.220264e-16, 
    1.220159e-16, 1.220083e-16, 1.219914e-16, 1.219647e-16, 1.219747e-16, 
    1.219561e-16, 1.219525e-16, 1.219805e-16, 1.219636e-16, 1.22019e-16, 
    1.220103e-16, 1.220153e-16, 1.220349e-16, 1.219728e-16, 1.220048e-16, 
    1.219454e-16, 1.219627e-16, 1.219123e-16, 1.219376e-16, 1.218883e-16, 
    1.21868e-16, 1.218476e-16, 1.218254e-16, 1.220201e-16, 1.220268e-16, 
    1.220146e-16, 1.219983e-16, 1.219824e-16, 1.219617e-16, 1.219594e-16, 
    1.219556e-16, 1.219454e-16, 1.21937e-16, 1.219547e-16, 1.219349e-16, 
    1.220089e-16, 1.219699e-16, 1.220296e-16, 1.220119e-16, 1.219991e-16, 
    1.220045e-16, 1.219757e-16, 1.219691e-16, 1.219421e-16, 1.219559e-16, 
    1.218732e-16, 1.219097e-16, 1.218076e-16, 1.218362e-16, 1.220292e-16, 
    1.2202e-16, 1.219886e-16, 1.220035e-16, 1.219601e-16, 1.219496e-16, 
    1.219408e-16, 1.2193e-16, 1.219287e-16, 1.219223e-16, 1.219328e-16, 
    1.219226e-16, 1.219616e-16, 1.219441e-16, 1.219918e-16, 1.219804e-16, 
    1.219855e-16, 1.219914e-16, 1.219733e-16, 1.219545e-16, 1.219536e-16, 
    1.219477e-16, 1.219317e-16, 1.2196e-16, 1.218693e-16, 1.21926e-16, 
    1.220101e-16, 1.21993e-16, 1.219901e-16, 1.219968e-16, 1.219507e-16, 
    1.219674e-16, 1.219224e-16, 1.219344e-16, 1.219146e-16, 1.219245e-16, 
    1.219259e-16, 1.219386e-16, 1.219466e-16, 1.219667e-16, 1.21983e-16, 
    1.219957e-16, 1.219927e-16, 1.219788e-16, 1.219532e-16, 1.219288e-16, 
    1.219342e-16, 1.219161e-16, 1.219633e-16, 1.219437e-16, 1.219514e-16, 
    1.219312e-16, 1.21975e-16, 1.21939e-16, 1.219844e-16, 1.219803e-16, 
    1.219677e-16, 1.219427e-16, 1.219365e-16, 1.219306e-16, 1.219341e-16, 
    1.219525e-16, 1.219553e-16, 1.21968e-16, 1.219717e-16, 1.219812e-16, 
    1.219893e-16, 1.21982e-16, 1.219744e-16, 1.219523e-16, 1.219326e-16, 
    1.219111e-16, 1.219056e-16, 1.218816e-16, 1.219017e-16, 1.218691e-16, 
    1.218978e-16, 1.218478e-16, 1.219363e-16, 1.218977e-16, 1.21967e-16, 
    1.219594e-16, 1.219462e-16, 1.219149e-16, 1.219313e-16, 1.219119e-16, 
    1.219554e-16, 1.219785e-16, 1.21984e-16, 1.21995e-16, 1.219837e-16, 
    1.219846e-16, 1.219738e-16, 1.219773e-16, 1.219516e-16, 1.219653e-16, 
    1.219261e-16, 1.219119e-16, 1.218715e-16, 1.218471e-16, 1.218216e-16, 
    1.218106e-16, 1.218072e-16, 1.218058e-16 ;

 MEG_carene_3 =
  4.84213e-17, 4.841163e-17, 4.841346e-17, 4.840577e-17, 4.840996e-17, 
    4.840498e-17, 4.841926e-17, 4.841131e-17, 4.841634e-17, 4.842032e-17, 
    4.83911e-17, 4.84054e-17, 4.837552e-17, 4.838474e-17, 4.836138e-17, 
    4.837706e-17, 4.835819e-17, 4.836164e-17, 4.835081e-17, 4.83539e-17, 
    4.834044e-17, 4.834938e-17, 4.833319e-17, 4.834248e-17, 4.834109e-17, 
    4.83497e-17, 4.840234e-17, 4.839294e-17, 4.840295e-17, 4.840159e-17, 
    4.840216e-17, 4.840994e-17, 4.841399e-17, 4.842192e-17, 4.842044e-17, 
    4.841455e-17, 4.840098e-17, 4.840546e-17, 4.839382e-17, 4.839408e-17, 
    4.838127e-17, 4.838704e-17, 4.836541e-17, 4.837151e-17, 4.835377e-17, 
    4.835825e-17, 4.835401e-17, 4.835527e-17, 4.835399e-17, 4.836056e-17, 
    4.835775e-17, 4.836347e-17, 4.8386e-17, 4.837943e-17, 4.839914e-17, 
    4.84113e-17, 4.841894e-17, 4.842451e-17, 4.842372e-17, 4.842226e-17, 
    4.841452e-17, 4.84071e-17, 4.840151e-17, 4.83978e-17, 4.839412e-17, 
    4.838347e-17, 4.837744e-17, 4.836427e-17, 4.836649e-17, 4.836261e-17, 
    4.835869e-17, 4.835232e-17, 4.835334e-17, 4.835057e-17, 4.83626e-17, 
    4.835466e-17, 4.83678e-17, 4.836421e-17, 4.839374e-17, 4.840422e-17, 
    4.840922e-17, 4.841313e-17, 4.842313e-17, 4.841626e-17, 4.841898e-17, 
    4.841238e-17, 4.840827e-17, 4.841027e-17, 4.83977e-17, 4.840261e-17, 
    4.837709e-17, 4.838806e-17, 4.835914e-17, 4.836602e-17, 4.835747e-17, 
    4.83618e-17, 4.835444e-17, 4.836106e-17, 4.834949e-17, 4.834705e-17, 
    4.834873e-17, 4.834206e-17, 4.836145e-17, 4.835407e-17, 4.841036e-17, 
    4.841004e-17, 4.840846e-17, 4.841541e-17, 4.84158e-17, 4.842199e-17, 
    4.841642e-17, 4.841411e-17, 4.840798e-17, 4.840448e-17, 4.840111e-17, 
    4.839371e-17, 4.838555e-17, 4.837398e-17, 4.836558e-17, 4.835999e-17, 
    4.836338e-17, 4.836039e-17, 4.836375e-17, 4.83653e-17, 4.834801e-17, 
    4.835776e-17, 4.834302e-17, 4.834381e-17, 4.835053e-17, 4.834372e-17, 
    4.84098e-17, 4.841168e-17, 4.841841e-17, 4.841314e-17, 4.842265e-17, 
    4.841741e-17, 4.841443e-17, 4.840264e-17, 4.83999e-17, 4.839756e-17, 
    4.839279e-17, 4.838675e-17, 4.837621e-17, 4.836695e-17, 4.835843e-17, 
    4.835905e-17, 4.835883e-17, 4.8357e-17, 4.836163e-17, 4.835623e-17, 
    4.835538e-17, 4.835769e-17, 4.834393e-17, 4.834784e-17, 4.834383e-17, 
    4.834637e-17, 4.841105e-17, 4.840786e-17, 4.840959e-17, 4.840637e-17, 
    4.840869e-17, 4.839856e-17, 4.839552e-17, 4.838118e-17, 4.838691e-17, 
    4.837762e-17, 4.838591e-17, 4.838448e-17, 4.837758e-17, 4.838542e-17, 
    4.836759e-17, 4.83799e-17, 4.835693e-17, 4.836945e-17, 4.835615e-17, 
    4.835847e-17, 4.835458e-17, 4.835116e-17, 4.834675e-17, 4.833881e-17, 
    4.834062e-17, 4.833388e-17, 4.840305e-17, 4.839898e-17, 4.839922e-17, 
    4.839488e-17, 4.83917e-17, 4.838466e-17, 4.837352e-17, 4.837767e-17, 
    4.836993e-17, 4.836842e-17, 4.838011e-17, 4.837304e-17, 4.839616e-17, 
    4.839254e-17, 4.839461e-17, 4.84028e-17, 4.837687e-17, 4.839023e-17, 
    4.836547e-17, 4.837267e-17, 4.835166e-17, 4.836221e-17, 4.834164e-17, 
    4.833318e-17, 4.832469e-17, 4.831541e-17, 4.839663e-17, 4.839941e-17, 
    4.839433e-17, 4.838752e-17, 4.838088e-17, 4.837225e-17, 4.837131e-17, 
    4.836972e-17, 4.836548e-17, 4.836198e-17, 4.836933e-17, 4.836109e-17, 
    4.839193e-17, 4.837566e-17, 4.840056e-17, 4.839321e-17, 4.838787e-17, 
    4.83901e-17, 4.837811e-17, 4.837534e-17, 4.836409e-17, 4.836983e-17, 
    4.833537e-17, 4.83506e-17, 4.830798e-17, 4.831992e-17, 4.840041e-17, 
    4.839658e-17, 4.838346e-17, 4.838969e-17, 4.837161e-17, 4.836723e-17, 
    4.836355e-17, 4.835906e-17, 4.835849e-17, 4.835582e-17, 4.836021e-17, 
    4.835595e-17, 4.837223e-17, 4.836493e-17, 4.838482e-17, 4.838004e-17, 
    4.83822e-17, 4.838466e-17, 4.83771e-17, 4.836925e-17, 4.83689e-17, 
    4.836641e-17, 4.835974e-17, 4.837153e-17, 4.833374e-17, 4.835736e-17, 
    4.839243e-17, 4.838533e-17, 4.838409e-17, 4.838688e-17, 4.836767e-17, 
    4.837465e-17, 4.835586e-17, 4.836089e-17, 4.83526e-17, 4.835673e-17, 
    4.835735e-17, 4.836262e-17, 4.836596e-17, 4.837436e-17, 4.838116e-17, 
    4.838645e-17, 4.838521e-17, 4.837938e-17, 4.836872e-17, 4.835853e-17, 
    4.836078e-17, 4.835323e-17, 4.837293e-17, 4.836475e-17, 4.836797e-17, 
    4.835955e-17, 4.837782e-17, 4.836282e-17, 4.838172e-17, 4.838003e-17, 
    4.837478e-17, 4.836432e-17, 4.836173e-17, 4.835931e-17, 4.836077e-17, 
    4.836842e-17, 4.836959e-17, 4.837487e-17, 4.837642e-17, 4.838038e-17, 
    4.838376e-17, 4.838072e-17, 4.837757e-17, 4.836834e-17, 4.836013e-17, 
    4.835114e-17, 4.834887e-17, 4.833885e-17, 4.834725e-17, 4.833365e-17, 
    4.834559e-17, 4.832474e-17, 4.836167e-17, 4.834558e-17, 4.837448e-17, 
    4.837132e-17, 4.836578e-17, 4.835275e-17, 4.835959e-17, 4.83515e-17, 
    4.836962e-17, 4.837927e-17, 4.838155e-17, 4.838616e-17, 4.838144e-17, 
    4.838181e-17, 4.837731e-17, 4.837875e-17, 4.836803e-17, 4.837378e-17, 
    4.835742e-17, 4.835151e-17, 4.833465e-17, 4.832447e-17, 4.831382e-17, 
    4.830923e-17, 4.830781e-17, 4.830723e-17 ;

 MEG_ethanol =
  3.916364e-18, 3.91493e-18, 3.915202e-18, 3.914062e-18, 3.914684e-18, 
    3.913945e-18, 3.916061e-18, 3.914884e-18, 3.915628e-18, 3.916218e-18, 
    3.911888e-18, 3.914007e-18, 3.909577e-18, 3.910943e-18, 3.907479e-18, 
    3.909805e-18, 3.907005e-18, 3.907518e-18, 3.905909e-18, 3.906368e-18, 
    3.90437e-18, 3.905697e-18, 3.903292e-18, 3.904672e-18, 3.904467e-18, 
    3.905745e-18, 3.913554e-18, 3.91216e-18, 3.913643e-18, 3.913443e-18, 
    3.913527e-18, 3.914681e-18, 3.915281e-18, 3.916455e-18, 3.916237e-18, 
    3.915364e-18, 3.913352e-18, 3.914016e-18, 3.91229e-18, 3.912328e-18, 
    3.910429e-18, 3.911285e-18, 3.908077e-18, 3.908982e-18, 3.906348e-18, 
    3.907014e-18, 3.906384e-18, 3.906572e-18, 3.906382e-18, 3.907356e-18, 
    3.90694e-18, 3.90779e-18, 3.91113e-18, 3.910156e-18, 3.913079e-18, 
    3.914882e-18, 3.916014e-18, 3.916839e-18, 3.916723e-18, 3.916506e-18, 
    3.915359e-18, 3.91426e-18, 3.91343e-18, 3.91288e-18, 3.912334e-18, 
    3.910756e-18, 3.909861e-18, 3.907908e-18, 3.908237e-18, 3.907662e-18, 
    3.907079e-18, 3.906133e-18, 3.906286e-18, 3.905874e-18, 3.90766e-18, 
    3.906481e-18, 3.90843e-18, 3.9079e-18, 3.912278e-18, 3.913833e-18, 
    3.914574e-18, 3.915153e-18, 3.916635e-18, 3.915617e-18, 3.91602e-18, 
    3.915041e-18, 3.914432e-18, 3.914729e-18, 3.912865e-18, 3.913593e-18, 
    3.909809e-18, 3.911436e-18, 3.907147e-18, 3.908167e-18, 3.906899e-18, 
    3.907542e-18, 3.906449e-18, 3.907432e-18, 3.905714e-18, 3.905351e-18, 
    3.905601e-18, 3.90461e-18, 3.907489e-18, 3.906393e-18, 3.914742e-18, 
    3.914694e-18, 3.914461e-18, 3.915491e-18, 3.915549e-18, 3.916466e-18, 
    3.915641e-18, 3.915298e-18, 3.91439e-18, 3.913871e-18, 3.913371e-18, 
    3.912273e-18, 3.911063e-18, 3.909348e-18, 3.908102e-18, 3.907273e-18, 
    3.907775e-18, 3.907333e-18, 3.907831e-18, 3.908061e-18, 3.905493e-18, 
    3.906942e-18, 3.904753e-18, 3.90487e-18, 3.905868e-18, 3.904857e-18, 
    3.91466e-18, 3.914938e-18, 3.915935e-18, 3.915155e-18, 3.916565e-18, 
    3.915787e-18, 3.915346e-18, 3.913598e-18, 3.913192e-18, 3.912844e-18, 
    3.912137e-18, 3.911242e-18, 3.909679e-18, 3.908306e-18, 3.907042e-18, 
    3.907132e-18, 3.907101e-18, 3.906828e-18, 3.907517e-18, 3.906714e-18, 
    3.906589e-18, 3.906931e-18, 3.904887e-18, 3.905469e-18, 3.904873e-18, 
    3.90525e-18, 3.914845e-18, 3.914372e-18, 3.914629e-18, 3.914151e-18, 
    3.914495e-18, 3.912993e-18, 3.912543e-18, 3.910415e-18, 3.911264e-18, 
    3.909888e-18, 3.911118e-18, 3.910905e-18, 3.909881e-18, 3.911045e-18, 
    3.908399e-18, 3.910226e-18, 3.906818e-18, 3.908676e-18, 3.906703e-18, 
    3.907047e-18, 3.906469e-18, 3.905962e-18, 3.905307e-18, 3.904127e-18, 
    3.904396e-18, 3.903395e-18, 3.913659e-18, 3.913055e-18, 3.913091e-18, 
    3.912447e-18, 3.911975e-18, 3.910931e-18, 3.90928e-18, 3.909895e-18, 
    3.908747e-18, 3.908522e-18, 3.910256e-18, 3.909208e-18, 3.912638e-18, 
    3.912101e-18, 3.912408e-18, 3.913621e-18, 3.909777e-18, 3.911758e-18, 
    3.908085e-18, 3.909153e-18, 3.906037e-18, 3.907602e-18, 3.904548e-18, 
    3.90329e-18, 3.902028e-18, 3.900648e-18, 3.912707e-18, 3.913119e-18, 
    3.912365e-18, 3.911356e-18, 3.910371e-18, 3.909091e-18, 3.908951e-18, 
    3.908716e-18, 3.908087e-18, 3.907568e-18, 3.908659e-18, 3.907436e-18, 
    3.91201e-18, 3.909597e-18, 3.913291e-18, 3.9122e-18, 3.911408e-18, 
    3.911738e-18, 3.909961e-18, 3.909548e-18, 3.90788e-18, 3.908732e-18, 
    3.903616e-18, 3.905879e-18, 3.899542e-18, 3.90132e-18, 3.913267e-18, 
    3.9127e-18, 3.910754e-18, 3.911677e-18, 3.908997e-18, 3.908346e-18, 
    3.907801e-18, 3.907135e-18, 3.90705e-18, 3.906654e-18, 3.907306e-18, 
    3.906673e-18, 3.909088e-18, 3.908005e-18, 3.910955e-18, 3.910247e-18, 
    3.910567e-18, 3.910931e-18, 3.90981e-18, 3.908646e-18, 3.908593e-18, 
    3.908225e-18, 3.907237e-18, 3.908985e-18, 3.903375e-18, 3.906883e-18, 
    3.912084e-18, 3.911031e-18, 3.910847e-18, 3.911261e-18, 3.908412e-18, 
    3.909447e-18, 3.906659e-18, 3.907406e-18, 3.906176e-18, 3.906789e-18, 
    3.906881e-18, 3.907663e-18, 3.908158e-18, 3.909404e-18, 3.910412e-18, 
    3.911197e-18, 3.911012e-18, 3.910149e-18, 3.908568e-18, 3.907055e-18, 
    3.90739e-18, 3.906269e-18, 3.909191e-18, 3.907979e-18, 3.908457e-18, 
    3.907207e-18, 3.909917e-18, 3.907693e-18, 3.910496e-18, 3.910244e-18, 
    3.909467e-18, 3.907916e-18, 3.907531e-18, 3.907172e-18, 3.907388e-18, 
    3.908523e-18, 3.908697e-18, 3.909479e-18, 3.909709e-18, 3.910297e-18, 
    3.910797e-18, 3.910347e-18, 3.90988e-18, 3.908511e-18, 3.907294e-18, 
    3.905959e-18, 3.905621e-18, 3.904134e-18, 3.905382e-18, 3.903361e-18, 
    3.905136e-18, 3.902036e-18, 3.907523e-18, 3.905133e-18, 3.909422e-18, 
    3.908952e-18, 3.908133e-18, 3.906197e-18, 3.907212e-18, 3.906012e-18, 
    3.908701e-18, 3.910133e-18, 3.910469e-18, 3.911154e-18, 3.910454e-18, 
    3.91051e-18, 3.909842e-18, 3.910055e-18, 3.908465e-18, 3.909317e-18, 
    3.906891e-18, 3.906014e-18, 3.90351e-18, 3.901995e-18, 3.900411e-18, 
    3.899728e-18, 3.899517e-18, 3.899431e-18 ;

 MEG_formaldehyde =
  7.832728e-19, 7.82986e-19, 7.830404e-19, 7.828124e-19, 7.829367e-19, 
    7.82789e-19, 7.832122e-19, 7.829768e-19, 7.831256e-19, 7.832436e-19, 
    7.823775e-19, 7.828014e-19, 7.819153e-19, 7.821887e-19, 7.814957e-19, 
    7.819609e-19, 7.81401e-19, 7.815036e-19, 7.811818e-19, 7.812736e-19, 
    7.80874e-19, 7.811394e-19, 7.806584e-19, 7.809343e-19, 7.808932e-19, 
    7.81149e-19, 7.827109e-19, 7.824319e-19, 7.827287e-19, 7.826885e-19, 
    7.827054e-19, 7.829361e-19, 7.830561e-19, 7.83291e-19, 7.832473e-19, 
    7.830728e-19, 7.826704e-19, 7.828033e-19, 7.82458e-19, 7.824657e-19, 
    7.820857e-19, 7.82257e-19, 7.816155e-19, 7.817964e-19, 7.812697e-19, 
    7.814028e-19, 7.812768e-19, 7.813143e-19, 7.812764e-19, 7.814713e-19, 
    7.81388e-19, 7.815579e-19, 7.82226e-19, 7.820312e-19, 7.826157e-19, 
    7.829763e-19, 7.832029e-19, 7.833679e-19, 7.833445e-19, 7.833012e-19, 
    7.830718e-19, 7.828518e-19, 7.826859e-19, 7.82576e-19, 7.824668e-19, 
    7.821511e-19, 7.819723e-19, 7.815816e-19, 7.816474e-19, 7.815323e-19, 
    7.814158e-19, 7.812267e-19, 7.81257e-19, 7.811749e-19, 7.815319e-19, 
    7.812962e-19, 7.816861e-19, 7.815799e-19, 7.824556e-19, 7.827665e-19, 
    7.829148e-19, 7.830306e-19, 7.83327e-19, 7.831233e-19, 7.83204e-19, 
    7.830082e-19, 7.828865e-19, 7.829459e-19, 7.825729e-19, 7.827185e-19, 
    7.819618e-19, 7.822871e-19, 7.814294e-19, 7.816335e-19, 7.813798e-19, 
    7.815083e-19, 7.812897e-19, 7.814863e-19, 7.811428e-19, 7.810702e-19, 
    7.811202e-19, 7.80922e-19, 7.814978e-19, 7.812786e-19, 7.829484e-19, 
    7.829389e-19, 7.828922e-19, 7.830981e-19, 7.831097e-19, 7.832931e-19, 
    7.831282e-19, 7.830595e-19, 7.82878e-19, 7.827741e-19, 7.826742e-19, 
    7.824546e-19, 7.822126e-19, 7.818696e-19, 7.816204e-19, 7.814546e-19, 
    7.81555e-19, 7.814665e-19, 7.815662e-19, 7.816122e-19, 7.810986e-19, 
    7.813883e-19, 7.809505e-19, 7.80974e-19, 7.811736e-19, 7.809714e-19, 
    7.829318e-19, 7.829875e-19, 7.83187e-19, 7.830309e-19, 7.833128e-19, 
    7.831573e-19, 7.830692e-19, 7.827196e-19, 7.826383e-19, 7.825688e-19, 
    7.824274e-19, 7.822484e-19, 7.819357e-19, 7.816612e-19, 7.814083e-19, 
    7.814265e-19, 7.814202e-19, 7.813657e-19, 7.815033e-19, 7.813429e-19, 
    7.813177e-19, 7.813862e-19, 7.809774e-19, 7.810938e-19, 7.809746e-19, 
    7.810499e-19, 7.829689e-19, 7.828744e-19, 7.829258e-19, 7.828302e-19, 
    7.828989e-19, 7.825985e-19, 7.825085e-19, 7.82083e-19, 7.822529e-19, 
    7.819775e-19, 7.822234e-19, 7.821809e-19, 7.819762e-19, 7.822089e-19, 
    7.816799e-19, 7.820452e-19, 7.813635e-19, 7.817352e-19, 7.813406e-19, 
    7.814093e-19, 7.812938e-19, 7.811923e-19, 7.810614e-19, 7.808253e-19, 
    7.808792e-19, 7.80679e-19, 7.827318e-19, 7.82611e-19, 7.826182e-19, 
    7.824894e-19, 7.82395e-19, 7.821862e-19, 7.818559e-19, 7.819789e-19, 
    7.817493e-19, 7.817044e-19, 7.820512e-19, 7.818416e-19, 7.825275e-19, 
    7.824202e-19, 7.824815e-19, 7.827242e-19, 7.819553e-19, 7.823516e-19, 
    7.81617e-19, 7.818305e-19, 7.812073e-19, 7.815204e-19, 7.809096e-19, 
    7.80658e-19, 7.804056e-19, 7.801296e-19, 7.825413e-19, 7.826237e-19, 
    7.824731e-19, 7.822712e-19, 7.820742e-19, 7.818182e-19, 7.817901e-19, 
    7.817432e-19, 7.816174e-19, 7.815135e-19, 7.817317e-19, 7.814872e-19, 
    7.824021e-19, 7.819194e-19, 7.826581e-19, 7.8244e-19, 7.822816e-19, 
    7.823476e-19, 7.819921e-19, 7.819096e-19, 7.815761e-19, 7.817465e-19, 
    7.807231e-19, 7.811757e-19, 7.799084e-19, 7.802639e-19, 7.826534e-19, 
    7.825399e-19, 7.821508e-19, 7.823353e-19, 7.817993e-19, 7.816691e-19, 
    7.815603e-19, 7.81427e-19, 7.814101e-19, 7.813307e-19, 7.814612e-19, 
    7.813345e-19, 7.818177e-19, 7.81601e-19, 7.821911e-19, 7.820494e-19, 
    7.821134e-19, 7.821862e-19, 7.81962e-19, 7.817292e-19, 7.817186e-19, 
    7.816449e-19, 7.814473e-19, 7.817969e-19, 7.806749e-19, 7.813766e-19, 
    7.824167e-19, 7.822062e-19, 7.821694e-19, 7.822521e-19, 7.816824e-19, 
    7.818893e-19, 7.813319e-19, 7.814812e-19, 7.812352e-19, 7.813578e-19, 
    7.813762e-19, 7.815325e-19, 7.816316e-19, 7.818808e-19, 7.820823e-19, 
    7.822394e-19, 7.822024e-19, 7.820298e-19, 7.817136e-19, 7.814111e-19, 
    7.81478e-19, 7.812538e-19, 7.818382e-19, 7.815958e-19, 7.816913e-19, 
    7.814414e-19, 7.819834e-19, 7.815385e-19, 7.820992e-19, 7.820489e-19, 
    7.818933e-19, 7.815831e-19, 7.815063e-19, 7.814343e-19, 7.814776e-19, 
    7.817045e-19, 7.817393e-19, 7.818958e-19, 7.819418e-19, 7.820594e-19, 
    7.821595e-19, 7.820694e-19, 7.81976e-19, 7.817022e-19, 7.814587e-19, 
    7.811917e-19, 7.811242e-19, 7.808267e-19, 7.810764e-19, 7.806721e-19, 
    7.810271e-19, 7.804071e-19, 7.815045e-19, 7.810267e-19, 7.818844e-19, 
    7.817905e-19, 7.816265e-19, 7.812395e-19, 7.814425e-19, 7.812023e-19, 
    7.817402e-19, 7.820266e-19, 7.820939e-19, 7.822308e-19, 7.820907e-19, 
    7.821019e-19, 7.819683e-19, 7.820109e-19, 7.81693e-19, 7.818635e-19, 
    7.813781e-19, 7.812028e-19, 7.807019e-19, 7.803989e-19, 7.800823e-19, 
    7.799455e-19, 7.799034e-19, 7.798861e-19 ;

 MEG_isoprene =
  6.252753e-19, 6.250062e-19, 6.250573e-19, 6.248433e-19, 6.2496e-19, 
    6.248214e-19, 6.252184e-19, 6.249976e-19, 6.251373e-19, 6.252479e-19, 
    6.244353e-19, 6.248331e-19, 6.240017e-19, 6.242582e-19, 6.23608e-19, 
    6.240445e-19, 6.235191e-19, 6.236154e-19, 6.233134e-19, 6.233996e-19, 
    6.230245e-19, 6.232736e-19, 6.228221e-19, 6.230811e-19, 6.230426e-19, 
    6.232826e-19, 6.247481e-19, 6.244864e-19, 6.247648e-19, 6.247272e-19, 
    6.247429e-19, 6.249594e-19, 6.25072e-19, 6.252923e-19, 6.252514e-19, 
    6.250876e-19, 6.247102e-19, 6.248348e-19, 6.245109e-19, 6.245181e-19, 
    6.241615e-19, 6.243223e-19, 6.237203e-19, 6.238901e-19, 6.233959e-19, 
    6.235208e-19, 6.234026e-19, 6.234378e-19, 6.234021e-19, 6.23585e-19, 
    6.23507e-19, 6.236664e-19, 6.242932e-19, 6.241104e-19, 6.246589e-19, 
    6.249972e-19, 6.252097e-19, 6.253644e-19, 6.253426e-19, 6.253019e-19, 
    6.250867e-19, 6.248804e-19, 6.247247e-19, 6.246216e-19, 6.245191e-19, 
    6.24223e-19, 6.240551e-19, 6.236885e-19, 6.237503e-19, 6.236423e-19, 
    6.23533e-19, 6.233555e-19, 6.23384e-19, 6.233069e-19, 6.23642e-19, 
    6.234208e-19, 6.237866e-19, 6.23687e-19, 6.245086e-19, 6.248003e-19, 
    6.249395e-19, 6.250481e-19, 6.253261e-19, 6.251351e-19, 6.252108e-19, 
    6.250271e-19, 6.249129e-19, 6.249686e-19, 6.246187e-19, 6.247553e-19, 
    6.240453e-19, 6.243505e-19, 6.235458e-19, 6.237372e-19, 6.234992e-19, 
    6.236198e-19, 6.234146e-19, 6.235992e-19, 6.232768e-19, 6.232086e-19, 
    6.232556e-19, 6.230696e-19, 6.236099e-19, 6.234043e-19, 6.24971e-19, 
    6.24962e-19, 6.249182e-19, 6.251114e-19, 6.251223e-19, 6.252944e-19, 
    6.251396e-19, 6.250752e-19, 6.249049e-19, 6.248075e-19, 6.247137e-19, 
    6.245077e-19, 6.242807e-19, 6.239588e-19, 6.23725e-19, 6.235694e-19, 
    6.236637e-19, 6.235806e-19, 6.236741e-19, 6.237172e-19, 6.232354e-19, 
    6.235072e-19, 6.230963e-19, 6.231184e-19, 6.233057e-19, 6.231159e-19, 
    6.249554e-19, 6.250077e-19, 6.251948e-19, 6.250483e-19, 6.253129e-19, 
    6.25167e-19, 6.250843e-19, 6.247562e-19, 6.2468e-19, 6.246149e-19, 
    6.244822e-19, 6.243142e-19, 6.240208e-19, 6.237633e-19, 6.235259e-19, 
    6.23543e-19, 6.235371e-19, 6.234859e-19, 6.236151e-19, 6.234646e-19, 
    6.23441e-19, 6.235053e-19, 6.231215e-19, 6.232309e-19, 6.231189e-19, 
    6.231897e-19, 6.249902e-19, 6.249016e-19, 6.249497e-19, 6.2486e-19, 
    6.249246e-19, 6.246427e-19, 6.245582e-19, 6.24159e-19, 6.243184e-19, 
    6.2406e-19, 6.242908e-19, 6.242509e-19, 6.240588e-19, 6.242772e-19, 
    6.237808e-19, 6.241236e-19, 6.23484e-19, 6.238327e-19, 6.234625e-19, 
    6.23527e-19, 6.234185e-19, 6.233233e-19, 6.232004e-19, 6.229788e-19, 
    6.230293e-19, 6.228415e-19, 6.247677e-19, 6.246544e-19, 6.246612e-19, 
    6.245403e-19, 6.244517e-19, 6.242559e-19, 6.23946e-19, 6.240613e-19, 
    6.238459e-19, 6.238038e-19, 6.241292e-19, 6.239325e-19, 6.245761e-19, 
    6.244754e-19, 6.245329e-19, 6.247606e-19, 6.240393e-19, 6.24411e-19, 
    6.237218e-19, 6.239222e-19, 6.233373e-19, 6.236312e-19, 6.23058e-19, 
    6.228218e-19, 6.225849e-19, 6.223257e-19, 6.24589e-19, 6.246664e-19, 
    6.24525e-19, 6.243356e-19, 6.241508e-19, 6.239106e-19, 6.238842e-19, 
    6.238402e-19, 6.237222e-19, 6.236247e-19, 6.238294e-19, 6.235999e-19, 
    6.244584e-19, 6.240055e-19, 6.246986e-19, 6.24494e-19, 6.243453e-19, 
    6.244073e-19, 6.240738e-19, 6.239964e-19, 6.236834e-19, 6.238433e-19, 
    6.228829e-19, 6.233076e-19, 6.22118e-19, 6.224518e-19, 6.246942e-19, 
    6.245877e-19, 6.242226e-19, 6.243957e-19, 6.238928e-19, 6.237707e-19, 
    6.236686e-19, 6.235435e-19, 6.235276e-19, 6.234531e-19, 6.235756e-19, 
    6.234567e-19, 6.239101e-19, 6.237068e-19, 6.242604e-19, 6.241275e-19, 
    6.241875e-19, 6.242558e-19, 6.240455e-19, 6.23827e-19, 6.238171e-19, 
    6.23748e-19, 6.235627e-19, 6.238906e-19, 6.228377e-19, 6.234962e-19, 
    6.244721e-19, 6.242747e-19, 6.242401e-19, 6.243177e-19, 6.237831e-19, 
    6.239773e-19, 6.234542e-19, 6.235943e-19, 6.233635e-19, 6.234786e-19, 
    6.234958e-19, 6.236425e-19, 6.237354e-19, 6.239694e-19, 6.241584e-19, 
    6.243057e-19, 6.24271e-19, 6.241091e-19, 6.238124e-19, 6.235285e-19, 
    6.235914e-19, 6.233809e-19, 6.239294e-19, 6.237019e-19, 6.237915e-19, 
    6.23557e-19, 6.240655e-19, 6.236482e-19, 6.241743e-19, 6.24127e-19, 
    6.239811e-19, 6.2369e-19, 6.236179e-19, 6.235504e-19, 6.23591e-19, 
    6.238039e-19, 6.238366e-19, 6.239834e-19, 6.240265e-19, 6.241369e-19, 
    6.242308e-19, 6.241463e-19, 6.240587e-19, 6.238018e-19, 6.235732e-19, 
    6.233227e-19, 6.232594e-19, 6.229801e-19, 6.232145e-19, 6.228351e-19, 
    6.231683e-19, 6.225863e-19, 6.236163e-19, 6.231678e-19, 6.239727e-19, 
    6.238845e-19, 6.237307e-19, 6.233675e-19, 6.235581e-19, 6.233327e-19, 
    6.238374e-19, 6.241061e-19, 6.241692e-19, 6.242977e-19, 6.241663e-19, 
    6.241767e-19, 6.240514e-19, 6.240913e-19, 6.237931e-19, 6.23953e-19, 
    6.234976e-19, 6.233331e-19, 6.22863e-19, 6.225786e-19, 6.222813e-19, 
    6.221529e-19, 6.221134e-19, 6.220972e-19 ;

 MEG_methanol =
  8.573298e-17, 8.571827e-17, 8.572106e-17, 8.570935e-17, 8.571574e-17, 
    8.570815e-17, 8.572988e-17, 8.571779e-17, 8.572543e-17, 8.573149e-17, 
    8.568704e-17, 8.57088e-17, 8.566333e-17, 8.567736e-17, 8.56418e-17, 
    8.566566e-17, 8.563694e-17, 8.56422e-17, 8.562571e-17, 8.563042e-17, 
    8.560994e-17, 8.562354e-17, 8.559891e-17, 8.561303e-17, 8.561093e-17, 
    8.562403e-17, 8.570414e-17, 8.568983e-17, 8.570506e-17, 8.5703e-17, 
    8.570387e-17, 8.57157e-17, 8.572186e-17, 8.573392e-17, 8.573168e-17, 
    8.572272e-17, 8.570207e-17, 8.570889e-17, 8.569117e-17, 8.569156e-17, 
    8.567208e-17, 8.568086e-17, 8.564794e-17, 8.565723e-17, 8.563022e-17, 
    8.563704e-17, 8.563058e-17, 8.56325e-17, 8.563056e-17, 8.564055e-17, 
    8.563628e-17, 8.564499e-17, 8.567928e-17, 8.566928e-17, 8.569927e-17, 
    8.571776e-17, 8.57294e-17, 8.573787e-17, 8.573667e-17, 8.573444e-17, 
    8.572267e-17, 8.571138e-17, 8.570287e-17, 8.569723e-17, 8.569162e-17, 
    8.567542e-17, 8.566625e-17, 8.56462e-17, 8.564958e-17, 8.564367e-17, 
    8.56377e-17, 8.562801e-17, 8.562957e-17, 8.562536e-17, 8.564366e-17, 
    8.563158e-17, 8.565157e-17, 8.564612e-17, 8.569104e-17, 8.5707e-17, 
    8.571461e-17, 8.572055e-17, 8.573577e-17, 8.572531e-17, 8.572946e-17, 
    8.57194e-17, 8.571316e-17, 8.571621e-17, 8.569707e-17, 8.570454e-17, 
    8.566572e-17, 8.568241e-17, 8.56384e-17, 8.564886e-17, 8.563586e-17, 
    8.564245e-17, 8.563124e-17, 8.564132e-17, 8.562372e-17, 8.562e-17, 
    8.562256e-17, 8.561241e-17, 8.564191e-17, 8.563067e-17, 8.571634e-17, 
    8.571585e-17, 8.571345e-17, 8.572402e-17, 8.572462e-17, 8.573403e-17, 
    8.572556e-17, 8.572204e-17, 8.571272e-17, 8.570739e-17, 8.570226e-17, 
    8.5691e-17, 8.567859e-17, 8.566098e-17, 8.564819e-17, 8.56397e-17, 
    8.564484e-17, 8.564031e-17, 8.564541e-17, 8.564777e-17, 8.562145e-17, 
    8.563629e-17, 8.561387e-17, 8.561507e-17, 8.562529e-17, 8.561494e-17, 
    8.571549e-17, 8.571834e-17, 8.572858e-17, 8.572057e-17, 8.573505e-17, 
    8.572706e-17, 8.572253e-17, 8.570459e-17, 8.570042e-17, 8.569686e-17, 
    8.568961e-17, 8.568042e-17, 8.566437e-17, 8.565028e-17, 8.563732e-17, 
    8.563825e-17, 8.563793e-17, 8.563514e-17, 8.564219e-17, 8.563397e-17, 
    8.563268e-17, 8.563619e-17, 8.561524e-17, 8.562121e-17, 8.56151e-17, 
    8.561896e-17, 8.571739e-17, 8.571254e-17, 8.571517e-17, 8.571027e-17, 
    8.57138e-17, 8.569838e-17, 8.569376e-17, 8.567193e-17, 8.568065e-17, 
    8.566652e-17, 8.567914e-17, 8.567696e-17, 8.566645e-17, 8.56784e-17, 
    8.565125e-17, 8.566999e-17, 8.563502e-17, 8.565408e-17, 8.563385e-17, 
    8.563737e-17, 8.563145e-17, 8.562625e-17, 8.561955e-17, 8.560746e-17, 
    8.561021e-17, 8.559997e-17, 8.570522e-17, 8.569902e-17, 8.569939e-17, 
    8.569279e-17, 8.568794e-17, 8.567723e-17, 8.566028e-17, 8.56666e-17, 
    8.565482e-17, 8.565251e-17, 8.567031e-17, 8.565954e-17, 8.569474e-17, 
    8.568923e-17, 8.569238e-17, 8.570483e-17, 8.566539e-17, 8.568571e-17, 
    8.564802e-17, 8.565899e-17, 8.562702e-17, 8.564306e-17, 8.561177e-17, 
    8.559889e-17, 8.558598e-17, 8.557186e-17, 8.569545e-17, 8.569968e-17, 
    8.569195e-17, 8.568159e-17, 8.567149e-17, 8.565835e-17, 8.565691e-17, 
    8.565451e-17, 8.564804e-17, 8.564271e-17, 8.565391e-17, 8.564136e-17, 
    8.56883e-17, 8.566354e-17, 8.570144e-17, 8.569025e-17, 8.568212e-17, 
    8.568551e-17, 8.566727e-17, 8.566304e-17, 8.564592e-17, 8.565467e-17, 
    8.560222e-17, 8.56254e-17, 8.556056e-17, 8.557873e-17, 8.57012e-17, 
    8.569538e-17, 8.567541e-17, 8.568488e-17, 8.565738e-17, 8.56507e-17, 
    8.564511e-17, 8.563828e-17, 8.563741e-17, 8.563334e-17, 8.564003e-17, 
    8.563354e-17, 8.565832e-17, 8.56472e-17, 8.567748e-17, 8.567021e-17, 
    8.56735e-17, 8.567723e-17, 8.566573e-17, 8.565378e-17, 8.565324e-17, 
    8.564945e-17, 8.563931e-17, 8.565726e-17, 8.559975e-17, 8.563569e-17, 
    8.568906e-17, 8.567826e-17, 8.567637e-17, 8.568061e-17, 8.565138e-17, 
    8.5662e-17, 8.56334e-17, 8.564105e-17, 8.562845e-17, 8.563473e-17, 
    8.563567e-17, 8.564369e-17, 8.564877e-17, 8.566156e-17, 8.56719e-17, 
    8.567996e-17, 8.567806e-17, 8.56692e-17, 8.565298e-17, 8.563746e-17, 
    8.564089e-17, 8.56294e-17, 8.565938e-17, 8.564693e-17, 8.565184e-17, 
    8.563901e-17, 8.566682e-17, 8.564399e-17, 8.567277e-17, 8.567018e-17, 
    8.56622e-17, 8.564628e-17, 8.564234e-17, 8.563865e-17, 8.564087e-17, 
    8.565252e-17, 8.56543e-17, 8.566233e-17, 8.566469e-17, 8.567073e-17, 
    8.567586e-17, 8.567124e-17, 8.566644e-17, 8.56524e-17, 8.56399e-17, 
    8.562622e-17, 8.562276e-17, 8.560752e-17, 8.562031e-17, 8.55996e-17, 
    8.561778e-17, 8.558605e-17, 8.564224e-17, 8.561776e-17, 8.566175e-17, 
    8.565693e-17, 8.56485e-17, 8.562866e-17, 8.563907e-17, 8.562677e-17, 
    8.565435e-17, 8.566904e-17, 8.567249e-17, 8.567952e-17, 8.567233e-17, 
    8.56729e-17, 8.566605e-17, 8.566824e-17, 8.565193e-17, 8.566067e-17, 
    8.563577e-17, 8.562679e-17, 8.560114e-17, 8.558564e-17, 8.556945e-17, 
    8.556246e-17, 8.556031e-17, 8.555943e-17 ;

 MEG_pinene_a =
  7.460954e-17, 7.459339e-17, 7.459646e-17, 7.458361e-17, 7.459062e-17, 
    7.45823e-17, 7.460613e-17, 7.459287e-17, 7.460126e-17, 7.46079e-17, 
    7.455914e-17, 7.4583e-17, 7.453313e-17, 7.454851e-17, 7.450951e-17, 
    7.453569e-17, 7.450419e-17, 7.450995e-17, 7.449186e-17, 7.449702e-17, 
    7.447456e-17, 7.448948e-17, 7.446245e-17, 7.447795e-17, 7.447564e-17, 
    7.449002e-17, 7.45779e-17, 7.45622e-17, 7.457891e-17, 7.457665e-17, 
    7.45776e-17, 7.459058e-17, 7.459734e-17, 7.461057e-17, 7.460811e-17, 
    7.459828e-17, 7.457563e-17, 7.45831e-17, 7.456368e-17, 7.456411e-17, 
    7.454272e-17, 7.455236e-17, 7.451625e-17, 7.452643e-17, 7.449681e-17, 
    7.450429e-17, 7.449721e-17, 7.449931e-17, 7.449718e-17, 7.450814e-17, 
    7.450346e-17, 7.451301e-17, 7.455061e-17, 7.453965e-17, 7.457255e-17, 
    7.459284e-17, 7.46056e-17, 7.461489e-17, 7.461358e-17, 7.461114e-17, 
    7.459822e-17, 7.458584e-17, 7.457651e-17, 7.457031e-17, 7.456416e-17, 
    7.45464e-17, 7.453633e-17, 7.451434e-17, 7.451805e-17, 7.451157e-17, 
    7.450502e-17, 7.449438e-17, 7.44961e-17, 7.449147e-17, 7.451155e-17, 
    7.449829e-17, 7.452023e-17, 7.451425e-17, 7.456353e-17, 7.458104e-17, 
    7.458938e-17, 7.459591e-17, 7.461259e-17, 7.460112e-17, 7.460567e-17, 
    7.459464e-17, 7.458779e-17, 7.459114e-17, 7.457014e-17, 7.457833e-17, 
    7.453574e-17, 7.455405e-17, 7.450579e-17, 7.451727e-17, 7.4503e-17, 
    7.451022e-17, 7.449793e-17, 7.450899e-17, 7.448967e-17, 7.448559e-17, 
    7.44884e-17, 7.447726e-17, 7.450963e-17, 7.449731e-17, 7.459128e-17, 
    7.459074e-17, 7.458811e-17, 7.459971e-17, 7.460036e-17, 7.461069e-17, 
    7.46014e-17, 7.459754e-17, 7.458731e-17, 7.458147e-17, 7.457584e-17, 
    7.456348e-17, 7.454986e-17, 7.453055e-17, 7.451653e-17, 7.45072e-17, 
    7.451285e-17, 7.450787e-17, 7.451348e-17, 7.451606e-17, 7.448718e-17, 
    7.450348e-17, 7.447887e-17, 7.448019e-17, 7.44914e-17, 7.448004e-17, 
    7.459034e-17, 7.459348e-17, 7.460472e-17, 7.459592e-17, 7.46118e-17, 
    7.460304e-17, 7.459808e-17, 7.457839e-17, 7.457382e-17, 7.456991e-17, 
    7.456195e-17, 7.455188e-17, 7.453427e-17, 7.451882e-17, 7.450459e-17, 
    7.450562e-17, 7.450527e-17, 7.45022e-17, 7.450994e-17, 7.450092e-17, 
    7.449951e-17, 7.450336e-17, 7.448037e-17, 7.448692e-17, 7.448022e-17, 
    7.448445e-17, 7.459243e-17, 7.458711e-17, 7.459001e-17, 7.458462e-17, 
    7.458849e-17, 7.457158e-17, 7.456651e-17, 7.454257e-17, 7.455213e-17, 
    7.453662e-17, 7.455047e-17, 7.454808e-17, 7.453655e-17, 7.454966e-17, 
    7.451988e-17, 7.454044e-17, 7.450208e-17, 7.452299e-17, 7.45008e-17, 
    7.450466e-17, 7.449816e-17, 7.449245e-17, 7.448509e-17, 7.447182e-17, 
    7.447485e-17, 7.446361e-17, 7.457908e-17, 7.457228e-17, 7.457269e-17, 
    7.456544e-17, 7.456013e-17, 7.454838e-17, 7.452979e-17, 7.453671e-17, 
    7.452379e-17, 7.452126e-17, 7.454078e-17, 7.452898e-17, 7.456759e-17, 
    7.456154e-17, 7.4565e-17, 7.457866e-17, 7.453538e-17, 7.455768e-17, 
    7.451634e-17, 7.452836e-17, 7.449329e-17, 7.45109e-17, 7.447656e-17, 
    7.446243e-17, 7.444825e-17, 7.443276e-17, 7.456836e-17, 7.4573e-17, 
    7.456452e-17, 7.455316e-17, 7.454208e-17, 7.452767e-17, 7.452608e-17, 
    7.452345e-17, 7.451636e-17, 7.451052e-17, 7.45228e-17, 7.450903e-17, 
    7.456052e-17, 7.453336e-17, 7.457493e-17, 7.456266e-17, 7.455374e-17, 
    7.455745e-17, 7.453745e-17, 7.453281e-17, 7.451403e-17, 7.452363e-17, 
    7.446608e-17, 7.449152e-17, 7.442034e-17, 7.444029e-17, 7.457467e-17, 
    7.456829e-17, 7.454638e-17, 7.455677e-17, 7.45266e-17, 7.451928e-17, 
    7.451314e-17, 7.450565e-17, 7.45047e-17, 7.450023e-17, 7.450757e-17, 
    7.450045e-17, 7.452764e-17, 7.451544e-17, 7.454865e-17, 7.454067e-17, 
    7.454428e-17, 7.454838e-17, 7.453576e-17, 7.452265e-17, 7.452206e-17, 
    7.451791e-17, 7.450679e-17, 7.452647e-17, 7.446337e-17, 7.450281e-17, 
    7.456135e-17, 7.45495e-17, 7.454743e-17, 7.455209e-17, 7.452002e-17, 
    7.453167e-17, 7.45003e-17, 7.45087e-17, 7.449487e-17, 7.450176e-17, 
    7.450279e-17, 7.451159e-17, 7.451715e-17, 7.453119e-17, 7.454253e-17, 
    7.455137e-17, 7.454929e-17, 7.453957e-17, 7.452178e-17, 7.450475e-17, 
    7.450852e-17, 7.449591e-17, 7.452879e-17, 7.451514e-17, 7.452052e-17, 
    7.450646e-17, 7.453696e-17, 7.451192e-17, 7.454348e-17, 7.454065e-17, 
    7.453189e-17, 7.451443e-17, 7.451011e-17, 7.450606e-17, 7.45085e-17, 
    7.452127e-17, 7.452323e-17, 7.453203e-17, 7.453462e-17, 7.454124e-17, 
    7.454687e-17, 7.45418e-17, 7.453654e-17, 7.452114e-17, 7.450743e-17, 
    7.449243e-17, 7.448863e-17, 7.44719e-17, 7.448593e-17, 7.446321e-17, 
    7.448316e-17, 7.444833e-17, 7.451001e-17, 7.448314e-17, 7.453139e-17, 
    7.452611e-17, 7.451687e-17, 7.449511e-17, 7.450652e-17, 7.449302e-17, 
    7.452328e-17, 7.453939e-17, 7.454318e-17, 7.455089e-17, 7.4543e-17, 
    7.454363e-17, 7.453611e-17, 7.453851e-17, 7.452062e-17, 7.453021e-17, 
    7.45029e-17, 7.449304e-17, 7.446489e-17, 7.444788e-17, 7.44301e-17, 
    7.442243e-17, 7.442006e-17, 7.44191e-17 ;

 MEG_thujene_a =
  1.797641e-18, 1.797282e-18, 1.79735e-18, 1.797064e-18, 1.79722e-18, 
    1.797035e-18, 1.797565e-18, 1.79727e-18, 1.797456e-18, 1.797604e-18, 
    1.79652e-18, 1.797051e-18, 1.795941e-18, 1.796283e-18, 1.795416e-18, 
    1.795998e-18, 1.795298e-18, 1.795426e-18, 1.795024e-18, 1.795138e-18, 
    1.794639e-18, 1.794971e-18, 1.79437e-18, 1.794714e-18, 1.794663e-18, 
    1.794983e-18, 1.796937e-18, 1.796588e-18, 1.796959e-18, 1.796909e-18, 
    1.79693e-18, 1.797219e-18, 1.797369e-18, 1.797664e-18, 1.797609e-18, 
    1.79739e-18, 1.796886e-18, 1.797053e-18, 1.796621e-18, 1.79663e-18, 
    1.796154e-18, 1.796369e-18, 1.795566e-18, 1.795792e-18, 1.795134e-18, 
    1.7953e-18, 1.795142e-18, 1.795189e-18, 1.795142e-18, 1.795386e-18, 
    1.795282e-18, 1.795494e-18, 1.79633e-18, 1.796086e-18, 1.796818e-18, 
    1.797269e-18, 1.797553e-18, 1.79776e-18, 1.797731e-18, 1.797676e-18, 
    1.797389e-18, 1.797114e-18, 1.796906e-18, 1.796768e-18, 1.796632e-18, 
    1.796236e-18, 1.796013e-18, 1.795524e-18, 1.795606e-18, 1.795462e-18, 
    1.795316e-18, 1.79508e-18, 1.795118e-18, 1.795015e-18, 1.795461e-18, 
    1.795167e-18, 1.795654e-18, 1.795521e-18, 1.796617e-18, 1.797007e-18, 
    1.797192e-18, 1.797338e-18, 1.797709e-18, 1.797454e-18, 1.797555e-18, 
    1.797309e-18, 1.797157e-18, 1.797231e-18, 1.796765e-18, 1.796947e-18, 
    1.795999e-18, 1.796407e-18, 1.795333e-18, 1.795588e-18, 1.795271e-18, 
    1.795432e-18, 1.795159e-18, 1.795404e-18, 1.794975e-18, 1.794884e-18, 
    1.794947e-18, 1.794699e-18, 1.795419e-18, 1.795145e-18, 1.797235e-18, 
    1.797223e-18, 1.797164e-18, 1.797422e-18, 1.797437e-18, 1.797666e-18, 
    1.79746e-18, 1.797374e-18, 1.797146e-18, 1.797016e-18, 1.796891e-18, 
    1.796616e-18, 1.796313e-18, 1.795884e-18, 1.795572e-18, 1.795365e-18, 
    1.79549e-18, 1.79538e-18, 1.795504e-18, 1.795562e-18, 1.79492e-18, 
    1.795282e-18, 1.794735e-18, 1.794764e-18, 1.795013e-18, 1.794761e-18, 
    1.797214e-18, 1.797284e-18, 1.797533e-18, 1.797338e-18, 1.797691e-18, 
    1.797496e-18, 1.797386e-18, 1.796948e-18, 1.796846e-18, 1.796759e-18, 
    1.796582e-18, 1.796358e-18, 1.795967e-18, 1.795623e-18, 1.795307e-18, 
    1.79533e-18, 1.795322e-18, 1.795253e-18, 1.795426e-18, 1.795225e-18, 
    1.795193e-18, 1.795279e-18, 1.794768e-18, 1.794914e-18, 1.794765e-18, 
    1.794859e-18, 1.79726e-18, 1.797142e-18, 1.797206e-18, 1.797086e-18, 
    1.797173e-18, 1.796796e-18, 1.796684e-18, 1.796151e-18, 1.796364e-18, 
    1.796019e-18, 1.796327e-18, 1.796274e-18, 1.796017e-18, 1.796309e-18, 
    1.795647e-18, 1.796104e-18, 1.795251e-18, 1.795716e-18, 1.795222e-18, 
    1.795308e-18, 1.795164e-18, 1.795037e-18, 1.794873e-18, 1.794578e-18, 
    1.794645e-18, 1.794395e-18, 1.796963e-18, 1.796812e-18, 1.796821e-18, 
    1.79666e-18, 1.796542e-18, 1.79628e-18, 1.795867e-18, 1.796021e-18, 
    1.795734e-18, 1.795678e-18, 1.796111e-18, 1.795849e-18, 1.796708e-18, 
    1.796573e-18, 1.79665e-18, 1.796954e-18, 1.795991e-18, 1.796487e-18, 
    1.795568e-18, 1.795835e-18, 1.795056e-18, 1.795447e-18, 1.794684e-18, 
    1.794369e-18, 1.794054e-18, 1.79371e-18, 1.796725e-18, 1.796828e-18, 
    1.796639e-18, 1.796387e-18, 1.79614e-18, 1.79582e-18, 1.795785e-18, 
    1.795726e-18, 1.795568e-18, 1.795438e-18, 1.795712e-18, 1.795405e-18, 
    1.79655e-18, 1.795946e-18, 1.796871e-18, 1.796598e-18, 1.7964e-18, 
    1.796482e-18, 1.796037e-18, 1.795934e-18, 1.795517e-18, 1.79573e-18, 
    1.79445e-18, 1.795016e-18, 1.793434e-18, 1.793877e-18, 1.796865e-18, 
    1.796723e-18, 1.796236e-18, 1.796467e-18, 1.795796e-18, 1.795633e-18, 
    1.795497e-18, 1.79533e-18, 1.795309e-18, 1.79521e-18, 1.795373e-18, 
    1.795215e-18, 1.795819e-18, 1.795548e-18, 1.796287e-18, 1.796109e-18, 
    1.796189e-18, 1.79628e-18, 1.796e-18, 1.795708e-18, 1.795695e-18, 
    1.795603e-18, 1.795355e-18, 1.795793e-18, 1.79439e-18, 1.795267e-18, 
    1.796569e-18, 1.796305e-18, 1.796259e-18, 1.796363e-18, 1.79565e-18, 
    1.795909e-18, 1.795211e-18, 1.795398e-18, 1.79509e-18, 1.795244e-18, 
    1.795267e-18, 1.795462e-18, 1.795586e-18, 1.795898e-18, 1.79615e-18, 
    1.796347e-18, 1.796301e-18, 1.796085e-18, 1.795689e-18, 1.79531e-18, 
    1.795394e-18, 1.795114e-18, 1.795845e-18, 1.795541e-18, 1.795661e-18, 
    1.795348e-18, 1.796026e-18, 1.79547e-18, 1.796172e-18, 1.796109e-18, 
    1.795914e-18, 1.795525e-18, 1.795429e-18, 1.795339e-18, 1.795393e-18, 
    1.795678e-18, 1.795721e-18, 1.795917e-18, 1.795974e-18, 1.796122e-18, 
    1.796247e-18, 1.796134e-18, 1.796017e-18, 1.795675e-18, 1.79537e-18, 
    1.795036e-18, 1.794952e-18, 1.79458e-18, 1.794892e-18, 1.794387e-18, 
    1.79483e-18, 1.794056e-18, 1.795427e-18, 1.79483e-18, 1.795903e-18, 
    1.795785e-18, 1.79558e-18, 1.795096e-18, 1.79535e-18, 1.795049e-18, 
    1.795722e-18, 1.796081e-18, 1.796165e-18, 1.796336e-18, 1.796161e-18, 
    1.796175e-18, 1.796008e-18, 1.796061e-18, 1.795663e-18, 1.795877e-18, 
    1.795269e-18, 1.79505e-18, 1.794424e-18, 1.794046e-18, 1.793651e-18, 
    1.79348e-18, 1.793428e-18, 1.793406e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -4.312828e-25, 1.730626e-25, -2.472314e-26, 1.648223e-26, 8.515785e-26, 
    -1.263631e-25, 2.884377e-25, -1.263631e-25, -1.126279e-25, 1.785567e-25, 
    2.472323e-25, -1.098809e-25, -2.499792e-25, -1.758095e-25, 2.197628e-26, 
    -4.010655e-25, -3.571131e-25, -3.021719e-26, -6.867554e-26, 
    -8.790471e-26, 3.57114e-26, 4.3403e-25, -7.966364e-26, 2.719555e-25, 
    -2.884375e-25, 1.813037e-25, 2.582204e-25, -8.790471e-26, 8.257562e-32, 
    -5.164406e-25, -1.593274e-25, 2.225091e-25, 4.120545e-26, -2.33497e-25, 
    1.620745e-25, -5.466578e-25, 1.785567e-25, -1.483393e-25, -5.768744e-26, 
    3.735955e-25, 1.098818e-26, -5.686341e-25, 2.032799e-25, -1.538333e-25, 
    -3.543661e-25, 2.911847e-25, 1.922926e-26, -2.911845e-25, -2.747016e-26, 
    4.395248e-26, -4.395231e-26, 1.098811e-25, 3.653544e-25, 5.603931e-25, 
    1.153751e-25, -4.56006e-25, 8.790487e-26, 4.120545e-26, 3.159079e-25, 
    8.257626e-32, 3.021735e-26, -2.692083e-25, -1.126279e-25, 3.296438e-26, 
    5.76876e-26, -4.257888e-25, -2.856905e-25, 1.813037e-25, 6.867563e-25, 
    -5.493967e-27, -4.285358e-25, 5.494132e-27, 4.395248e-26, 1.208692e-25, 
    8.515785e-26, 3.653544e-25, 2.417383e-25, -3.268959e-25, 1.730626e-25, 
    -4.202947e-25, -7.142256e-26, -8.515768e-26, -2.197612e-26, 2.829436e-25, 
    1.758097e-25, 9.06519e-26, 2.307502e-25, 3.159079e-25, 4.66995e-26, 
    -4.779822e-25, -2.554732e-25, -7.966364e-26, -1.565803e-25, 1.263632e-25, 
    -8.241066e-26, -2.637143e-25, -1.565803e-25, -3.076667e-25, 
    -1.648214e-25, 2.032799e-25, 1.703156e-25, -1.895446e-25, 1.922918e-25, 
    -5.65887e-25, -2.774494e-25, -3.296421e-26, 1.346043e-25, -2.747024e-25, 
    -2.856905e-25, -4.395231e-26, 2.719555e-25, -1.043869e-25, -4.120529e-26, 
    -4.093066e-25, -1.23616e-25, -2.554732e-25, -7.691661e-26, 3.818365e-25, 
    -4.175477e-25, 3.049198e-25, 2.582204e-25, 3.131609e-25, 3.18655e-25, 
    -5.219339e-26, -6.318148e-26, 2.225091e-25, 1.346043e-25, -2.197612e-26, 
    1.867978e-25, 5.027056e-25, -6.043446e-26, -2.060268e-25, 1.455924e-25, 
    -9.614578e-26, -1.950387e-25, -3.296421e-26, 3.351371e-25, 8.790487e-26, 
    -6.592851e-26, 2.637145e-25, -3.296421e-26, -1.758095e-25, -7.416958e-26, 
    2.939317e-25, -3.928245e-25, 8.241157e-27, 8.241083e-26, -1.703155e-25, 
    -4.669934e-26, -3.955715e-25, -1.840506e-25, -5.988513e-25, 1.291103e-25, 
    7.691677e-26, -4.889703e-25, -1.428452e-25, -5.466578e-25, 2.747107e-27, 
    -2.225089e-25, 2.225091e-25, -1.922909e-26, 2.08774e-25, 4.31283e-25, 
    -1.895446e-25, -3.296421e-26, 8.79048e-25, 1.922918e-25, -1.895446e-25, 
    -1.373504e-26, -7.416958e-26, 1.648223e-26, -1.648214e-25, 4.120545e-26, 
    2.389912e-25, 1.208692e-25, -4.395239e-25, 3.021735e-26, -1.016398e-25, 
    3.21402e-25, 4.395248e-26, 2.060269e-25, -5.219339e-26, 2.307502e-25, 
    5.219355e-26, 4.944653e-26, 5.384169e-25, -1.428452e-25, 2.197621e-25, 
    3.296438e-26, 3.378841e-25, 2.362442e-25, -2.719554e-25, -5.521519e-25, 
    8.257461e-32, -5.851162e-25, 1.346043e-25, -3.488721e-25, -1.593274e-25, 
    -2.911845e-25, -2.142679e-25, -3.46125e-25, -9.065174e-26, -4.202947e-25, 
    4.834764e-25, -5.493967e-27, 2.389912e-25, -1.675684e-25, -4.120536e-25, 
    4.944653e-26, -2.856905e-25, -1.538333e-25, 6.592867e-26, -3.845834e-25, 
    2.005329e-25, -1.950387e-25, -4.257888e-25, -7.334556e-25, -2.582203e-25, 
    1.483394e-25, -2.801964e-25, -1.977857e-25, 1.346043e-25, -1.071339e-25, 
    -1.538333e-25, -2.747024e-25, -6.043446e-26, -3.626072e-25, 
    -2.966786e-25, -4.340298e-25, -2.472314e-26, -1.043869e-25, 7.96638e-26, 
    -1.922909e-26, -4.285358e-25, 2.472323e-25, -3.818364e-25, -7.966364e-26, 
    2.637145e-25, 1.04387e-25, -6.592851e-26, -1.18122e-25, 3.433782e-25, 
    -4.340298e-25, 4.120538e-25, 4.944653e-26, 2.994258e-25, 2.856907e-25, 
    8.241157e-27, 2.582204e-25, -5.494041e-26, -3.516191e-25, -2.774494e-25, 
    1.126281e-25, 5.494132e-27, -8.241066e-26, 2.032799e-25, -4.752352e-25, 
    -2.087738e-25, 6.043463e-26, 8.241083e-26, -1.565803e-25, 2.939317e-25, 
    -3.104137e-25, -1.593274e-25, -3.955715e-25, 8.257467e-32, 3.845843e-26, 
    -3.516191e-25, 3.21402e-25, -1.620744e-25, -1.263631e-25, -4.175477e-25, 
    -1.867976e-25, -2.829435e-25, 2.747033e-26, -1.703155e-25, 4.395241e-25, 
    -1.620744e-25, -8.515768e-26, 8.790487e-26, -3.571124e-26, 1.098811e-25, 
    1.730626e-25, 1.208692e-25, 5.76876e-26, 4.3403e-25, 1.04387e-25, 
    -4.944636e-26, 2.362442e-25, -3.488721e-25, 3.461252e-25, -7.691661e-26, 
    -6.867554e-26, -4.312828e-25, -2.25256e-25, 2.032799e-25, -1.785565e-25, 
    -9.889281e-26, 1.181221e-25, -2.747024e-25, 3.159079e-25, -2.36244e-25, 
    -3.818364e-25, -3.735953e-25, -2.829435e-25, 1.977859e-25, -1.346041e-25, 
    -2.747024e-25, -2.527262e-25, 3.21402e-25, 1.922918e-25, 8.257297e-32, 
    -3.681012e-25, -1.977857e-25, 7.416975e-26, -1.950387e-25, -4.779822e-25, 
    1.181221e-25, 3.076668e-25, 4.587532e-25, 2.252561e-25, -2.389911e-25, 
    7.142273e-26, -1.098809e-25, -1.016398e-25, -1.126279e-25, 4.642473e-25, 
    -9.614578e-26, 2.197628e-26, 2.911847e-25, -4.50512e-25, -2.36244e-25, 
    2.11521e-25, 2.692085e-25, -2.554732e-25, -2.28003e-25, -3.571124e-26, 
    -1.593274e-25 ;

 M_LITR2C_TO_LEACHING =
  -1.15375e-25, -8.790474e-26, -8.515771e-26, -1.071339e-25, -1.428452e-25, 
    -2.527262e-25, 2.747078e-27, -7.966367e-26, 6.867567e-26, -1.483393e-25, 
    -4.944639e-26, 2.087739e-25, -7.416961e-26, 1.510864e-25, 1.758096e-25, 
    1.922923e-26, -1.922912e-26, 6.867567e-26, 4.120543e-26, -8.241021e-27, 
    -1.895447e-25, -9.339879e-26, 3.84584e-26, 1.07134e-25, -1.758095e-25, 
    4.669947e-26, -1.098805e-26, -1.758095e-25, 2.884376e-25, -9.339879e-26, 
    -1.867976e-25, -1.648209e-26, -1.291101e-25, -1.098809e-25, 
    -3.845829e-26, -6.318152e-26, -1.922912e-26, 3.021733e-26, 5.494055e-26, 
    -7.142259e-26, -7.691664e-26, -5.219342e-26, -1.510863e-25, 
    -2.472322e-25, -4.395234e-26, -1.12628e-25, 5.494055e-26, 3.021733e-26, 
    -1.895447e-25, -1.12628e-25, -3.076667e-25, 9.889295e-26, 1.620745e-25, 
    1.098815e-26, 5.494055e-26, -1.950387e-25, -4.120532e-26, 2.74703e-26, 
    -2.554732e-25, -5.493996e-27, -5.493996e-27, -1.318571e-25, 3.296435e-26, 
    -2.142679e-25, -2.115208e-25, -1.675685e-25, -4.120532e-26, 
    -2.197614e-26, 3.433782e-25, 4.94465e-26, 8.241128e-27, 1.09881e-25, 
    -3.296424e-26, 2.74703e-26, -2.774495e-25, 5.494103e-27, -3.461251e-25, 
    5.494055e-26, -9.889284e-26, 1.208691e-25, -6.592854e-26, -2.25256e-25, 
    -1.813036e-25, -1.098809e-25, -5.494044e-26, -2.142679e-25, 
    -5.219342e-26, -4.944639e-26, 6.592865e-26, 5.768757e-26, 1.098815e-26, 
    -1.098805e-26, -1.098805e-26, -1.400982e-25, -7.416961e-26, 3.296435e-26, 
    -1.236161e-25, 5.768757e-26, -1.648214e-25, 1.510864e-25, -2.362441e-25, 
    -5.494044e-26, 1.867977e-25, -9.339879e-26, 1.153751e-25, -1.12628e-25, 
    1.098815e-26, -5.494044e-26, -9.614581e-26, 8.241128e-27, 2.197625e-26, 
    -3.021727e-25, 1.153751e-25, -6.043449e-26, -8.790474e-26, -3.186548e-25, 
    -6.867557e-26, -3.049197e-25, -3.571127e-26, 1.318572e-25, 2.14268e-25, 
    -1.895447e-25, 1.922918e-25, -1.922912e-26, 2.307501e-25, -1.20869e-25, 
    -2.746971e-27, 8.241128e-27, -2.197614e-26, 1.813037e-25, 1.07134e-25, 
    3.296435e-26, 1.318572e-25, -2.499792e-25, 1.181221e-25, -4.944639e-26, 
    1.428453e-25, 2.692085e-25, -8.241069e-26, -1.428452e-25, -1.840506e-25, 
    1.620745e-25, 5.494055e-26, 3.735954e-25, -6.043449e-26, 3.296435e-26, 
    -1.098805e-26, 2.197625e-26, -8.241069e-26, 6.592865e-26, 1.922923e-26, 
    -1.098805e-26, 5.768757e-26, 5.768757e-26, -4.944639e-26, 1.675686e-25, 
    1.0164e-25, -2.3075e-25, -1.648209e-26, -6.592854e-26, 3.296435e-26, 
    2.307501e-25, -5.493996e-27, 3.296435e-26, -1.373507e-26, 5.494055e-26, 
    4.779824e-25, -6.043449e-26, -1.730625e-25, 1.04387e-25, -9.339879e-26, 
    -9.889284e-26, -1.071339e-25, 9.889295e-26, 1.840507e-25, -1.20869e-25, 
    -5.219342e-26, -1.098809e-25, 3.296435e-26, 1.703156e-25, 1.373513e-25, 
    -2.746971e-27, -2.637143e-25, 1.565805e-25, -8.241069e-26, -3.296424e-26, 
    1.098815e-26, -1.043869e-25, -1.098809e-25, 2.527263e-25, -3.845829e-26, 
    -7.691664e-26, 3.571138e-26, 6.592865e-26, -2.444852e-25, -3.571132e-25, 
    5.351449e-32, 6.04346e-26, 1.153751e-25, -1.867976e-25, -1.977857e-25, 
    1.181221e-25, -2.334971e-25, 1.758096e-25, 1.400983e-25, -5.494044e-26, 
    -2.692084e-25, -1.15375e-25, -1.20869e-25, -1.098805e-26, -2.746971e-27, 
    3.84584e-26, 8.241128e-27, -3.049197e-25, -5.493996e-27, -4.395234e-26, 
    2.472328e-26, -8.790474e-26, 1.153751e-25, -8.515771e-26, -2.087738e-25, 
    -1.236161e-25, 1.09881e-25, 1.04387e-25, -1.400982e-25, 1.620745e-25, 
    -9.339879e-26, 1.565805e-25, -2.197614e-26, -5.494044e-26, -4.395234e-26, 
    1.703156e-25, -3.571132e-25, -6.592854e-26, 1.922923e-26, 1.126281e-25, 
    -9.889284e-26, -6.592854e-26, -4.944639e-26, -9.339879e-26, 
    -9.339879e-26, -1.455923e-25, -1.016399e-25, -1.043869e-25, 
    -2.115208e-25, -1.043869e-25, -1.483393e-25, 1.181221e-25, 1.703156e-25, 
    -3.598602e-25, 3.84584e-26, 5.494055e-26, 1.098815e-26, -1.428452e-25, 
    1.538334e-25, -6.043449e-26, 1.181221e-25, -8.790474e-26, -1.373512e-25, 
    5.494055e-26, -1.483393e-25, -1.098805e-26, -4.395234e-26, 3.735954e-25, 
    4.94465e-26, 1.675686e-25, 1.538334e-25, 1.428453e-25, -2.142679e-25, 
    -3.461251e-25, 1.593275e-25, -3.845829e-26, 1.373513e-25, 4.120543e-26, 
    -1.483393e-25, -8.790474e-26, 5.351443e-32, -3.296424e-26, -4.395234e-26, 
    6.592865e-26, 2.74703e-26, -1.867976e-25, -1.483393e-25, -2.362441e-25, 
    4.148008e-25, -1.538333e-25, -1.565804e-25, 1.181221e-25, -3.735953e-25, 
    -3.845829e-26, -2.197614e-26, -8.790474e-26, 3.021733e-26, 9.889295e-26, 
    -3.845829e-26, -6.043449e-26, -8.515771e-26, 1.153751e-25, -1.098809e-25, 
    8.24108e-26, 1.483394e-25, 9.339889e-26, 2.692085e-25, 1.813037e-25, 
    -2.005328e-25, -2.25256e-25, -2.74702e-26, 2.19762e-25, -1.098805e-26, 
    -1.318571e-25, -3.818364e-25, -5.494044e-26, -1.620744e-25, 6.592865e-26, 
    2.362442e-25, 1.620745e-25, -2.417381e-25, -3.241489e-25, 1.922918e-25, 
    4.669947e-26, -1.922912e-26, -1.098809e-25, 5.494103e-27, -1.620744e-25, 
    1.09881e-25, -4.45018e-25, 1.153751e-25, 1.950388e-25, 1.538334e-25, 
    -2.197614e-26, -2.25256e-25, 3.928246e-25, -3.049197e-25, -2.472322e-25, 
    -1.400982e-25, -1.098805e-26, -1.840506e-25, 2.856906e-25 ;

 M_LITR3C_TO_LEACHING =
  1.291102e-25, 2.032799e-25, 2.747028e-26, 1.785569e-26, -1.263631e-25, 
    -3.983183e-26, 4.807296e-26, -1.071339e-25, -1.208691e-25, 1.332307e-25, 
    -5.906101e-26, -5.768749e-26, 2.675718e-32, 9.065185e-26, 3.708486e-26, 
    4.944647e-26, -1.483393e-25, 5.494052e-26, 1.428453e-25, -6.592857e-26, 
    -1.277366e-25, 1.400983e-25, 1.428453e-25, -4.395237e-26, 1.12628e-25, 
    1.236161e-25, -1.236161e-25, -6.318154e-26, -1.346042e-25, -1.71689e-25, 
    -5.494023e-27, -8.241047e-27, 2.060269e-25, 3.708486e-26, -6.043452e-26, 
    7.416969e-26, -3.57113e-26, -3.845832e-26, 9.614614e-27, 6.592862e-26, 
    1.167486e-25, 5.494076e-27, -1.37351e-26, -2.128944e-25, -1.098807e-26, 
    9.614614e-27, -1.085074e-25, -9.339881e-26, 2.197622e-26, -7.829018e-26, 
    -1.043869e-25, -1.291101e-25, 1.414718e-25, 5.494052e-26, -4.395237e-26, 
    -8.241071e-26, 4.944647e-26, 6.867565e-26, -4.120535e-26, -3.57113e-26, 
    -1.37351e-26, -2.060266e-26, -3.296427e-26, 7.966375e-26, -6.043452e-26, 
    -5.768749e-26, -9.614584e-26, 5.494052e-26, -1.112545e-25, -1.09881e-25, 
    -6.592857e-26, -1.510861e-26, -5.906101e-26, -2.334968e-26, 
    -1.414718e-25, -6.318154e-26, -7.279613e-26, 1.373515e-26, 1.510864e-25, 
    -4.395237e-26, -2.128944e-25, 8.241101e-27, -4.532588e-26, -4.120511e-27, 
    -1.09881e-25, -1.579539e-25, 4.532594e-26, -1.098807e-26, 2.747052e-27, 
    5.768755e-26, 1.236164e-26, 7.142267e-26, -1.318572e-25, -1.785563e-26, 
    -6.592857e-26, -8.515774e-26, -1.346042e-25, 8.241101e-27, 1.373515e-26, 
    -3.296427e-26, 3.02173e-26, 2.197622e-26, -8.653126e-26, 1.785569e-26, 
    -9.614584e-26, -1.167485e-25, -9.751935e-26, 3.845837e-26, -1.785563e-26, 
    -3.845832e-26, 1.07134e-25, -1.648212e-26, -6.592857e-26, -6.043452e-26, 
    8.241077e-26, 3.02173e-26, -7.142262e-26, 7.279618e-26, -1.510861e-26, 
    -1.304836e-25, -1.098807e-26, 2.884379e-26, 1.68942e-25, -8.790477e-26, 
    4.807296e-26, -3.296427e-26, -8.241047e-27, -2.183885e-25, -8.790477e-26, 
    -1.291101e-25, -1.098807e-26, 1.208691e-25, -1.346042e-25, 8.790482e-26, 
    -2.060266e-26, -8.653126e-26, -8.10372e-26, 1.648217e-26, 8.241101e-27, 
    6.592862e-26, -2.197617e-26, 6.867565e-26, -1.043869e-25, -1.37351e-26, 
    -2.22509e-25, -3.296427e-26, 3.571135e-26, -4.532588e-26, -1.236158e-26, 
    -1.208691e-25, -7.00491e-26, -9.20253e-26, -3.57113e-26, 6.592862e-26, 
    -1.112545e-25, 5.081998e-26, -1.236158e-26, -6.318154e-26, -1.002664e-25, 
    -2.884373e-26, -6.867535e-27, 5.356701e-26, -4.807291e-26, 3.433784e-26, 
    -4.120511e-27, -1.098807e-26, -7.279613e-26, -2.362441e-25, 
    -5.356696e-26, 8.927833e-26, 8.103726e-26, -2.747022e-26, 7.416969e-26, 
    9.614614e-27, -1.867977e-25, -1.140015e-25, -5.906101e-26, 6.867565e-26, 
    1.648217e-26, 2.675708e-32, -1.922915e-26, -1.785563e-26, 3.708486e-26, 
    -7.416964e-26, -4.944642e-26, -4.807291e-26, -8.653126e-26, 
    -5.906101e-26, 8.241101e-27, 1.648217e-26, 1.318572e-25, -6.867535e-27, 
    -5.219344e-26, 9.75194e-26, -5.768749e-26, 2.675723e-32, -2.747022e-26, 
    2.675726e-32, 3.571135e-26, 7.142267e-26, 4.395242e-26, 5.494052e-26, 
    -4.257886e-26, 5.356701e-26, -3.021725e-26, -1.428453e-25, -1.922915e-26, 
    -1.291101e-25, 1.098813e-26, -8.927828e-26, 3.571135e-26, 2.675721e-32, 
    -5.494023e-27, -8.241071e-26, 5.494076e-27, -1.648212e-26, 7.554321e-26, 
    -1.510863e-25, -5.219344e-26, 1.373515e-26, 5.356701e-26, -4.532588e-26, 
    -4.395237e-26, 1.153751e-25, -2.197617e-26, -1.332307e-25, -2.527263e-25, 
    -8.241047e-27, 8.103726e-26, -2.884373e-26, 3.845837e-26, -1.194956e-25, 
    -2.746998e-27, -6.043452e-26, -5.631398e-26, 2.675724e-32, -3.296427e-26, 
    7.142267e-26, 7.691672e-26, -3.845832e-26, -2.197617e-26, -2.060266e-26, 
    -3.296427e-26, 1.236161e-25, 7.554321e-26, 1.950388e-25, -5.768749e-26, 
    -8.515774e-26, 5.494076e-27, -6.867559e-26, -5.906101e-26, -5.494047e-26, 
    -1.37351e-26, -5.081993e-26, 3.02173e-26, 8.790482e-26, 1.483394e-25, 
    -5.768749e-26, -1.043869e-25, -1.565804e-25, 4.669945e-26, 2.675721e-32, 
    -1.15375e-25, -4.257886e-26, 4.532594e-26, -4.669939e-26, -5.494047e-26, 
    -4.257886e-26, -4.669939e-26, -3.983183e-26, -4.807291e-26, 
    -4.395237e-26, -1.359777e-25, 6.455511e-26, 2.747028e-26, -3.021725e-26, 
    -4.395237e-26, -3.845832e-26, 1.140016e-25, 9.889292e-26, 4.669945e-26, 
    -6.455506e-26, 8.241077e-26, 6.867589e-27, -3.296427e-26, 2.197622e-26, 
    6.31816e-26, -2.087739e-25, 4.944647e-26, 5.768755e-26, -5.494047e-26, 
    6.31816e-26, 4.12054e-26, 4.532594e-26, 7.279618e-26, 9.065185e-26, 
    -6.867559e-26, 3.02173e-26, -1.922915e-26, -2.884373e-26, -1.236158e-26, 
    5.21935e-26, 3.296432e-26, -1.318572e-25, 9.339887e-26, -2.884373e-26, 
    1.92292e-26, -1.400982e-25, 3.845837e-26, 2.197622e-26, -6.730208e-26, 
    -7.416964e-26, 3.845837e-26, 7.004916e-26, 6.043457e-26, -2.746998e-27, 
    1.002664e-25, 5.768755e-26, -1.043869e-25, -5.494023e-27, 2.307501e-25, 
    -1.346042e-25, 6.043457e-26, 1.648217e-26, -6.867535e-27, -7.416964e-26, 
    -4.120535e-26, -1.071339e-25, -2.47232e-26, -5.219344e-26, -1.648212e-26, 
    -1.648212e-26, -9.20253e-26, 8.653131e-26, -2.046533e-25, -8.241047e-27, 
    -1.236158e-26, -1.15375e-25 ;

 M_SOIL1C_TO_LEACHING =
  2.751366e-20, 5.717381e-21, -1.131751e-21, -7.471725e-21, 1.108026e-21, 
    -4.213791e-20, -4.400816e-20, -1.00703e-20, 1.885191e-20, 1.257867e-21, 
    -2.457438e-20, 1.463754e-20, -6.327817e-21, -1.392366e-20, 1.667715e-20, 
    -1.002423e-20, 8.377319e-21, -1.336299e-20, -2.471547e-20, 8.481635e-21, 
    1.095864e-20, -1.688949e-20, 1.148171e-20, 1.924208e-20, 3.074017e-20, 
    4.103567e-21, 2.694934e-20, 4.328635e-22, 1.693758e-20, -2.453285e-20, 
    1.035416e-20, 7.783292e-21, 2.495412e-20, 2.459503e-20, 3.343317e-21, 
    -9.825767e-21, 3.654802e-20, -8.315957e-21, -2.168064e-20, -2.305074e-20, 
    -1.030584e-20, 1.362745e-21, -1.294397e-20, 3.551183e-20, 1.113988e-20, 
    -1.174491e-20, 5.214133e-21, -6.572085e-21, -4.678334e-21, 1.45708e-20, 
    2.136116e-20, 1.57761e-20, -6.575743e-21, 7.81168e-22, -2.755493e-21, 
    6.517707e-20, -4.886981e-21, -1.797292e-20, -2.319524e-20, 2.551916e-21, 
    -3.783616e-20, -5.549735e-21, 3.009951e-20, 4.989236e-20, 1.474695e-20, 
    -2.039394e-20, 5.92027e-22, 2.224721e-20, -3.590088e-20, -4.769374e-21, 
    1.833848e-20, -1.701389e-20, 7.355793e-21, -2.242989e-20, -2.299307e-20, 
    2.95992e-21, 4.114017e-21, 1.705236e-20, -2.387518e-20, -7.06769e-21, 
    -3.626391e-20, 2.482998e-20, -9.124002e-21, 5.624079e-21, 1.340115e-20, 
    2.204157e-21, -1.518309e-22, -1.006011e-20, 4.894067e-21, -2.33434e-20, 
    7.315665e-21, -7.777634e-21, -9.228627e-21, -2.07864e-21, 5.388572e-21, 
    1.630705e-20, 1.115544e-20, 2.275161e-20, 3.463084e-20, 2.207026e-20, 
    4.875949e-20, -1.721596e-22, -1.209834e-20, -4.514084e-21, 5.517773e-21, 
    5.464677e-20, 1.21283e-20, 1.818665e-20, 6.300386e-21, -9.646199e-21, 
    -3.053266e-20, -2.671239e-21, 2.860839e-20, -4.857875e-21, -3.64505e-20, 
    1.62867e-20, 2.960475e-20, 4.120516e-21, 9.107624e-21, -1.402683e-20, 
    8.395697e-21, 1.897632e-20, -2.374909e-20, -2.186697e-20, 3.052078e-20, 
    -4.12487e-20, -3.782933e-22, 7.363704e-21, 2.032579e-20, 2.574602e-20, 
    3.544961e-20, 1.932154e-20, 3.729331e-20, 2.016152e-20, -4.435877e-20, 
    -2.4599e-20, 4.588716e-21, 2.149122e-20, -3.885009e-21, 2.624318e-21, 
    -1.098577e-20, -1.125841e-21, 4.362196e-20, 7.503967e-21, 2.011009e-20, 
    8.967379e-21, -2.209683e-20, -6.716561e-21, -3.106872e-20, 1.081303e-20, 
    3.342613e-20, -4.505343e-20, 1.627851e-20, -4.45298e-20, -6.407787e-21, 
    -1.965826e-21, 4.170555e-21, 4.869698e-20, -1.296349e-20, -2.116438e-20, 
    -2.301145e-20, -2.975686e-20, -1.459654e-20, -1.156654e-21, 
    -1.778629e-20, -5.750943e-20, 4.022297e-20, 2.007945e-21, 4.205084e-20, 
    1.714452e-20, -3.129915e-20, -3.647821e-20, -2.595103e-20, -1.479249e-20, 
    -2.119123e-20, -5.595234e-21, 3.33922e-20, -7.241011e-21, 5.104715e-21, 
    -1.818183e-20, -1.763223e-20, -6.11379e-21, -7.322728e-22, 7.354397e-21, 
    3.907617e-21, -2.622583e-20, -1.265784e-20, 1.09903e-20, 2.523344e-20, 
    -1.840267e-20, 2.40454e-20, -1.007655e-20, -2.195122e-20, -1.206497e-20, 
    -1.371132e-20, 2.899518e-20, 1.526266e-20, 1.297162e-21, 8.152253e-21, 
    2.539629e-20, 5.00885e-21, 7.970744e-21, 2.812493e-20, -4.074942e-20, 
    -5.663154e-20, -1.360755e-20, -3.562136e-21, -3.788166e-20, -7.59983e-22, 
    1.420752e-20, 3.897166e-21, -9.544163e-21, 1.298724e-20, -3.48491e-20, 
    -1.522987e-20, 7.799418e-21, -1.62101e-20, -1.237426e-20, -3.108595e-20, 
    1.351283e-20, 6.251337e-22, -2.620123e-20, 2.615003e-20, -8.087494e-21, 
    1.011017e-20, 1.176556e-20, 1.785927e-20, -1.595872e-20, 8.869855e-21, 
    2.227466e-20, -8.267099e-22, 4.021647e-20, -3.626417e-20, 1.539241e-20, 
    4.812948e-21, -2.549974e-21, -1.366297e-20, -6.397084e-21, 2.153251e-20, 
    1.860963e-20, 3.711887e-20, -2.640197e-20, 1.034146e-20, 2.89751e-20, 
    6.086914e-21, -1.248482e-20, 5.138689e-20, -2.466345e-20, -9.666283e-21, 
    -1.186988e-20, 3.049254e-21, 9.275549e-21, 5.913593e-21, -3.390112e-20, 
    3.60575e-20, 3.603205e-20, -2.699341e-20, 2.103714e-20, -3.054541e-20, 
    -1.232648e-20, 1.837353e-20, -2.103829e-20, 4.736646e-20, -2.478135e-21, 
    -4.093378e-21, -1.703792e-20, -2.864911e-21, -1.414955e-20, 
    -2.643616e-20, 3.475037e-21, 4.119866e-20, 2.160093e-20, 2.234927e-20, 
    -3.221799e-20, -1.561521e-20, 1.309607e-20, -9.418619e-21, 3.479485e-20, 
    3.021346e-20, 1.907133e-20, 1.285353e-20, -1.086023e-20, 2.870171e-20, 
    -3.503798e-20, -1.684085e-20, 2.408583e-20, 3.373089e-22, 2.884673e-20, 
    -1.598221e-20, -1.439297e-20, 3.547732e-20, 1.692059e-20, -1.038047e-20, 
    2.245447e-20, 1.101547e-20, 2.705652e-22, 2.629452e-20, 6.911345e-21, 
    2.830276e-20, -1.812418e-20, 2.394149e-21, -5.991905e-21, 2.566352e-21, 
    -2.25263e-20, -2.535539e-21, 9.360064e-21, 3.254656e-20, 7.208215e-21, 
    6.822011e-21, 3.374952e-21, 5.151375e-21, 2.528235e-20, 2.106515e-20, 
    -1.341134e-20, 1.381789e-20, -2.669833e-21, 3.697279e-21, -3.524238e-20, 
    1.81598e-20, 1.162616e-20, 8.250086e-21, -3.128188e-20, -2.225957e-21, 
    1.971199e-20, 4.024107e-20, -8.069973e-21, -9.794088e-21, -1.594827e-20, 
    -1.038357e-20, -2.133912e-20, -1.078787e-20, -1.293887e-20, 4.746195e-21, 
    1.84086e-20, 2.298205e-20, -2.686141e-20, 1.769779e-20, -4.102395e-20 ;

 M_SOIL2C_TO_LEACHING =
  2.031223e-20, -2.538442e-20, 2.515173e-20, 3.857974e-20, 1.386824e-20, 
    4.764692e-20, 9.999606e-21, -9.368018e-21, 1.659064e-20, -2.071568e-20, 
    2.078665e-20, -1.067303e-21, 8.698503e-21, 1.962774e-20, 1.001404e-20, 
    8.006097e-21, 2.045217e-20, 1.746171e-20, -2.950294e-20, 3.694739e-21, 
    6.948673e-21, 1.539977e-20, 4.684707e-20, -3.195876e-20, 1.095637e-20, 
    -2.325572e-20, -1.691013e-20, 5.379462e-20, 2.41367e-21, 1.21266e-20, 
    -2.865562e-20, -2.527442e-20, 1.5812e-20, -1.801392e-20, 7.738601e-21, 
    -6.688557e-21, 2.001791e-20, 3.578235e-21, -1.411308e-20, -4.424597e-20, 
    1.890423e-20, 3.563058e-20, 4.260478e-21, -1.733394e-20, -6.104174e-21, 
    1.403447e-20, 4.730453e-20, -1.020969e-20, 4.286766e-21, 1.530365e-20, 
    -2.292354e-20, -2.924623e-20, 1.275059e-20, 4.094281e-20, 2.557244e-20, 
    -1.367682e-20, -2.076291e-20, 8.955221e-21, -3.685401e-21, -5.274067e-21, 
    -5.794003e-21, 4.559429e-20, -3.925434e-20, 5.149096e-21, 8.35837e-21, 
    -4.231489e-20, -4.86133e-20, -9.988696e-22, 1.473139e-20, -5.703501e-20, 
    -9.819258e-21, -8.664278e-21, -2.127069e-20, 1.72135e-20, 1.75997e-20, 
    1.958984e-20, 2.025188e-21, 1.388858e-20, -8.103904e-21, 1.347353e-20, 
    -8.321043e-21, 2.371258e-21, -1.67467e-20, -1.532542e-20, -1.657989e-20, 
    -2.432417e-20, -8.621015e-21, -9.252663e-21, -1.56873e-20, -1.379643e-20, 
    -2.246466e-20, -2.44206e-20, -3.912719e-21, 3.059853e-20, -1.684511e-20, 
    -1.288632e-20, -1.820194e-20, 2.869141e-21, -1.49836e-20, -3.401957e-20, 
    3.080918e-20, -2.013806e-20, -2.422494e-20, -1.278678e-20, 2.809498e-20, 
    7.959437e-21, -4.860708e-20, -1.207316e-20, -2.697527e-21, -3.142864e-20, 
    -2.251074e-20, 1.690276e-20, 9.01007e-21, 1.831228e-21, -1.606985e-20, 
    -1.48632e-21, 2.191898e-20, -2.658603e-20, 2.618114e-20, -4.042767e-20, 
    -4.419591e-20, 1.965545e-20, 1.12391e-20, -3.04764e-20, -9.477964e-21, 
    -6.729836e-21, 1.114579e-20, 7.027556e-21, 1.85398e-20, 3.580391e-20, 
    8.677302e-21, 6.401043e-21, 2.432391e-20, 3.269327e-20, -1.326687e-20, 
    -2.70121e-20, 2.003486e-20, -3.460082e-21, -2.557329e-20, 3.9273e-20, 
    3.104959e-21, -1.349956e-20, 3.673096e-20, 1.138981e-20, 7.959437e-21, 
    5.749344e-21, -4.044265e-20, 1.986721e-20, -1.258123e-20, 3.047156e-20, 
    9.897832e-21, -2.908394e-20, -8.497188e-21, -4.161287e-20, 3.763824e-20, 
    -2.853828e-20, 2.699033e-20, -5.944471e-20, 2.185396e-20, -4.807639e-20, 
    -4.412183e-20, -7.353253e-21, -1.354733e-20, -2.828269e-20, 
    -2.579947e-20, 1.240169e-20, 1.199257e-20, -1.286509e-20, -1.010395e-20, 
    7.42083e-21, -5.009989e-20, -1.234743e-20, -1.359114e-20, 2.705366e-20, 
    -4.445149e-20, -1.152723e-20, 5.596603e-23, 2.242198e-20, 5.297531e-21, 
    -1.896756e-20, 3.728766e-20, -4.653013e-20, -2.871965e-21, 1.188883e-20, 
    1.994671e-21, -1.301777e-20, -5.453019e-21, -3.506715e-21, -1.432202e-20, 
    1.939053e-20, -2.452434e-20, -2.890837e-20, -1.587024e-20, -3.742778e-21, 
    -2.885523e-20, 7.620733e-21, -3.81715e-20, -9.64423e-21, 5.733245e-21, 
    5.475082e-21, 1.421374e-20, 1.578089e-20, -1.344414e-20, -2.569741e-20, 
    -2.129783e-20, 1.228012e-20, -2.186526e-20, -1.568928e-20, 4.131884e-20, 
    -2.227127e-20, 4.665986e-23, -2.434765e-20, 1.477071e-20, 2.589815e-21, 
    1.152975e-20, 3.321437e-20, -1.46415e-20, -1.444302e-20, -7.795449e-21, 
    -1.064878e-20, -1.419308e-20, 9.287989e-21, 2.882158e-20, 1.605884e-20, 
    -1.807131e-20, 1.989096e-20, -3.772252e-20, -2.516898e-20, 1.91471e-20, 
    -1.60628e-20, 5.913511e-20, -1.238673e-20, -1.508652e-20, -1.862404e-20, 
    1.306102e-20, -2.161959e-20, -3.965016e-20, -9.822916e-21, -3.759132e-20, 
    -2.255316e-20, -1.028152e-20, 1.709108e-20, -5.971698e-20, 1.753751e-20, 
    1.238656e-21, -1.42157e-20, 1.360078e-20, 1.212605e-20, 2.30697e-20, 
    8.209364e-21, -4.867664e-20, 3.387959e-21, -5.680338e-21, -9.925263e-21, 
    2.588766e-20, 4.349524e-21, 1.120912e-20, 3.576289e-20, -6.658595e-21, 
    -1.145991e-20, 4.355468e-20, -2.625436e-21, 4.198584e-20, -8.873513e-21, 
    -4.025859e-20, -3.672163e-20, -1.296914e-20, -1.99031e-20, -2.936216e-20, 
    4.448502e-21, -5.805649e-20, -1.199145e-20, -2.750979e-21, -9.276094e-21, 
    -7.390654e-22, -1.207716e-20, 9.611697e-21, -9.06718e-21, 1.978639e-20, 
    -1.291795e-20, -2.60378e-20, -3.440976e-20, -7.684913e-21, 3.337608e-20, 
    -1.564829e-20, -1.379303e-20, 3.803152e-20, -4.263071e-20, 8.023962e-22, 
    -2.875768e-20, 1.714226e-20, 2.44777e-20, 2.801581e-21, -4.010931e-20, 
    -2.771384e-20, -1.159478e-20, 1.17896e-20, -2.391339e-20, -5.848573e-21, 
    -1.893533e-20, -2.257238e-20, 1.422929e-20, -9.27358e-21, 1.046415e-20, 
    -9.860815e-21, -2.222828e-20, 7.464933e-21, 1.764748e-20, 2.652184e-20, 
    1.976007e-20, 3.065312e-20, 8.954649e-21, -1.212913e-21, -2.947453e-21, 
    -6.431839e-21, -2.487436e-20, 3.00164e-20, -1.419875e-20, -7.08531e-22, 
    -6.712047e-21, -1.934728e-20, 6.172591e-21, -1.283232e-20, 3.69778e-20, 
    -3.134806e-20, 1.380517e-20, 2.985593e-22, -2.27166e-20, -2.88993e-20, 
    8.015404e-21, -2.796433e-20, -3.14261e-20, 8.006669e-21, 2.032891e-20, 
    -3.097737e-20, -4.083567e-20, -3.689495e-20, 1.273731e-20 ;

 M_SOIL3C_TO_LEACHING =
  2.017028e-20, 2.545114e-20, 7.843243e-21, 6.710886e-21, -4.062843e-21, 
    8.019944e-21, 2.631799e-20, -7.725327e-21, -3.890277e-22, -4.361992e-21, 
    2.74147e-20, 2.063537e-20, -5.494593e-21, -1.632714e-20, 7.927197e-21, 
    2.823095e-20, 3.469589e-20, 2.406351e-20, -2.817638e-20, 3.340605e-20, 
    -2.827451e-20, -7.396375e-22, 1.769725e-20, 3.10591e-20, -2.338466e-20, 
    -1.438648e-20, -2.268179e-20, -8.190837e-22, 1.200618e-20, -2.348758e-20, 
    -1.346957e-20, 4.379614e-20, 5.974751e-20, -1.326855e-20, -1.603762e-20, 
    1.029676e-20, -3.97605e-21, -2.955497e-20, 6.847654e-20, 2.823943e-20, 
    1.774049e-20, 3.258195e-21, 1.741282e-20, 1.577916e-21, -1.943095e-20, 
    1.720692e-21, 1.884117e-20, 1.279245e-20, 3.526981e-20, 2.991349e-20, 
    2.085535e-20, -6.173414e-21, -1.012175e-20, -5.216252e-22, -4.652902e-21, 
    -3.814858e-20, 3.264496e-20, 6.546065e-21, -2.501657e-20, 9.087247e-21, 
    -2.661966e-20, -4.640745e-21, 9.38495e-21, -6.793928e-22, -3.540335e-21, 
    5.361e-20, -8.414646e-21, 1.500255e-20, -2.362158e-20, -1.592115e-20, 
    -6.925503e-21, 3.723845e-21, -3.322625e-20, -1.41798e-20, 2.610161e-21, 
    -6.544947e-21, -1.828705e-20, 1.055718e-21, 2.402789e-20, 6.469149e-21, 
    -7.676977e-21, 8.067721e-21, 3.458308e-20, -2.387097e-20, -1.293409e-20, 
    -4.384728e-20, -7.89271e-21, -2.824498e-21, -2.747324e-20, 6.334048e-20, 
    -5.550853e-21, 2.806388e-20, -2.411693e-20, -1.594827e-20, -2.421109e-20, 
    3.563254e-21, 1.057979e-20, -6.599778e-21, 2.550628e-20, -1.579901e-20, 
    9.050204e-21, -3.094797e-20, 1.362538e-20, -2.157801e-20, 1.578317e-20, 
    6.378681e-21, 2.515992e-20, -7.140942e-21, 4.422188e-21, -8.013151e-21, 
    -1.686403e-20, 2.667482e-20, -1.6734e-20, -1.377805e-20, 1.58971e-20, 
    1.316959e-20, -2.205074e-20, -3.435291e-22, -3.21332e-20, -6.31366e-21, 
    -3.648978e-20, 3.334782e-20, 2.479718e-20, 7.178252e-21, -1.831474e-20, 
    -1.61654e-20, 8.146605e-21, 3.852213e-21, -1.766249e-20, 1.979878e-20, 
    -2.790846e-21, -3.125251e-20, -1.859633e-20, 6.668212e-21, -3.505013e-20, 
    -1.260783e-20, 1.450386e-22, -1.617502e-20, 4.768802e-21, -1.253485e-20, 
    -1.761448e-22, -1.161995e-20, 2.184384e-21, 1.805914e-20, -4.408933e-20, 
    3.582173e-20, -1.733206e-22, 1.705405e-20, -6.667838e-20, -4.196434e-20, 
    8.913926e-21, -2.467392e-20, 4.906821e-20, 9.957487e-21, -2.830504e-20, 
    9.164441e-21, 2.21549e-21, 4.053244e-21, -5.749033e-21, -2.389752e-20, 
    -1.002649e-20, 2.072966e-21, 1.684793e-20, 7.738911e-21, 6.820011e-21, 
    -2.571438e-21, 4.292702e-21, 1.198438e-20, 3.063783e-20, -4.309807e-20, 
    -2.03651e-20, 1.966761e-20, 7.946735e-21, 2.584451e-21, 2.211747e-20, 
    1.768143e-20, -2.920071e-20, 1.272848e-21, -8.123425e-21, -9.548676e-21, 
    1.71021e-20, 2.020564e-20, -4.996693e-21, -4.715661e-21, 2.513756e-21, 
    -4.093998e-22, -3.639227e-20, -1.697402e-20, 1.752675e-20, 1.077799e-20, 
    5.908507e-21, -4.075e-21, -9.626132e-21, 3.879906e-21, -7.458141e-21, 
    -1.009832e-20, 3.47465e-20, -4.313904e-21, -1.003977e-20, 2.514807e-20, 
    6.387174e-21, -6.325817e-21, 2.341745e-20, 2.941558e-20, 4.124051e-20, 
    7.749907e-20, -2.453567e-20, -7.045627e-22, 2.084065e-20, 1.948949e-20, 
    -3.788845e-20, 1.308619e-20, -1.427198e-20, 1.412635e-20, -1.210796e-20, 
    5.693067e-21, -1.647777e-21, 2.007048e-20, -3.021798e-20, 3.264416e-21, 
    -1.430615e-21, 2.210134e-20, 6.339664e-21, -2.087855e-20, -1.782627e-21, 
    -2.940452e-22, 6.314233e-21, -3.13342e-20, 4.115655e-20, -7.812137e-21, 
    1.106976e-20, 4.949226e-21, -1.84154e-20, -1.052322e-21, -2.267226e-21, 
    7.130754e-21, 1.744621e-20, -2.890075e-20, 4.37246e-20, -9.88316e-21, 
    -4.578549e-21, -1.2536e-20, -1.385183e-20, 1.748098e-20, 1.757399e-20, 
    1.444414e-20, -1.476535e-20, 2.034303e-20, 2.263826e-20, 2.03648e-20, 
    9.041159e-21, 2.310192e-20, 1.189744e-21, -1.892714e-20, -1.802972e-21, 
    -1.839023e-20, -8.843655e-22, -3.429269e-20, -1.210822e-20, 
    -3.404219e-20, -7.952644e-21, 2.459186e-21, 1.64278e-20, 1.041872e-21, 
    1.234036e-20, 1.478393e-21, -6.781026e-21, 2.549403e-21, 7.62329e-21, 
    3.607531e-20, -1.53353e-20, -1.71889e-20, 3.076114e-21, 2.163745e-21, 
    -1.245514e-20, 7.331506e-21, 3.236928e-20, -8.520079e-21, 3.123525e-20, 
    1.475205e-20, 1.016474e-20, 3.203765e-20, -1.147209e-20, 1.830908e-20, 
    2.714301e-20, -2.333669e-21, 3.088833e-21, 2.285765e-20, 8.979535e-21, 
    1.787594e-20, -1.412072e-20, 5.357465e-21, 1.316847e-20, 2.166907e-20, 
    2.22034e-20, 1.739642e-21, 9.184508e-21, 1.676055e-20, 1.307431e-20, 
    1.684002e-20, 7.695076e-21, -4.073584e-20, -2.949453e-21, -2.682665e-20, 
    -9.064328e-21, 4.995559e-21, -3.483412e-20, -3.341906e-20, 1.575082e-21, 
    -3.300288e-21, 3.609603e-21, -2.847722e-20, 3.64102e-21, 2.300385e-20, 
    7.287098e-21, 1.216958e-20, 7.917318e-21, 5.315052e-21, -2.265918e-20, 
    2.808591e-20, 3.529047e-20, -2.049401e-20, 1.702973e-20, -8.287086e-21, 
    2.206233e-20, -9.841293e-21, -1.953048e-20, -1.181643e-20, -8.870117e-21, 
    -2.319578e-20, -6.359185e-21, -1.392138e-20, 2.101397e-20, 5.553132e-21, 
    7.547214e-21, 3.321437e-20, -2.504571e-20, -3.902363e-20 ;

 NBP =
  -6.356978e-08, -6.384934e-08, -6.379499e-08, -6.402048e-08, -6.389539e-08, 
    -6.404304e-08, -6.362645e-08, -6.386044e-08, -6.371106e-08, 
    -6.359494e-08, -6.445807e-08, -6.403054e-08, -6.490213e-08, 
    -6.462948e-08, -6.531439e-08, -6.485971e-08, -6.540607e-08, 
    -6.530126e-08, -6.561668e-08, -6.552632e-08, -6.592977e-08, 
    -6.565838e-08, -6.61389e-08, -6.586495e-08, -6.590781e-08, -6.564943e-08, 
    -6.411657e-08, -6.440485e-08, -6.409949e-08, -6.41406e-08, -6.412215e-08, 
    -6.389798e-08, -6.378502e-08, -6.354841e-08, -6.359136e-08, 
    -6.376514e-08, -6.415908e-08, -6.402535e-08, -6.436237e-08, 
    -6.435476e-08, -6.472996e-08, -6.456079e-08, -6.51914e-08, -6.501217e-08, 
    -6.553009e-08, -6.539984e-08, -6.552398e-08, -6.548633e-08, 
    -6.552447e-08, -6.533344e-08, -6.541529e-08, -6.524719e-08, 
    -6.459248e-08, -6.478489e-08, -6.421101e-08, -6.386593e-08, 
    -6.363672e-08, -6.347406e-08, -6.349706e-08, -6.35409e-08, -6.376616e-08, 
    -6.397794e-08, -6.413933e-08, -6.42473e-08, -6.435366e-08, -6.467567e-08, 
    -6.484608e-08, -6.522765e-08, -6.515878e-08, -6.527544e-08, 
    -6.538689e-08, -6.557399e-08, -6.55432e-08, -6.562563e-08, -6.527236e-08, 
    -6.550714e-08, -6.511956e-08, -6.522556e-08, -6.438261e-08, 
    -6.406143e-08, -6.392494e-08, -6.380544e-08, -6.351474e-08, 
    -6.371549e-08, -6.363636e-08, -6.382462e-08, -6.394425e-08, 
    -6.388508e-08, -6.425024e-08, -6.410828e-08, -6.485618e-08, 
    -6.453404e-08, -6.537388e-08, -6.517291e-08, -6.542206e-08, 
    -6.529492e-08, -6.551276e-08, -6.53167e-08, -6.565631e-08, -6.573026e-08, 
    -6.567973e-08, -6.587384e-08, -6.530584e-08, -6.552398e-08, 
    -6.388343e-08, -6.389308e-08, -6.393803e-08, -6.374042e-08, 
    -6.372833e-08, -6.354723e-08, -6.370837e-08, -6.377699e-08, 
    -6.395118e-08, -6.405422e-08, -6.415217e-08, -6.436752e-08, 
    -6.460803e-08, -6.494434e-08, -6.518594e-08, -6.53479e-08, -6.524859e-08, 
    -6.533626e-08, -6.523825e-08, -6.519231e-08, -6.570255e-08, 
    -6.541605e-08, -6.584592e-08, -6.582213e-08, -6.562759e-08, 
    -6.582481e-08, -6.389985e-08, -6.384432e-08, -6.365153e-08, -6.38024e-08, 
    -6.352751e-08, -6.368138e-08, -6.376987e-08, -6.411125e-08, 
    -6.418625e-08, -6.425581e-08, -6.439316e-08, -6.456945e-08, 
    -6.487869e-08, -6.514775e-08, -6.539337e-08, -6.537537e-08, 
    -6.538171e-08, -6.543657e-08, -6.530066e-08, -6.545889e-08, 
    -6.548544e-08, -6.541601e-08, -6.581894e-08, -6.570383e-08, 
    -6.582162e-08, -6.574668e-08, -6.386237e-08, -6.395581e-08, 
    -6.390532e-08, -6.400027e-08, -6.393338e-08, -6.42308e-08, -6.431998e-08, 
    -6.473723e-08, -6.456598e-08, -6.483852e-08, -6.459366e-08, 
    -6.463705e-08, -6.484741e-08, -6.460689e-08, -6.513292e-08, -6.47763e-08, 
    -6.543871e-08, -6.50826e-08, -6.546102e-08, -6.53923e-08, -6.550608e-08, 
    -6.560798e-08, -6.573618e-08, -6.597273e-08, -6.591795e-08, 
    -6.611577e-08, -6.40951e-08, -6.42163e-08, -6.420562e-08, -6.433245e-08, 
    -6.442625e-08, -6.462955e-08, -6.49556e-08, -6.483299e-08, -6.505808e-08, 
    -6.510327e-08, -6.476129e-08, -6.497127e-08, -6.42974e-08, -6.440629e-08, 
    -6.434146e-08, -6.410467e-08, -6.486125e-08, -6.447298e-08, 
    -6.518994e-08, -6.49796e-08, -6.559345e-08, -6.528818e-08, -6.58878e-08, 
    -6.614415e-08, -6.638538e-08, -6.666732e-08, -6.428244e-08, 
    -6.420009e-08, -6.434753e-08, -6.455154e-08, -6.47408e-08, -6.499243e-08, 
    -6.501818e-08, -6.506531e-08, -6.518741e-08, -6.529008e-08, 
    -6.508023e-08, -6.531582e-08, -6.443155e-08, -6.489495e-08, 
    -6.416896e-08, -6.438758e-08, -6.453951e-08, -6.447286e-08, 
    -6.481897e-08, -6.490055e-08, -6.523204e-08, -6.506068e-08, 
    -6.608088e-08, -6.562952e-08, -6.688197e-08, -6.653197e-08, 
    -6.417132e-08, -6.428215e-08, -6.466789e-08, -6.448436e-08, 
    -6.500922e-08, -6.513842e-08, -6.524344e-08, -6.53777e-08, -6.539219e-08, 
    -6.547174e-08, -6.534139e-08, -6.546659e-08, -6.499297e-08, 
    -6.520462e-08, -6.46238e-08, -6.476517e-08, -6.470013e-08, -6.46288e-08, 
    -6.484896e-08, -6.508353e-08, -6.508854e-08, -6.516375e-08, 
    -6.537572e-08, -6.501136e-08, -6.613915e-08, -6.544267e-08, 
    -6.440301e-08, -6.461651e-08, -6.464699e-08, -6.456429e-08, 
    -6.512547e-08, -6.492213e-08, -6.54698e-08, -6.532179e-08, -6.55643e-08, 
    -6.544379e-08, -6.542606e-08, -6.527128e-08, -6.517492e-08, 
    -6.493146e-08, -6.473337e-08, -6.457628e-08, -6.461281e-08, 
    -6.478536e-08, -6.509788e-08, -6.539351e-08, -6.532875e-08, 
    -6.554587e-08, -6.497117e-08, -6.521216e-08, -6.511902e-08, 
    -6.536187e-08, -6.482973e-08, -6.52829e-08, -6.471389e-08, -6.476378e-08, 
    -6.49181e-08, -6.522851e-08, -6.529717e-08, -6.53705e-08, -6.532525e-08, 
    -6.510581e-08, -6.506986e-08, -6.491435e-08, -6.487141e-08, 
    -6.475292e-08, -6.465483e-08, -6.474446e-08, -6.483858e-08, -6.51059e-08, 
    -6.53468e-08, -6.560944e-08, -6.567371e-08, -6.59806e-08, -6.573079e-08, 
    -6.614304e-08, -6.579257e-08, -6.639924e-08, -6.530915e-08, 
    -6.578225e-08, -6.492512e-08, -6.501746e-08, -6.518448e-08, 
    -6.556754e-08, -6.536073e-08, -6.560259e-08, -6.506844e-08, 
    -6.479132e-08, -6.471961e-08, -6.458583e-08, -6.472267e-08, 
    -6.471154e-08, -6.484247e-08, -6.48004e-08, -6.511478e-08, -6.494591e-08, 
    -6.542562e-08, -6.560068e-08, -6.609504e-08, -6.63981e-08, -6.670659e-08, 
    -6.684278e-08, -6.688423e-08, -6.690156e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.356978e-08, 6.384934e-08, 6.379499e-08, 6.402048e-08, 6.389539e-08, 
    6.404304e-08, 6.362645e-08, 6.386044e-08, 6.371106e-08, 6.359494e-08, 
    6.445807e-08, 6.403054e-08, 6.490213e-08, 6.462948e-08, 6.531439e-08, 
    6.485971e-08, 6.540607e-08, 6.530126e-08, 6.561668e-08, 6.552632e-08, 
    6.592977e-08, 6.565838e-08, 6.61389e-08, 6.586495e-08, 6.590781e-08, 
    6.564943e-08, 6.411657e-08, 6.440485e-08, 6.409949e-08, 6.41406e-08, 
    6.412215e-08, 6.389798e-08, 6.378502e-08, 6.354841e-08, 6.359136e-08, 
    6.376514e-08, 6.415908e-08, 6.402535e-08, 6.436237e-08, 6.435476e-08, 
    6.472996e-08, 6.456079e-08, 6.51914e-08, 6.501217e-08, 6.553009e-08, 
    6.539984e-08, 6.552398e-08, 6.548633e-08, 6.552447e-08, 6.533344e-08, 
    6.541529e-08, 6.524719e-08, 6.459248e-08, 6.478489e-08, 6.421101e-08, 
    6.386593e-08, 6.363672e-08, 6.347406e-08, 6.349706e-08, 6.35409e-08, 
    6.376616e-08, 6.397794e-08, 6.413933e-08, 6.42473e-08, 6.435366e-08, 
    6.467567e-08, 6.484608e-08, 6.522765e-08, 6.515878e-08, 6.527544e-08, 
    6.538689e-08, 6.557399e-08, 6.55432e-08, 6.562563e-08, 6.527236e-08, 
    6.550714e-08, 6.511956e-08, 6.522556e-08, 6.438261e-08, 6.406143e-08, 
    6.392494e-08, 6.380544e-08, 6.351474e-08, 6.371549e-08, 6.363636e-08, 
    6.382462e-08, 6.394425e-08, 6.388508e-08, 6.425024e-08, 6.410828e-08, 
    6.485618e-08, 6.453404e-08, 6.537388e-08, 6.517291e-08, 6.542206e-08, 
    6.529492e-08, 6.551276e-08, 6.53167e-08, 6.565631e-08, 6.573026e-08, 
    6.567973e-08, 6.587384e-08, 6.530584e-08, 6.552398e-08, 6.388343e-08, 
    6.389308e-08, 6.393803e-08, 6.374042e-08, 6.372833e-08, 6.354723e-08, 
    6.370837e-08, 6.377699e-08, 6.395118e-08, 6.405422e-08, 6.415217e-08, 
    6.436752e-08, 6.460803e-08, 6.494434e-08, 6.518594e-08, 6.53479e-08, 
    6.524859e-08, 6.533626e-08, 6.523825e-08, 6.519231e-08, 6.570255e-08, 
    6.541605e-08, 6.584592e-08, 6.582213e-08, 6.562759e-08, 6.582481e-08, 
    6.389985e-08, 6.384432e-08, 6.365153e-08, 6.38024e-08, 6.352751e-08, 
    6.368138e-08, 6.376987e-08, 6.411125e-08, 6.418625e-08, 6.425581e-08, 
    6.439316e-08, 6.456945e-08, 6.487869e-08, 6.514775e-08, 6.539337e-08, 
    6.537537e-08, 6.538171e-08, 6.543657e-08, 6.530066e-08, 6.545889e-08, 
    6.548544e-08, 6.541601e-08, 6.581894e-08, 6.570383e-08, 6.582162e-08, 
    6.574668e-08, 6.386237e-08, 6.395581e-08, 6.390532e-08, 6.400027e-08, 
    6.393338e-08, 6.42308e-08, 6.431998e-08, 6.473723e-08, 6.456598e-08, 
    6.483852e-08, 6.459366e-08, 6.463705e-08, 6.484741e-08, 6.460689e-08, 
    6.513292e-08, 6.47763e-08, 6.543871e-08, 6.50826e-08, 6.546102e-08, 
    6.53923e-08, 6.550608e-08, 6.560798e-08, 6.573618e-08, 6.597273e-08, 
    6.591795e-08, 6.611577e-08, 6.40951e-08, 6.42163e-08, 6.420562e-08, 
    6.433245e-08, 6.442625e-08, 6.462955e-08, 6.49556e-08, 6.483299e-08, 
    6.505808e-08, 6.510327e-08, 6.476129e-08, 6.497127e-08, 6.42974e-08, 
    6.440629e-08, 6.434146e-08, 6.410467e-08, 6.486125e-08, 6.447298e-08, 
    6.518994e-08, 6.49796e-08, 6.559345e-08, 6.528818e-08, 6.58878e-08, 
    6.614415e-08, 6.638538e-08, 6.666732e-08, 6.428244e-08, 6.420009e-08, 
    6.434753e-08, 6.455154e-08, 6.47408e-08, 6.499243e-08, 6.501818e-08, 
    6.506531e-08, 6.518741e-08, 6.529008e-08, 6.508023e-08, 6.531582e-08, 
    6.443155e-08, 6.489495e-08, 6.416896e-08, 6.438758e-08, 6.453951e-08, 
    6.447286e-08, 6.481897e-08, 6.490055e-08, 6.523204e-08, 6.506068e-08, 
    6.608088e-08, 6.562952e-08, 6.688197e-08, 6.653197e-08, 6.417132e-08, 
    6.428215e-08, 6.466789e-08, 6.448436e-08, 6.500922e-08, 6.513842e-08, 
    6.524344e-08, 6.53777e-08, 6.539219e-08, 6.547174e-08, 6.534139e-08, 
    6.546659e-08, 6.499297e-08, 6.520462e-08, 6.46238e-08, 6.476517e-08, 
    6.470013e-08, 6.46288e-08, 6.484896e-08, 6.508353e-08, 6.508854e-08, 
    6.516375e-08, 6.537572e-08, 6.501136e-08, 6.613915e-08, 6.544267e-08, 
    6.440301e-08, 6.461651e-08, 6.464699e-08, 6.456429e-08, 6.512547e-08, 
    6.492213e-08, 6.54698e-08, 6.532179e-08, 6.55643e-08, 6.544379e-08, 
    6.542606e-08, 6.527128e-08, 6.517492e-08, 6.493146e-08, 6.473337e-08, 
    6.457628e-08, 6.461281e-08, 6.478536e-08, 6.509788e-08, 6.539351e-08, 
    6.532875e-08, 6.554587e-08, 6.497117e-08, 6.521216e-08, 6.511902e-08, 
    6.536187e-08, 6.482973e-08, 6.52829e-08, 6.471389e-08, 6.476378e-08, 
    6.49181e-08, 6.522851e-08, 6.529717e-08, 6.53705e-08, 6.532525e-08, 
    6.510581e-08, 6.506986e-08, 6.491435e-08, 6.487141e-08, 6.475292e-08, 
    6.465483e-08, 6.474446e-08, 6.483858e-08, 6.51059e-08, 6.53468e-08, 
    6.560944e-08, 6.567371e-08, 6.59806e-08, 6.573079e-08, 6.614304e-08, 
    6.579257e-08, 6.639924e-08, 6.530915e-08, 6.578225e-08, 6.492512e-08, 
    6.501746e-08, 6.518448e-08, 6.556754e-08, 6.536073e-08, 6.560259e-08, 
    6.506844e-08, 6.479132e-08, 6.471961e-08, 6.458583e-08, 6.472267e-08, 
    6.471154e-08, 6.484247e-08, 6.48004e-08, 6.511478e-08, 6.494591e-08, 
    6.542562e-08, 6.560068e-08, 6.609504e-08, 6.63981e-08, 6.670659e-08, 
    6.684278e-08, 6.688423e-08, 6.690156e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.356978e-08, -6.384934e-08, -6.379499e-08, -6.402048e-08, -6.389539e-08, 
    -6.404304e-08, -6.362645e-08, -6.386044e-08, -6.371106e-08, 
    -6.359494e-08, -6.445807e-08, -6.403054e-08, -6.490213e-08, 
    -6.462948e-08, -6.531439e-08, -6.485971e-08, -6.540607e-08, 
    -6.530126e-08, -6.561668e-08, -6.552632e-08, -6.592977e-08, 
    -6.565838e-08, -6.61389e-08, -6.586495e-08, -6.590781e-08, -6.564943e-08, 
    -6.411657e-08, -6.440485e-08, -6.409949e-08, -6.41406e-08, -6.412215e-08, 
    -6.389798e-08, -6.378502e-08, -6.354841e-08, -6.359136e-08, 
    -6.376514e-08, -6.415908e-08, -6.402535e-08, -6.436237e-08, 
    -6.435476e-08, -6.472996e-08, -6.456079e-08, -6.51914e-08, -6.501217e-08, 
    -6.553009e-08, -6.539984e-08, -6.552398e-08, -6.548633e-08, 
    -6.552447e-08, -6.533344e-08, -6.541529e-08, -6.524719e-08, 
    -6.459248e-08, -6.478489e-08, -6.421101e-08, -6.386593e-08, 
    -6.363672e-08, -6.347406e-08, -6.349706e-08, -6.35409e-08, -6.376616e-08, 
    -6.397794e-08, -6.413933e-08, -6.42473e-08, -6.435366e-08, -6.467567e-08, 
    -6.484608e-08, -6.522765e-08, -6.515878e-08, -6.527544e-08, 
    -6.538689e-08, -6.557399e-08, -6.55432e-08, -6.562563e-08, -6.527236e-08, 
    -6.550714e-08, -6.511956e-08, -6.522556e-08, -6.438261e-08, 
    -6.406143e-08, -6.392494e-08, -6.380544e-08, -6.351474e-08, 
    -6.371549e-08, -6.363636e-08, -6.382462e-08, -6.394425e-08, 
    -6.388508e-08, -6.425024e-08, -6.410828e-08, -6.485618e-08, 
    -6.453404e-08, -6.537388e-08, -6.517291e-08, -6.542206e-08, 
    -6.529492e-08, -6.551276e-08, -6.53167e-08, -6.565631e-08, -6.573026e-08, 
    -6.567973e-08, -6.587384e-08, -6.530584e-08, -6.552398e-08, 
    -6.388343e-08, -6.389308e-08, -6.393803e-08, -6.374042e-08, 
    -6.372833e-08, -6.354723e-08, -6.370837e-08, -6.377699e-08, 
    -6.395118e-08, -6.405422e-08, -6.415217e-08, -6.436752e-08, 
    -6.460803e-08, -6.494434e-08, -6.518594e-08, -6.53479e-08, -6.524859e-08, 
    -6.533626e-08, -6.523825e-08, -6.519231e-08, -6.570255e-08, 
    -6.541605e-08, -6.584592e-08, -6.582213e-08, -6.562759e-08, 
    -6.582481e-08, -6.389985e-08, -6.384432e-08, -6.365153e-08, -6.38024e-08, 
    -6.352751e-08, -6.368138e-08, -6.376987e-08, -6.411125e-08, 
    -6.418625e-08, -6.425581e-08, -6.439316e-08, -6.456945e-08, 
    -6.487869e-08, -6.514775e-08, -6.539337e-08, -6.537537e-08, 
    -6.538171e-08, -6.543657e-08, -6.530066e-08, -6.545889e-08, 
    -6.548544e-08, -6.541601e-08, -6.581894e-08, -6.570383e-08, 
    -6.582162e-08, -6.574668e-08, -6.386237e-08, -6.395581e-08, 
    -6.390532e-08, -6.400027e-08, -6.393338e-08, -6.42308e-08, -6.431998e-08, 
    -6.473723e-08, -6.456598e-08, -6.483852e-08, -6.459366e-08, 
    -6.463705e-08, -6.484741e-08, -6.460689e-08, -6.513292e-08, -6.47763e-08, 
    -6.543871e-08, -6.50826e-08, -6.546102e-08, -6.53923e-08, -6.550608e-08, 
    -6.560798e-08, -6.573618e-08, -6.597273e-08, -6.591795e-08, 
    -6.611577e-08, -6.40951e-08, -6.42163e-08, -6.420562e-08, -6.433245e-08, 
    -6.442625e-08, -6.462955e-08, -6.49556e-08, -6.483299e-08, -6.505808e-08, 
    -6.510327e-08, -6.476129e-08, -6.497127e-08, -6.42974e-08, -6.440629e-08, 
    -6.434146e-08, -6.410467e-08, -6.486125e-08, -6.447298e-08, 
    -6.518994e-08, -6.49796e-08, -6.559345e-08, -6.528818e-08, -6.58878e-08, 
    -6.614415e-08, -6.638538e-08, -6.666732e-08, -6.428244e-08, 
    -6.420009e-08, -6.434753e-08, -6.455154e-08, -6.47408e-08, -6.499243e-08, 
    -6.501818e-08, -6.506531e-08, -6.518741e-08, -6.529008e-08, 
    -6.508023e-08, -6.531582e-08, -6.443155e-08, -6.489495e-08, 
    -6.416896e-08, -6.438758e-08, -6.453951e-08, -6.447286e-08, 
    -6.481897e-08, -6.490055e-08, -6.523204e-08, -6.506068e-08, 
    -6.608088e-08, -6.562952e-08, -6.688197e-08, -6.653197e-08, 
    -6.417132e-08, -6.428215e-08, -6.466789e-08, -6.448436e-08, 
    -6.500922e-08, -6.513842e-08, -6.524344e-08, -6.53777e-08, -6.539219e-08, 
    -6.547174e-08, -6.534139e-08, -6.546659e-08, -6.499297e-08, 
    -6.520462e-08, -6.46238e-08, -6.476517e-08, -6.470013e-08, -6.46288e-08, 
    -6.484896e-08, -6.508353e-08, -6.508854e-08, -6.516375e-08, 
    -6.537572e-08, -6.501136e-08, -6.613915e-08, -6.544267e-08, 
    -6.440301e-08, -6.461651e-08, -6.464699e-08, -6.456429e-08, 
    -6.512547e-08, -6.492213e-08, -6.54698e-08, -6.532179e-08, -6.55643e-08, 
    -6.544379e-08, -6.542606e-08, -6.527128e-08, -6.517492e-08, 
    -6.493146e-08, -6.473337e-08, -6.457628e-08, -6.461281e-08, 
    -6.478536e-08, -6.509788e-08, -6.539351e-08, -6.532875e-08, 
    -6.554587e-08, -6.497117e-08, -6.521216e-08, -6.511902e-08, 
    -6.536187e-08, -6.482973e-08, -6.52829e-08, -6.471389e-08, -6.476378e-08, 
    -6.49181e-08, -6.522851e-08, -6.529717e-08, -6.53705e-08, -6.532525e-08, 
    -6.510581e-08, -6.506986e-08, -6.491435e-08, -6.487141e-08, 
    -6.475292e-08, -6.465483e-08, -6.474446e-08, -6.483858e-08, -6.51059e-08, 
    -6.53468e-08, -6.560944e-08, -6.567371e-08, -6.59806e-08, -6.573079e-08, 
    -6.614304e-08, -6.579257e-08, -6.639924e-08, -6.530915e-08, 
    -6.578225e-08, -6.492512e-08, -6.501746e-08, -6.518448e-08, 
    -6.556754e-08, -6.536073e-08, -6.560259e-08, -6.506844e-08, 
    -6.479132e-08, -6.471961e-08, -6.458583e-08, -6.472267e-08, 
    -6.471154e-08, -6.484247e-08, -6.48004e-08, -6.511478e-08, -6.494591e-08, 
    -6.542562e-08, -6.560068e-08, -6.609504e-08, -6.63981e-08, -6.670659e-08, 
    -6.684278e-08, -6.688423e-08, -6.690156e-08 ;

 NET_NMIN =
  8.955569e-09, 8.994951e-09, 8.987294e-09, 9.019058e-09, 9.001438e-09, 
    9.022237e-09, 8.963553e-09, 8.996515e-09, 8.975472e-09, 8.959113e-09, 
    9.080702e-09, 9.020475e-09, 9.143255e-09, 9.104847e-09, 9.201329e-09, 
    9.137279e-09, 9.214243e-09, 9.199479e-09, 9.243911e-09, 9.231182e-09, 
    9.288014e-09, 9.249786e-09, 9.317473e-09, 9.278884e-09, 9.284921e-09, 
    9.248525e-09, 9.032595e-09, 9.073204e-09, 9.030189e-09, 9.03598e-09, 
    9.033381e-09, 9.001802e-09, 8.985889e-09, 8.952559e-09, 8.958609e-09, 
    8.98309e-09, 9.038583e-09, 9.019745e-09, 9.06722e-09, 9.066148e-09, 
    9.119002e-09, 9.095171e-09, 9.184004e-09, 9.158756e-09, 9.231713e-09, 
    9.213365e-09, 9.230852e-09, 9.225549e-09, 9.230921e-09, 9.204012e-09, 
    9.215541e-09, 9.191861e-09, 9.099635e-09, 9.12674e-09, 9.045897e-09, 
    8.997288e-09, 8.964999e-09, 8.942086e-09, 8.945325e-09, 8.951501e-09, 
    8.983233e-09, 9.013066e-09, 9.035801e-09, 9.05101e-09, 9.065994e-09, 
    9.111353e-09, 9.135358e-09, 9.189109e-09, 9.179408e-09, 9.195842e-09, 
    9.21154e-09, 9.237898e-09, 9.233559e-09, 9.245172e-09, 9.195407e-09, 
    9.228481e-09, 9.173883e-09, 9.188816e-09, 9.070072e-09, 9.024827e-09, 
    9.0056e-09, 8.988766e-09, 8.947816e-09, 8.976095e-09, 8.964948e-09, 
    8.991469e-09, 9.008321e-09, 8.999986e-09, 9.051425e-09, 9.031427e-09, 
    9.136781e-09, 9.091402e-09, 9.209709e-09, 9.181399e-09, 9.216494e-09, 
    9.198586e-09, 9.229272e-09, 9.201655e-09, 9.249494e-09, 9.25991e-09, 
    9.252791e-09, 9.280136e-09, 9.200124e-09, 9.230852e-09, 8.999752e-09, 
    9.001112e-09, 9.007445e-09, 8.979607e-09, 8.977905e-09, 8.952393e-09, 
    8.975093e-09, 8.98476e-09, 9.009297e-09, 9.023812e-09, 9.03761e-09, 
    9.067946e-09, 9.101826e-09, 9.149201e-09, 9.183235e-09, 9.206048e-09, 
    9.192059e-09, 9.20441e-09, 9.190603e-09, 9.184132e-09, 9.256008e-09, 
    9.215649e-09, 9.276203e-09, 9.272852e-09, 9.245448e-09, 9.273229e-09, 
    9.002067e-09, 8.994244e-09, 8.967085e-09, 8.988339e-09, 8.949614e-09, 
    8.971291e-09, 8.983755e-09, 9.031846e-09, 9.042411e-09, 9.052209e-09, 
    9.071559e-09, 9.096391e-09, 9.139953e-09, 9.177854e-09, 9.212453e-09, 
    9.209918e-09, 9.210811e-09, 9.218541e-09, 9.199394e-09, 9.221684e-09, 
    9.225425e-09, 9.215643e-09, 9.272403e-09, 9.256187e-09, 9.272781e-09, 
    9.262222e-09, 8.996786e-09, 9.009949e-09, 9.002837e-09, 9.016211e-09, 
    9.006789e-09, 9.048687e-09, 9.061249e-09, 9.120026e-09, 9.095903e-09, 
    9.134293e-09, 9.099802e-09, 9.105913e-09, 9.135547e-09, 9.101665e-09, 
    9.175766e-09, 9.12553e-09, 9.218841e-09, 9.168677e-09, 9.221984e-09, 
    9.212304e-09, 9.228331e-09, 9.242686e-09, 9.260744e-09, 9.294066e-09, 
    9.28635e-09, 9.314216e-09, 9.029571e-09, 9.046643e-09, 9.04514e-09, 
    9.063005e-09, 9.076219e-09, 9.104856e-09, 9.150787e-09, 9.133514e-09, 
    9.165222e-09, 9.171588e-09, 9.123416e-09, 9.152994e-09, 9.058069e-09, 
    9.073406e-09, 9.064274e-09, 9.030918e-09, 9.137496e-09, 9.082801e-09, 
    9.183797e-09, 9.154168e-09, 9.240639e-09, 9.197636e-09, 9.282102e-09, 
    9.318213e-09, 9.352194e-09, 9.391909e-09, 9.05596e-09, 9.04436e-09, 
    9.06513e-09, 9.093868e-09, 9.120529e-09, 9.155976e-09, 9.159601e-09, 
    9.166242e-09, 9.183442e-09, 9.197904e-09, 9.168343e-09, 9.201529e-09, 
    9.076965e-09, 9.142243e-09, 9.039975e-09, 9.070772e-09, 9.092173e-09, 
    9.082784e-09, 9.13154e-09, 9.143032e-09, 9.189728e-09, 9.165588e-09, 
    9.309301e-09, 9.245719e-09, 9.422147e-09, 9.372844e-09, 9.040307e-09, 
    9.05592e-09, 9.110259e-09, 9.084404e-09, 9.158341e-09, 9.17654e-09, 
    9.191334e-09, 9.210247e-09, 9.212288e-09, 9.223493e-09, 9.205132e-09, 
    9.222767e-09, 9.156051e-09, 9.185865e-09, 9.104047e-09, 9.123962e-09, 
    9.1148e-09, 9.104751e-09, 9.135765e-09, 9.168808e-09, 9.169513e-09, 
    9.180108e-09, 9.209967e-09, 9.158641e-09, 9.317509e-09, 9.219399e-09, 
    9.072945e-09, 9.10302e-09, 9.107313e-09, 9.095664e-09, 9.174716e-09, 
    9.146073e-09, 9.22322e-09, 9.20237e-09, 9.236532e-09, 9.219557e-09, 
    9.217059e-09, 9.195255e-09, 9.181681e-09, 9.147387e-09, 9.119482e-09, 
    9.097353e-09, 9.102498e-09, 9.126806e-09, 9.170829e-09, 9.212473e-09, 
    9.203351e-09, 9.233936e-09, 9.15298e-09, 9.186927e-09, 9.173807e-09, 
    9.208017e-09, 9.133056e-09, 9.196893e-09, 9.116738e-09, 9.123767e-09, 
    9.145504e-09, 9.189231e-09, 9.198903e-09, 9.209232e-09, 9.202858e-09, 
    9.171946e-09, 9.166881e-09, 9.144975e-09, 9.138928e-09, 9.122236e-09, 
    9.108417e-09, 9.121043e-09, 9.134303e-09, 9.171959e-09, 9.205893e-09, 
    9.242891e-09, 9.251944e-09, 9.295174e-09, 9.259985e-09, 9.318057e-09, 
    9.268687e-09, 9.354146e-09, 9.200591e-09, 9.267233e-09, 9.146493e-09, 
    9.159501e-09, 9.183029e-09, 9.236989e-09, 9.207856e-09, 9.241926e-09, 
    9.166683e-09, 9.127645e-09, 9.117544e-09, 9.098699e-09, 9.117975e-09, 
    9.116407e-09, 9.134851e-09, 9.128924e-09, 9.173209e-09, 9.149421e-09, 
    9.216997e-09, 9.241656e-09, 9.311296e-09, 9.353987e-09, 9.397441e-09, 
    9.416627e-09, 9.422465e-09, 9.424906e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.484872e-14, 4.497019e-14, 4.49466e-14, 4.504447e-14, 4.49902e-14, 
    4.505427e-14, 4.487338e-14, 4.497499e-14, 4.491014e-14, 4.485969e-14, 
    4.523413e-14, 4.504884e-14, 4.542646e-14, 4.530849e-14, 4.560464e-14, 
    4.540809e-14, 4.564424e-14, 4.559901e-14, 4.573518e-14, 4.569619e-14, 
    4.587009e-14, 4.575318e-14, 4.59602e-14, 4.584221e-14, 4.586065e-14, 
    4.574931e-14, 4.508619e-14, 4.521107e-14, 4.507878e-14, 4.50966e-14, 
    4.508862e-14, 4.499131e-14, 4.494222e-14, 4.483946e-14, 4.485813e-14, 
    4.493362e-14, 4.510461e-14, 4.504662e-14, 4.51928e-14, 4.51895e-14, 
    4.5352e-14, 4.527876e-14, 4.555155e-14, 4.547411e-14, 4.569782e-14, 
    4.564159e-14, 4.569517e-14, 4.567893e-14, 4.569538e-14, 4.56129e-14, 
    4.564825e-14, 4.557566e-14, 4.529247e-14, 4.537577e-14, 4.512715e-14, 
    4.497733e-14, 4.487783e-14, 4.480714e-14, 4.481714e-14, 4.483618e-14, 
    4.493406e-14, 4.502604e-14, 4.509608e-14, 4.514291e-14, 4.518903e-14, 
    4.532841e-14, 4.540221e-14, 4.556718e-14, 4.553746e-14, 4.558784e-14, 
    4.563599e-14, 4.571675e-14, 4.570347e-14, 4.573903e-14, 4.558653e-14, 
    4.568789e-14, 4.552054e-14, 4.556632e-14, 4.520142e-14, 4.506227e-14, 
    4.500296e-14, 4.495113e-14, 4.482482e-14, 4.491205e-14, 4.487767e-14, 
    4.495948e-14, 4.501142e-14, 4.498574e-14, 4.514419e-14, 4.508261e-14, 
    4.540658e-14, 4.526715e-14, 4.563038e-14, 4.554357e-14, 4.565118e-14, 
    4.559629e-14, 4.569032e-14, 4.560569e-14, 4.575227e-14, 4.578414e-14, 
    4.576236e-14, 4.584606e-14, 4.5601e-14, 4.569516e-14, 4.498502e-14, 
    4.49892e-14, 4.500873e-14, 4.492288e-14, 4.491763e-14, 4.483895e-14, 
    4.490898e-14, 4.493877e-14, 4.501444e-14, 4.505915e-14, 4.510164e-14, 
    4.519502e-14, 4.529919e-14, 4.544474e-14, 4.554919e-14, 4.561917e-14, 
    4.557627e-14, 4.561414e-14, 4.55718e-14, 4.555196e-14, 4.577219e-14, 
    4.564857e-14, 4.583403e-14, 4.582378e-14, 4.573986e-14, 4.582493e-14, 
    4.499214e-14, 4.496804e-14, 4.488427e-14, 4.494983e-14, 4.483037e-14, 
    4.489724e-14, 4.493566e-14, 4.508386e-14, 4.511643e-14, 4.514659e-14, 
    4.520614e-14, 4.528251e-14, 4.541635e-14, 4.553267e-14, 4.56388e-14, 
    4.563103e-14, 4.563376e-14, 4.565745e-14, 4.559876e-14, 4.566708e-14, 
    4.567853e-14, 4.564857e-14, 4.582241e-14, 4.577277e-14, 4.582356e-14, 
    4.579125e-14, 4.497588e-14, 4.501644e-14, 4.499452e-14, 4.503573e-14, 
    4.500669e-14, 4.513571e-14, 4.517436e-14, 4.535511e-14, 4.5281e-14, 
    4.539896e-14, 4.5293e-14, 4.531177e-14, 4.540274e-14, 4.529874e-14, 
    4.552626e-14, 4.5372e-14, 4.565837e-14, 4.550447e-14, 4.5668e-14, 
    4.563834e-14, 4.568746e-14, 4.573142e-14, 4.578672e-14, 4.588865e-14, 
    4.586506e-14, 4.595027e-14, 4.507689e-14, 4.512944e-14, 4.512484e-14, 
    4.517983e-14, 4.522047e-14, 4.530854e-14, 4.544963e-14, 4.53966e-14, 
    4.549396e-14, 4.551349e-14, 4.536558e-14, 4.545639e-14, 4.516461e-14, 
    4.521178e-14, 4.518372e-14, 4.508102e-14, 4.540879e-14, 4.524068e-14, 
    4.555091e-14, 4.546002e-14, 4.572515e-14, 4.559333e-14, 4.585207e-14, 
    4.596242e-14, 4.60663e-14, 4.618743e-14, 4.515814e-14, 4.512244e-14, 
    4.518637e-14, 4.527471e-14, 4.53567e-14, 4.546556e-14, 4.547671e-14, 
    4.549708e-14, 4.554984e-14, 4.559419e-14, 4.550349e-14, 4.560531e-14, 
    4.522266e-14, 4.542338e-14, 4.510892e-14, 4.520366e-14, 4.526952e-14, 
    4.524066e-14, 4.539055e-14, 4.542584e-14, 4.556909e-14, 4.549509e-14, 
    4.593517e-14, 4.574066e-14, 4.627966e-14, 4.612929e-14, 4.510996e-14, 
    4.515802e-14, 4.532512e-14, 4.524565e-14, 4.547284e-14, 4.552868e-14, 
    4.557405e-14, 4.563201e-14, 4.563829e-14, 4.567262e-14, 4.561636e-14, 
    4.567041e-14, 4.546579e-14, 4.555727e-14, 4.530606e-14, 4.536724e-14, 
    4.533911e-14, 4.530823e-14, 4.540352e-14, 4.550492e-14, 4.550713e-14, 
    4.553958e-14, 4.5631e-14, 4.547376e-14, 4.596017e-14, 4.565993e-14, 
    4.521041e-14, 4.530284e-14, 4.531609e-14, 4.528029e-14, 4.552308e-14, 
    4.543516e-14, 4.567179e-14, 4.560789e-14, 4.571258e-14, 4.566056e-14, 
    4.565291e-14, 4.558607e-14, 4.554443e-14, 4.543919e-14, 4.535347e-14, 
    4.528549e-14, 4.53013e-14, 4.537598e-14, 4.551112e-14, 4.563884e-14, 
    4.561086e-14, 4.570463e-14, 4.545638e-14, 4.55605e-14, 4.552027e-14, 
    4.562519e-14, 4.539518e-14, 4.559095e-14, 4.534507e-14, 4.536666e-14, 
    4.543342e-14, 4.556753e-14, 4.559726e-14, 4.56289e-14, 4.560939e-14, 
    4.551456e-14, 4.549904e-14, 4.54318e-14, 4.541321e-14, 4.536197e-14, 
    4.53195e-14, 4.535829e-14, 4.5399e-14, 4.551462e-14, 4.561866e-14, 
    4.573204e-14, 4.575978e-14, 4.589195e-14, 4.578431e-14, 4.596183e-14, 
    4.581083e-14, 4.607213e-14, 4.560234e-14, 4.580648e-14, 4.543647e-14, 
    4.54764e-14, 4.554852e-14, 4.571391e-14, 4.56247e-14, 4.572905e-14, 
    4.549843e-14, 4.537853e-14, 4.534754e-14, 4.528962e-14, 4.534887e-14, 
    4.534405e-14, 4.540072e-14, 4.538251e-14, 4.551846e-14, 4.544546e-14, 
    4.56527e-14, 4.572824e-14, 4.594133e-14, 4.607172e-14, 4.620437e-14, 
    4.626286e-14, 4.628066e-14, 4.628809e-14 ;

 POT_F_DENIT =
  1.021877e-12, 1.024722e-12, 1.024168e-12, 1.026462e-12, 1.025188e-12, 
    1.02669e-12, 1.022451e-12, 1.024832e-12, 1.023311e-12, 1.022128e-12, 
    1.03091e-12, 1.02656e-12, 1.03542e-12, 1.032648e-12, 1.039606e-12, 
    1.034989e-12, 1.040536e-12, 1.03947e-12, 1.042671e-12, 1.041753e-12, 
    1.045848e-12, 1.043093e-12, 1.047967e-12, 1.045189e-12, 1.045623e-12, 
    1.043e-12, 1.027438e-12, 1.030373e-12, 1.027264e-12, 1.027682e-12, 
    1.027493e-12, 1.025213e-12, 1.024064e-12, 1.021654e-12, 1.022091e-12, 
    1.02386e-12, 1.027867e-12, 1.026505e-12, 1.029931e-12, 1.029854e-12, 
    1.033667e-12, 1.031948e-12, 1.038354e-12, 1.036532e-12, 1.041791e-12, 
    1.040468e-12, 1.041728e-12, 1.041345e-12, 1.041731e-12, 1.039793e-12, 
    1.040622e-12, 1.038916e-12, 1.032276e-12, 1.034231e-12, 1.028397e-12, 
    1.024888e-12, 1.022553e-12, 1.020898e-12, 1.021131e-12, 1.021577e-12, 
    1.023869e-12, 1.026022e-12, 1.027663e-12, 1.028761e-12, 1.029841e-12, 
    1.033117e-12, 1.034847e-12, 1.038721e-12, 1.038021e-12, 1.039206e-12, 
    1.040336e-12, 1.042235e-12, 1.041922e-12, 1.042758e-12, 1.039171e-12, 
    1.041555e-12, 1.037618e-12, 1.038695e-12, 1.030145e-12, 1.026874e-12, 
    1.025487e-12, 1.02427e-12, 1.02131e-12, 1.023354e-12, 1.022548e-12, 
    1.024462e-12, 1.025679e-12, 1.025076e-12, 1.02879e-12, 1.027346e-12, 
    1.034949e-12, 1.031675e-12, 1.040205e-12, 1.038163e-12, 1.040692e-12, 
    1.039402e-12, 1.041612e-12, 1.039622e-12, 1.043068e-12, 1.043819e-12, 
    1.043305e-12, 1.045274e-12, 1.039508e-12, 1.041723e-12, 1.025063e-12, 
    1.025161e-12, 1.025617e-12, 1.023607e-12, 1.023483e-12, 1.021639e-12, 
    1.023278e-12, 1.023977e-12, 1.025748e-12, 1.026796e-12, 1.027791e-12, 
    1.029981e-12, 1.032426e-12, 1.035842e-12, 1.038295e-12, 1.039939e-12, 
    1.03893e-12, 1.039819e-12, 1.038824e-12, 1.038357e-12, 1.043536e-12, 
    1.040629e-12, 1.044989e-12, 1.044748e-12, 1.042774e-12, 1.044774e-12, 
    1.025229e-12, 1.024663e-12, 1.022701e-12, 1.024235e-12, 1.021437e-12, 
    1.023004e-12, 1.023904e-12, 1.027376e-12, 1.028137e-12, 1.028845e-12, 
    1.03024e-12, 1.032032e-12, 1.035175e-12, 1.037907e-12, 1.0404e-12, 
    1.040216e-12, 1.04028e-12, 1.040837e-12, 1.039457e-12, 1.041062e-12, 
    1.041331e-12, 1.040626e-12, 1.044714e-12, 1.043546e-12, 1.044741e-12, 
    1.043979e-12, 1.024846e-12, 1.025796e-12, 1.025281e-12, 1.026248e-12, 
    1.025566e-12, 1.028592e-12, 1.029498e-12, 1.033739e-12, 1.031997e-12, 
    1.034767e-12, 1.032277e-12, 1.032718e-12, 1.034857e-12, 1.03241e-12, 
    1.037755e-12, 1.034132e-12, 1.040858e-12, 1.037243e-12, 1.041083e-12, 
    1.040385e-12, 1.041539e-12, 1.042574e-12, 1.043873e-12, 1.046274e-12, 
    1.045716e-12, 1.047723e-12, 1.027212e-12, 1.028444e-12, 1.028335e-12, 
    1.029624e-12, 1.030577e-12, 1.032643e-12, 1.035956e-12, 1.034709e-12, 
    1.036995e-12, 1.037454e-12, 1.033979e-12, 1.036113e-12, 1.029264e-12, 
    1.030371e-12, 1.02971e-12, 1.027302e-12, 1.034993e-12, 1.031046e-12, 
    1.03833e-12, 1.036193e-12, 1.042425e-12, 1.039327e-12, 1.04541e-12, 
    1.048012e-12, 1.050455e-12, 1.053312e-12, 1.029116e-12, 1.028277e-12, 
    1.029776e-12, 1.031851e-12, 1.033773e-12, 1.036329e-12, 1.03659e-12, 
    1.037068e-12, 1.038307e-12, 1.03935e-12, 1.037219e-12, 1.039609e-12, 
    1.030628e-12, 1.035335e-12, 1.027955e-12, 1.030179e-12, 1.031721e-12, 
    1.031043e-12, 1.03456e-12, 1.035388e-12, 1.038755e-12, 1.037014e-12, 
    1.047369e-12, 1.04279e-12, 1.055484e-12, 1.05194e-12, 1.027984e-12, 
    1.02911e-12, 1.033032e-12, 1.031166e-12, 1.036498e-12, 1.037811e-12, 
    1.038875e-12, 1.040239e-12, 1.040385e-12, 1.041193e-12, 1.039868e-12, 
    1.041139e-12, 1.036329e-12, 1.038479e-12, 1.032577e-12, 1.034013e-12, 
    1.033352e-12, 1.032626e-12, 1.034863e-12, 1.037247e-12, 1.037296e-12, 
    1.03806e-12, 1.040215e-12, 1.03651e-12, 1.04796e-12, 1.040893e-12, 
    1.030339e-12, 1.032509e-12, 1.032817e-12, 1.031977e-12, 1.037678e-12, 
    1.035612e-12, 1.041173e-12, 1.039669e-12, 1.04213e-12, 1.040907e-12, 
    1.040726e-12, 1.039155e-12, 1.038176e-12, 1.035703e-12, 1.033689e-12, 
    1.032092e-12, 1.032463e-12, 1.034217e-12, 1.037391e-12, 1.040392e-12, 
    1.039735e-12, 1.041937e-12, 1.036101e-12, 1.038549e-12, 1.037602e-12, 
    1.040068e-12, 1.034674e-12, 1.039281e-12, 1.033496e-12, 1.034002e-12, 
    1.03557e-12, 1.038724e-12, 1.039418e-12, 1.040164e-12, 1.039702e-12, 
    1.037475e-12, 1.037109e-12, 1.035528e-12, 1.035092e-12, 1.033887e-12, 
    1.032889e-12, 1.0338e-12, 1.034756e-12, 1.037471e-12, 1.039917e-12, 
    1.042582e-12, 1.043234e-12, 1.046349e-12, 1.043814e-12, 1.047997e-12, 
    1.044443e-12, 1.050592e-12, 1.039544e-12, 1.044346e-12, 1.035641e-12, 
    1.036578e-12, 1.038275e-12, 1.042164e-12, 1.040062e-12, 1.042519e-12, 
    1.037094e-12, 1.034279e-12, 1.033548e-12, 1.032189e-12, 1.033578e-12, 
    1.033465e-12, 1.034795e-12, 1.034367e-12, 1.03756e-12, 1.035845e-12, 
    1.040715e-12, 1.042493e-12, 1.047507e-12, 1.050579e-12, 1.053703e-12, 
    1.055082e-12, 1.055501e-12, 1.055676e-12 ;

 POT_F_NIT =
  4.013708e-11, 4.04835e-11, 4.041602e-11, 4.069631e-11, 4.05407e-11, 
    4.07244e-11, 4.020716e-11, 4.049725e-11, 4.031193e-11, 4.016816e-11, 
    4.124308e-11, 4.07088e-11, 4.180183e-11, 4.145828e-11, 4.232403e-11, 
    4.174826e-11, 4.244061e-11, 4.230734e-11, 4.270907e-11, 4.259377e-11, 
    4.310976e-11, 4.276232e-11, 4.337848e-11, 4.302664e-11, 4.308158e-11, 
    4.275086e-11, 4.081606e-11, 4.11764e-11, 4.079475e-11, 4.084602e-11, 
    4.0823e-11, 4.054389e-11, 4.040362e-11, 4.011063e-11, 4.016373e-11, 
    4.037896e-11, 4.086906e-11, 4.070233e-11, 4.112315e-11, 4.111363e-11, 
    4.15847e-11, 4.137196e-11, 4.216787e-11, 4.194085e-11, 4.259857e-11, 
    4.243266e-11, 4.259077e-11, 4.254279e-11, 4.259138e-11, 4.234819e-11, 
    4.245229e-11, 4.223862e-11, 4.141181e-11, 4.165395e-11, 4.09339e-11, 
    4.050408e-11, 4.021985e-11, 4.00188e-11, 4.004718e-11, 4.010134e-11, 
    4.038021e-11, 4.06433e-11, 4.08444e-11, 4.09792e-11, 4.111224e-11, 
    4.151636e-11, 4.173105e-11, 4.221384e-11, 4.212649e-11, 4.227451e-11, 
    4.241617e-11, 4.265455e-11, 4.261526e-11, 4.272046e-11, 4.227058e-11, 
    4.25693e-11, 4.207674e-11, 4.221117e-11, 4.114853e-11, 4.074729e-11, 
    4.057739e-11, 4.042895e-11, 4.006902e-11, 4.03174e-11, 4.021939e-11, 
    4.045275e-11, 4.060139e-11, 4.052783e-11, 4.098288e-11, 4.080565e-11, 
    4.174378e-11, 4.133835e-11, 4.239964e-11, 4.21444e-11, 4.246092e-11, 
    4.229925e-11, 4.257645e-11, 4.232692e-11, 4.275963e-11, 4.285416e-11, 
    4.278954e-11, 4.3038e-11, 4.231309e-11, 4.259073e-11, 4.052579e-11, 
    4.053779e-11, 4.059367e-11, 4.034829e-11, 4.03333e-11, 4.010915e-11, 
    4.030856e-11, 4.039363e-11, 4.061e-11, 4.073827e-11, 4.086039e-11, 
    4.112958e-11, 4.143129e-11, 4.185508e-11, 4.216092e-11, 4.236657e-11, 
    4.22404e-11, 4.235177e-11, 4.222727e-11, 4.216897e-11, 4.281872e-11, 
    4.245325e-11, 4.30022e-11, 4.297173e-11, 4.272293e-11, 4.297515e-11, 
    4.05462e-11, 4.04772e-11, 4.023816e-11, 4.042516e-11, 4.008477e-11, 
    4.027512e-11, 4.038479e-11, 4.080936e-11, 4.090293e-11, 4.098982e-11, 
    4.116169e-11, 4.13828e-11, 4.177218e-11, 4.211249e-11, 4.24244e-11, 
    4.24015e-11, 4.240956e-11, 4.247938e-11, 4.230651e-11, 4.250779e-11, 
    4.254161e-11, 4.245319e-11, 4.296764e-11, 4.282033e-11, 4.297107e-11, 
    4.287511e-11, 4.049962e-11, 4.061576e-11, 4.055297e-11, 4.067108e-11, 
    4.058785e-11, 4.095858e-11, 4.107007e-11, 4.159383e-11, 4.137844e-11, 
    4.172148e-11, 4.141321e-11, 4.146775e-11, 4.17327e-11, 4.142982e-11, 
    4.209368e-11, 4.164302e-11, 4.248209e-11, 4.202992e-11, 4.25105e-11, 
    4.242301e-11, 4.25679e-11, 4.269789e-11, 4.286169e-11, 4.316482e-11, 
    4.309452e-11, 4.334865e-11, 4.078923e-11, 4.094046e-11, 4.092713e-11, 
    4.108568e-11, 4.120313e-11, 4.145832e-11, 4.186931e-11, 4.17145e-11, 
    4.19989e-11, 4.205612e-11, 4.162412e-11, 4.188909e-11, 4.104179e-11, 
    4.117808e-11, 4.10969e-11, 4.080108e-11, 4.175012e-11, 4.126166e-11, 
    4.216593e-11, 4.189959e-11, 4.267933e-11, 4.229062e-11, 4.305585e-11, 
    4.338517e-11, 4.369625e-11, 4.406129e-11, 4.102312e-11, 4.09202e-11, 
    4.110454e-11, 4.136031e-11, 4.159832e-11, 4.191586e-11, 4.194841e-11, 
    4.200806e-11, 4.216276e-11, 4.229308e-11, 4.202692e-11, 4.232576e-11, 
    4.120973e-11, 4.179266e-11, 4.088128e-11, 4.115464e-11, 4.134515e-11, 
    4.126151e-11, 4.169677e-11, 4.17997e-11, 4.221933e-11, 4.200213e-11, 
    4.330376e-11, 4.272535e-11, 4.434026e-11, 4.388584e-11, 4.088428e-11, 
    4.102274e-11, 4.150654e-11, 4.127598e-11, 4.193709e-11, 4.210066e-11, 
    4.223385e-11, 4.240445e-11, 4.242288e-11, 4.252415e-11, 4.235826e-11, 
    4.251758e-11, 4.191649e-11, 4.218455e-11, 4.145104e-11, 4.162896e-11, 
    4.154705e-11, 4.145731e-11, 4.173459e-11, 4.203106e-11, 4.203739e-11, 
    4.213269e-11, 4.240186e-11, 4.19397e-11, 4.337871e-11, 4.248706e-11, 
    4.1174e-11, 4.144191e-11, 4.148023e-11, 4.13763e-11, 4.208423e-11, 
    4.1827e-11, 4.252168e-11, 4.233334e-11, 4.264214e-11, 4.248855e-11, 
    4.246596e-11, 4.226916e-11, 4.214687e-11, 4.183875e-11, 4.158889e-11, 
    4.139131e-11, 4.14372e-11, 4.165439e-11, 4.204922e-11, 4.24245e-11, 
    4.234214e-11, 4.261858e-11, 4.188888e-11, 4.219407e-11, 4.207597e-11, 
    4.238424e-11, 4.171038e-11, 4.228396e-11, 4.156442e-11, 4.162724e-11, 
    4.182189e-11, 4.221488e-11, 4.230205e-11, 4.239527e-11, 4.233773e-11, 
    4.20593e-11, 4.201376e-11, 4.181713e-11, 4.176292e-11, 4.161351e-11, 
    4.149003e-11, 4.160284e-11, 4.172148e-11, 4.205938e-11, 4.236508e-11, 
    4.269969e-11, 4.278177e-11, 4.317487e-11, 4.285474e-11, 4.338369e-11, 
    4.293379e-11, 4.37141e-11, 4.23173e-11, 4.292066e-11, 4.183076e-11, 
    4.194747e-11, 4.215902e-11, 4.264626e-11, 4.238284e-11, 4.269099e-11, 
    4.201197e-11, 4.166191e-11, 4.157156e-11, 4.140331e-11, 4.15754e-11, 
    4.156139e-11, 4.172639e-11, 4.167332e-11, 4.20706e-11, 4.185696e-11, 
    4.246534e-11, 4.26885e-11, 4.332194e-11, 4.371265e-11, 4.411221e-11, 
    4.428921e-11, 4.434316e-11, 4.436572e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001208392, 0.00120832, 0.001208334, 0.001208277, 0.001208308, 
    0.001208271, 0.001208376, 0.001208318, 0.001208355, 0.001208384, 
    0.001208168, 0.001208274, 0.001208053, 0.001208121, 0.001207947, 
    0.001208064, 0.001207923, 0.001207949, 0.001207868, 0.001207891, 
    0.001207791, 0.001207858, 0.001207737, 0.001207807, 0.001207796, 
    0.00120786, 0.001208252, 0.001208182, 0.001208256, 0.001208246, 
    0.00120825, 0.001208308, 0.001208338, 0.001208396, 0.001208385, 
    0.001208342, 0.001208241, 0.001208275, 0.001208188, 0.00120819, 
    0.001208096, 0.001208138, 0.001207977, 0.001208024, 0.00120789, 
    0.001207924, 0.001207892, 0.001207902, 0.001207892, 0.001207941, 
    0.00120792, 0.001207962, 0.001208131, 0.001208082, 0.001208228, 
    0.001208318, 0.001208374, 0.001208415, 0.001208409, 0.001208399, 
    0.001208341, 0.001208287, 0.001208245, 0.001208218, 0.001208191, 
    0.001208112, 0.001208067, 0.001207968, 0.001207985, 0.001207956, 
    0.001207927, 0.00120788, 0.001207887, 0.001207867, 0.001207956, 
    0.001207897, 0.001207996, 0.001207968, 0.001208188, 0.001208265, 
    0.001208302, 0.001208331, 0.001208405, 0.001208354, 0.001208374, 
    0.001208326, 0.001208295, 0.00120831, 0.001208217, 0.001208253, 
    0.001208065, 0.001208146, 0.00120793, 0.001207981, 0.001207918, 
    0.00120795, 0.001207895, 0.001207944, 0.001207859, 0.001207841, 
    0.001207853, 0.001207803, 0.001207947, 0.001207893, 0.001208311, 
    0.001208308, 0.001208297, 0.001208348, 0.001208351, 0.001208397, 
    0.001208356, 0.001208338, 0.001208293, 0.001208267, 0.001208242, 
    0.001208188, 0.001208127, 0.001208042, 0.001207978, 0.001207937, 
    0.001207962, 0.001207939, 0.001207964, 0.001207976, 0.001207848, 
    0.00120792, 0.001207811, 0.001207816, 0.001207866, 0.001207816, 
    0.001208307, 0.00120832, 0.00120837, 0.001208331, 0.001208402, 
    0.001208363, 0.001208341, 0.001208254, 0.001208233, 0.001208216, 
    0.001208181, 0.001208136, 0.001208058, 0.001207988, 0.001207925, 
    0.001207929, 0.001207928, 0.001207914, 0.001207949, 0.001207909, 
    0.001207902, 0.001207919, 0.001207817, 0.001207846, 0.001207817, 
    0.001207835, 0.001208316, 0.001208292, 0.001208305, 0.001208281, 
    0.001208298, 0.001208224, 0.001208201, 0.001208095, 0.001208137, 
    0.001208069, 0.00120813, 0.001208119, 0.001208068, 0.001208126, 
    0.001207994, 0.001208086, 0.001207914, 0.001208008, 0.001207908, 
    0.001207925, 0.001207896, 0.001207871, 0.001207838, 0.001207779, 
    0.001207793, 0.001207743, 0.001208257, 0.001208227, 0.001208228, 
    0.001208196, 0.001208173, 0.001208121, 0.001208038, 0.001208069, 
    0.001208012, 0.001208001, 0.001208087, 0.001208035, 0.001208206, 
    0.001208179, 0.001208194, 0.001208255, 0.001208063, 0.001208162, 
    0.001207977, 0.001208032, 0.001207875, 0.001207953, 0.0012078, 
    0.001207737, 0.001207674, 0.001207605, 0.001208209, 0.00120823, 
    0.001208192, 0.001208142, 0.001208093, 0.001208029, 0.001208022, 
    0.00120801, 0.001207977, 0.001207951, 0.001208007, 0.001207945, 
    0.001208175, 0.001208054, 0.001208238, 0.001208184, 0.001208144, 
    0.001208161, 0.001208072, 0.001208052, 0.001207967, 0.001208011, 
    0.001207754, 0.001207867, 0.00120755, 0.001207639, 0.001208237, 
    0.001208209, 0.001208112, 0.001208158, 0.001208024, 0.001207992, 
    0.001207963, 0.00120793, 0.001207925, 0.001207906, 0.001207938, 
    0.001207907, 0.001208029, 0.001207973, 0.001208122, 0.001208087, 
    0.001208103, 0.001208121, 0.001208065, 0.001208007, 0.001208004, 
    0.001207984, 0.001207935, 0.001208024, 0.001207742, 0.001207917, 
    0.001208178, 0.001208126, 0.001208117, 0.001208137, 0.001207995, 
    0.001208047, 0.001207906, 0.001207943, 0.001207882, 0.001207912, 
    0.001207917, 0.001207956, 0.001207981, 0.001208045, 0.001208095, 
    0.001208134, 0.001208125, 0.001208082, 0.001208003, 0.001207926, 
    0.001207942, 0.001207886, 0.001208034, 0.001207972, 0.001207997, 
    0.001207933, 0.00120807, 0.001207958, 0.001208099, 0.001208086, 
    0.001208048, 0.001207969, 0.001207949, 0.001207931, 0.001207942, 
    0.001208001, 0.001208009, 0.001208048, 0.00120806, 0.001208089, 
    0.001208114, 0.001208092, 0.001208068, 0.001208, 0.001207938, 
    0.001207871, 0.001207854, 0.00120778, 0.001207842, 0.001207741, 
    0.00120783, 0.001207675, 0.001207949, 0.00120783, 0.001208045, 
    0.001208022, 0.00120798, 0.001207883, 0.001207934, 0.001207874, 
    0.001208009, 0.001208081, 0.001208098, 0.001208132, 0.001208097, 
    0.0012081, 0.001208066, 0.001208077, 0.001207998, 0.00120804, 
    0.001207917, 0.001207874, 0.001207748, 0.001207673, 0.001207593, 
    0.001207559, 0.001207548, 0.001207544 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  -1.484414e-07, -1.486925e-07, -1.486433e-07, -1.488465e-07, -1.487332e-07, 
    -1.488666e-07, -1.484916e-07, -1.487031e-07, -1.485677e-07, 
    -1.484631e-07, -1.49241e-07, -1.488553e-07, -1.496338e-07, -1.493898e-07, 
    -1.500032e-07, -1.495968e-07, -1.50084e-07, -1.4999e-07, -1.502689e-07, 
    -1.501889e-07, -1.505482e-07, -1.503057e-07, -1.507315e-07, 
    -1.504895e-07, -1.50528e-07, -1.50298e-07, -1.489315e-07, -1.491936e-07, 
    -1.489164e-07, -1.489537e-07, -1.489366e-07, -1.487361e-07, 
    -1.486359e-07, -1.484211e-07, -1.484599e-07, -1.48617e-07, -1.489704e-07, 
    -1.488497e-07, -1.491507e-07, -1.491439e-07, -1.494792e-07, 
    -1.493282e-07, -1.498926e-07, -1.497297e-07, -1.501922e-07, 
    -1.500771e-07, -1.501871e-07, -1.501536e-07, -1.501875e-07, 
    -1.500186e-07, -1.500911e-07, -1.499418e-07, -1.493568e-07, 
    -1.495285e-07, -1.490164e-07, -1.487095e-07, -1.485012e-07, 
    -1.483544e-07, -1.483752e-07, -1.484151e-07, -1.48618e-07, -1.488072e-07, 
    -1.489514e-07, -1.49048e-07, -1.491429e-07, -1.494337e-07, -1.495839e-07, 
    -1.499256e-07, -1.498633e-07, -1.499678e-07, -1.500656e-07, 
    -1.502315e-07, -1.50204e-07, -1.502774e-07, -1.49964e-07, -1.501729e-07, 
    -1.498247e-07, -1.499226e-07, -1.49174e-07, -1.48882e-07, -1.487621e-07, 
    -1.48653e-07, -1.483912e-07, -1.485723e-07, -1.485011e-07, -1.486694e-07, 
    -1.48777e-07, -1.487236e-07, -1.490507e-07, -1.489239e-07, -1.495929e-07, 
    -1.493051e-07, -1.500542e-07, -1.498759e-07, -1.500967e-07, 
    -1.499838e-07, -1.501776e-07, -1.500032e-07, -1.503043e-07, 
    -1.503703e-07, -1.503253e-07, -1.504964e-07, -1.499937e-07, 
    -1.501876e-07, -1.487223e-07, -1.487311e-07, -1.487712e-07, 
    -1.485948e-07, -1.485838e-07, -1.484203e-07, -1.485653e-07, 
    -1.486274e-07, -1.487828e-07, -1.488756e-07, -1.489633e-07, 
    -1.491559e-07, -1.493713e-07, -1.496706e-07, -1.498876e-07, 
    -1.500308e-07, -1.499427e-07, -1.500206e-07, -1.499337e-07, 
    -1.498927e-07, -1.503459e-07, -1.500921e-07, -1.504718e-07, 
    -1.504506e-07, -1.502793e-07, -1.50453e-07, -1.487371e-07, -1.48687e-07, 
    -1.485143e-07, -1.486494e-07, -1.484024e-07, -1.485414e-07, 
    -1.486217e-07, -1.489277e-07, -1.489935e-07, -1.490561e-07, 
    -1.491785e-07, -1.493359e-07, -1.49612e-07, -1.498542e-07, -1.500711e-07, 
    -1.500551e-07, -1.500608e-07, -1.501097e-07, -1.499892e-07, 
    -1.501295e-07, -1.501535e-07, -1.500914e-07, -1.504478e-07, 
    -1.503461e-07, -1.504502e-07, -1.503838e-07, -1.487031e-07, 
    -1.487873e-07, -1.487419e-07, -1.488275e-07, -1.487676e-07, 
    -1.490349e-07, -1.491149e-07, -1.49487e-07, -1.493331e-07, -1.495765e-07, 
    -1.493574e-07, -1.493966e-07, -1.495866e-07, -1.493689e-07, 
    -1.498387e-07, -1.495224e-07, -1.501116e-07, -1.497952e-07, 
    -1.501313e-07, -1.500702e-07, -1.501709e-07, -1.502617e-07, 
    -1.503747e-07, -1.505847e-07, -1.505359e-07, -1.507103e-07, 
    -1.489121e-07, -1.490213e-07, -1.490107e-07, -1.491242e-07, 
    -1.492084e-07, -1.493892e-07, -1.496799e-07, -1.495704e-07, 
    -1.497703e-07, -1.498108e-07, -1.495064e-07, -1.496943e-07, 
    -1.490936e-07, -1.491919e-07, -1.491327e-07, -1.489212e-07, -1.49597e-07, 
    -1.492513e-07, -1.498913e-07, -1.49701e-07, -1.502489e-07, -1.499794e-07, 
    -1.505092e-07, -1.507375e-07, -1.509475e-07, -1.511976e-07, 
    -1.490798e-07, -1.490057e-07, -1.491374e-07, -1.493213e-07, 
    -1.494887e-07, -1.497126e-07, -1.49735e-07, -1.497771e-07, -1.498884e-07, 
    -1.499796e-07, -1.497914e-07, -1.500024e-07, -1.492167e-07, 
    -1.496265e-07, -1.489786e-07, -1.491754e-07, -1.4931e-07, -1.4925e-07, 
    -1.495576e-07, -1.496304e-07, -1.499292e-07, -1.497726e-07, 
    -1.506821e-07, -1.502822e-07, -1.513844e-07, -1.510781e-07, 
    -1.489801e-07, -1.490791e-07, -1.494245e-07, -1.492601e-07, -1.49727e-07, 
    -1.498421e-07, -1.499381e-07, -1.50058e-07, -1.500702e-07, -1.501411e-07, 
    -1.500251e-07, -1.501361e-07, -1.497131e-07, -1.49904e-07, -1.493838e-07, 
    -1.495104e-07, -1.494519e-07, -1.493883e-07, -1.495844e-07, 
    -1.497946e-07, -1.497975e-07, -1.498684e-07, -1.500615e-07, 
    -1.497289e-07, -1.507365e-07, -1.5012e-07, -1.49187e-07, -1.493795e-07, 
    -1.494051e-07, -1.493309e-07, -1.498307e-07, -1.4965e-07, -1.501391e-07, 
    -1.500077e-07, -1.502226e-07, -1.50116e-07, -1.501004e-07, -1.499629e-07, 
    -1.498777e-07, -1.496586e-07, -1.494823e-07, -1.493414e-07, 
    -1.493741e-07, -1.495287e-07, -1.498071e-07, -1.500721e-07, -1.50015e-07, 
    -1.502062e-07, -1.496933e-07, -1.499114e-07, -1.498256e-07, 
    -1.500435e-07, -1.495678e-07, -1.499783e-07, -1.494641e-07, 
    -1.495086e-07, -1.496464e-07, -1.49927e-07, -1.499859e-07, -1.500516e-07, 
    -1.500108e-07, -1.498138e-07, -1.497814e-07, -1.496427e-07, 
    -1.496051e-07, -1.494988e-07, -1.494115e-07, -1.494917e-07, 
    -1.495762e-07, -1.498133e-07, -1.500307e-07, -1.502632e-07, 
    -1.503194e-07, -1.505943e-07, -1.503727e-07, -1.507403e-07, 
    -1.504311e-07, -1.509641e-07, -1.499995e-07, -1.504189e-07, 
    -1.496521e-07, -1.497342e-07, -1.498876e-07, -1.502276e-07, 
    -1.500425e-07, -1.502582e-07, -1.4978e-07, -1.495348e-07, -1.494693e-07, 
    -1.493503e-07, -1.49472e-07, -1.494621e-07, -1.495785e-07, -1.49541e-07, 
    -1.498211e-07, -1.496707e-07, -1.501004e-07, -1.502561e-07, 
    -1.506926e-07, -1.509604e-07, -1.512298e-07, -1.513494e-07, 
    -1.513856e-07, -1.514008e-07 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_NODYNLNDUSE =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_R =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.2567e-06, 3.26279e-06, 3.261605e-06, 3.266526e-06, 3.263796e-06, 
    3.267019e-06, 3.257934e-06, 3.263032e-06, 3.259777e-06, 3.257248e-06, 
    3.276056e-06, 3.266745e-06, 3.285764e-06, 3.279803e-06, 3.295445e-06, 
    3.284834e-06, 3.297464e-06, 3.295159e-06, 3.302109e-06, 3.300116e-06, 
    3.309019e-06, 3.303029e-06, 3.313651e-06, 3.307589e-06, 3.308535e-06, 
    3.302831e-06, 3.268619e-06, 3.274895e-06, 3.268247e-06, 3.269141e-06, 
    3.268741e-06, 3.263851e-06, 3.261386e-06, 3.256236e-06, 3.25717e-06, 
    3.260954e-06, 3.269543e-06, 3.266634e-06, 3.273975e-06, 3.273809e-06, 
    3.281998e-06, 3.278304e-06, 3.292744e-06, 3.288177e-06, 3.3002e-06, 
    3.297329e-06, 3.300064e-06, 3.299235e-06, 3.300075e-06, 3.295867e-06, 
    3.297669e-06, 3.29397e-06, 3.278995e-06, 3.2832e-06, 3.270675e-06, 
    3.263149e-06, 3.258157e-06, 3.254619e-06, 3.255119e-06, 3.256072e-06, 
    3.260976e-06, 3.265598e-06, 3.269115e-06, 3.271466e-06, 3.273785e-06, 
    3.280808e-06, 3.284536e-06, 3.293539e-06, 3.292027e-06, 3.29459e-06, 
    3.297044e-06, 3.301167e-06, 3.300488e-06, 3.302305e-06, 3.294524e-06, 
    3.299692e-06, 3.290533e-06, 3.293495e-06, 3.274409e-06, 3.26742e-06, 
    3.264437e-06, 3.261833e-06, 3.255503e-06, 3.259872e-06, 3.258149e-06, 
    3.262252e-06, 3.264862e-06, 3.263571e-06, 3.27153e-06, 3.268439e-06, 
    3.284758e-06, 3.277719e-06, 3.296758e-06, 3.292338e-06, 3.297819e-06, 
    3.29502e-06, 3.299816e-06, 3.2955e-06, 3.302983e-06, 3.304614e-06, 
    3.303499e-06, 3.307788e-06, 3.29526e-06, 3.300063e-06, 3.263535e-06, 
    3.263745e-06, 3.264727e-06, 3.260415e-06, 3.260152e-06, 3.25621e-06, 
    3.259718e-06, 3.261213e-06, 3.265015e-06, 3.267263e-06, 3.269394e-06, 
    3.274087e-06, 3.279334e-06, 3.286689e-06, 3.292624e-06, 3.296186e-06, 
    3.294002e-06, 3.29593e-06, 3.293774e-06, 3.292765e-06, 3.304002e-06, 
    3.297685e-06, 3.30717e-06, 3.306645e-06, 3.302348e-06, 3.306704e-06, 
    3.263893e-06, 3.262682e-06, 3.25848e-06, 3.261768e-06, 3.255781e-06, 
    3.259129e-06, 3.261056e-06, 3.268502e-06, 3.270137e-06, 3.271651e-06, 
    3.274646e-06, 3.278493e-06, 3.285252e-06, 3.291784e-06, 3.297187e-06, 
    3.296791e-06, 3.296931e-06, 3.298138e-06, 3.295146e-06, 3.29863e-06, 
    3.299214e-06, 3.297685e-06, 3.306574e-06, 3.304032e-06, 3.306634e-06, 
    3.304978e-06, 3.263076e-06, 3.265115e-06, 3.264013e-06, 3.266085e-06, 
    3.264624e-06, 3.271105e-06, 3.273047e-06, 3.282156e-06, 3.278417e-06, 
    3.284372e-06, 3.279021e-06, 3.279968e-06, 3.284563e-06, 3.279311e-06, 
    3.290822e-06, 3.283009e-06, 3.298185e-06, 3.289716e-06, 3.298677e-06, 
    3.297164e-06, 3.29967e-06, 3.301916e-06, 3.304746e-06, 3.309973e-06, 
    3.308762e-06, 3.313141e-06, 3.268152e-06, 3.27079e-06, 3.270559e-06, 
    3.273322e-06, 3.275367e-06, 3.279805e-06, 3.286937e-06, 3.284253e-06, 
    3.289184e-06, 3.290174e-06, 3.282685e-06, 3.287279e-06, 3.272557e-06, 
    3.27493e-06, 3.273518e-06, 3.268359e-06, 3.28487e-06, 3.276385e-06, 
    3.292712e-06, 3.287463e-06, 3.301596e-06, 3.294869e-06, 3.308095e-06, 
    3.313764e-06, 3.319121e-06, 3.325383e-06, 3.272232e-06, 3.270438e-06, 
    3.273651e-06, 3.2781e-06, 3.282236e-06, 3.287744e-06, 3.288309e-06, 
    3.289342e-06, 3.292657e-06, 3.294914e-06, 3.289667e-06, 3.29548e-06, 
    3.275478e-06, 3.285608e-06, 3.269759e-06, 3.274522e-06, 3.277838e-06, 
    3.276385e-06, 3.283947e-06, 3.285732e-06, 3.293636e-06, 3.289241e-06, 
    3.312362e-06, 3.302388e-06, 3.330168e-06, 3.322374e-06, 3.269811e-06, 
    3.272226e-06, 3.280642e-06, 3.276636e-06, 3.288113e-06, 3.290945e-06, 
    3.293889e-06, 3.296841e-06, 3.297161e-06, 3.298913e-06, 3.296043e-06, 
    3.2988e-06, 3.287756e-06, 3.293035e-06, 3.27968e-06, 3.282769e-06, 
    3.281348e-06, 3.279789e-06, 3.284603e-06, 3.289739e-06, 3.289852e-06, 
    3.292135e-06, 3.296787e-06, 3.288159e-06, 3.313646e-06, 3.298263e-06, 
    3.274861e-06, 3.279518e-06, 3.280186e-06, 3.278381e-06, 3.290661e-06, 
    3.286204e-06, 3.29887e-06, 3.295612e-06, 3.300954e-06, 3.298297e-06, 
    3.297907e-06, 3.2945e-06, 3.292382e-06, 3.286408e-06, 3.282073e-06, 
    3.278643e-06, 3.27944e-06, 3.28321e-06, 3.290054e-06, 3.297189e-06, 
    3.295763e-06, 3.300547e-06, 3.287279e-06, 3.293199e-06, 3.290518e-06, 
    3.296493e-06, 3.284181e-06, 3.294747e-06, 3.281649e-06, 3.282739e-06, 
    3.286116e-06, 3.293557e-06, 3.29507e-06, 3.296683e-06, 3.295688e-06, 
    3.290229e-06, 3.289441e-06, 3.286034e-06, 3.285093e-06, 3.282502e-06, 
    3.280358e-06, 3.282316e-06, 3.284374e-06, 3.290232e-06, 3.29616e-06, 
    3.301948e-06, 3.303367e-06, 3.310141e-06, 3.304621e-06, 3.313732e-06, 
    3.305978e-06, 3.319418e-06, 3.295328e-06, 3.305757e-06, 3.28627e-06, 
    3.288294e-06, 3.29259e-06, 3.301021e-06, 3.296468e-06, 3.301795e-06, 
    3.289411e-06, 3.283339e-06, 3.281773e-06, 3.278851e-06, 3.28184e-06, 
    3.281597e-06, 3.284461e-06, 3.283541e-06, 3.290427e-06, 3.286726e-06, 
    3.297896e-06, 3.301753e-06, 3.31268e-06, 3.319399e-06, 3.326263e-06, 
    3.329296e-06, 3.33022e-06, 3.330607e-06 ;

 QVEGE =
  -6.482253e-07, -6.477864e-07, -6.478697e-07, -6.475194e-07, -6.477105e-07, 
    -6.474834e-07, -6.481324e-07, -6.477725e-07, -6.480001e-07, 
    -6.481803e-07, -6.468475e-07, -6.475028e-07, -6.461315e-07, 
    -6.465538e-07, -6.454798e-07, -6.462028e-07, -6.453311e-07, 
    -6.454915e-07, -6.449849e-07, -6.451298e-07, -6.444979e-07, 
    -6.449179e-07, -6.44153e-07, -6.445934e-07, -6.445282e-07, -6.449332e-07, 
    -6.473625e-07, -6.469323e-07, -6.4739e-07, -6.473283e-07, -6.473539e-07, 
    -6.477098e-07, -6.478945e-07, -6.482525e-07, -6.48186e-07, -6.479195e-07, 
    -6.473003e-07, -6.47505e-07, -6.469705e-07, -6.469824e-07, -6.463948e-07, 
    -6.466591e-07, -6.456664e-07, -6.459459e-07, -6.451236e-07, 
    -6.453332e-07, -6.451351e-07, -6.45194e-07, -6.451343e-07, -6.454409e-07, 
    -6.453101e-07, -6.455764e-07, -6.466113e-07, -6.463105e-07, 
    -6.472156e-07, -6.477728e-07, -6.481183e-07, -6.483695e-07, 
    -6.483341e-07, -6.482683e-07, -6.479181e-07, -6.475797e-07, 
    -6.473238e-07, -6.471536e-07, -6.469842e-07, -6.464973e-07, -6.4622e-07, 
    -6.456138e-07, -6.457162e-07, -6.455367e-07, -6.453536e-07, 
    -6.450559e-07, -6.451039e-07, -6.449743e-07, -6.455357e-07, 
    -6.451659e-07, -6.457741e-07, -6.456107e-07, -6.469694e-07, 
    -6.474484e-07, -6.476779e-07, -6.478548e-07, -6.483075e-07, 
    -6.479968e-07, -6.481201e-07, -6.478199e-07, -6.476332e-07, 
    -6.477243e-07, -6.471489e-07, -6.473742e-07, -6.462035e-07, 
    -6.467061e-07, -6.453749e-07, -6.456945e-07, -6.45297e-07, -6.454986e-07, 
    -6.451554e-07, -6.454642e-07, -6.449235e-07, -6.448088e-07, 
    -6.448879e-07, -6.445732e-07, -6.454821e-07, -6.45138e-07, -6.477283e-07, 
    -6.477137e-07, -6.476416e-07, -6.479584e-07, -6.479759e-07, 
    -6.482559e-07, -6.48004e-07, -6.478991e-07, -6.476199e-07, -6.474601e-07, 
    -6.473059e-07, -6.469655e-07, -6.465912e-07, -6.4606e-07, -6.456742e-07, 
    -6.454143e-07, -6.455717e-07, -6.45433e-07, -6.455892e-07, -6.45661e-07, 
    -6.448539e-07, -6.453108e-07, -6.446186e-07, -6.44656e-07, -6.449724e-07, 
    -6.446517e-07, -6.477028e-07, -6.477882e-07, -6.48094e-07, -6.478547e-07, 
    -6.482859e-07, -6.480487e-07, -6.479144e-07, -6.473763e-07, 
    -6.472502e-07, -6.471428e-07, -6.469231e-07, -6.466457e-07, 
    -6.461627e-07, -6.457379e-07, -6.453416e-07, -6.453701e-07, 
    -6.453604e-07, -6.452748e-07, -6.454909e-07, -6.45239e-07, -6.451996e-07, 
    -6.453072e-07, -6.446612e-07, -6.448459e-07, -6.446568e-07, 
    -6.447764e-07, -6.477597e-07, -6.476145e-07, -6.476935e-07, 
    -6.475466e-07, -6.476525e-07, -6.471893e-07, -6.470501e-07, 
    -6.463912e-07, -6.466529e-07, -6.462275e-07, -6.466072e-07, 
    -6.465418e-07, -6.462267e-07, -6.465847e-07, -6.457654e-07, 
    -6.463333e-07, -6.452714e-07, -6.458523e-07, -6.452355e-07, 
    -6.453434e-07, -6.451615e-07, -6.450018e-07, -6.447945e-07, 
    -6.444197e-07, -6.445053e-07, -6.441857e-07, -6.473946e-07, 
    -6.472083e-07, -6.472189e-07, -6.470194e-07, -6.468728e-07, 
    -6.465497e-07, -6.460385e-07, -6.462292e-07, -6.458726e-07, 
    -6.458029e-07, -6.463412e-07, -6.460165e-07, -6.470789e-07, 
    -6.469127e-07, -6.470074e-07, -6.473834e-07, -6.461934e-07, -6.46806e-07, 
    -6.456688e-07, -6.459991e-07, -6.450254e-07, -6.455184e-07, 
    -6.445539e-07, -6.441533e-07, -6.437466e-07, -6.433011e-07, 
    -6.471001e-07, -6.472276e-07, -6.46994e-07, -6.466817e-07, -6.463771e-07, 
    -6.4598e-07, -6.459362e-07, -6.458634e-07, -6.456692e-07, -6.455067e-07, 
    -6.45846e-07, -6.454653e-07, -6.468858e-07, -6.461373e-07, -6.472811e-07, 
    -6.469436e-07, -6.466975e-07, -6.46799e-07, -6.462495e-07, -6.461217e-07, 
    -6.456052e-07, -6.458683e-07, -6.442576e-07, -6.449763e-07, 
    -6.429402e-07, -6.435185e-07, -6.472735e-07, -6.470977e-07, 
    -6.464956e-07, -6.4678e-07, -6.459504e-07, -6.457479e-07, -6.455799e-07, 
    -6.453714e-07, -6.453445e-07, -6.452199e-07, -6.454247e-07, 
    -6.452258e-07, -6.459792e-07, -6.456438e-07, -6.465571e-07, 
    -6.463385e-07, -6.464372e-07, -6.465496e-07, -6.46203e-07, -6.458421e-07, 
    -6.458249e-07, -6.457126e-07, -6.45406e-07, -6.459468e-07, -6.441819e-07, 
    -6.452947e-07, -6.469064e-07, -6.465815e-07, -6.465239e-07, 
    -6.466513e-07, -6.457686e-07, -6.460903e-07, -6.452216e-07, -6.45456e-07, 
    -6.450691e-07, -6.452625e-07, -6.452913e-07, -6.455365e-07, 
    -6.456914e-07, -6.460774e-07, -6.463896e-07, -6.466316e-07, 
    -6.465746e-07, -6.463084e-07, -6.458178e-07, -6.453463e-07, 
    -6.454516e-07, -6.450985e-07, -6.460111e-07, -6.456359e-07, -6.45783e-07, 
    -6.453938e-07, -6.462364e-07, -6.455484e-07, -6.464153e-07, 
    -6.463375e-07, -6.460966e-07, -6.456166e-07, -6.454954e-07, 
    -6.453829e-07, -6.454504e-07, -6.458035e-07, -6.458574e-07, 
    -6.461002e-07, -6.461719e-07, -6.463537e-07, -6.465084e-07, 
    -6.463695e-07, -6.462253e-07, -6.457995e-07, -6.454213e-07, 
    -6.450009e-07, -6.44894e-07, -6.444232e-07, -6.448198e-07, -6.441776e-07, 
    -6.447437e-07, -6.437511e-07, -6.454943e-07, -6.44741e-07, -6.460825e-07, 
    -6.459367e-07, -6.456844e-07, -6.45077e-07, -6.453955e-07, -6.450182e-07, 
    -6.458587e-07, -6.463039e-07, -6.464071e-07, -6.466186e-07, 
    -6.464023e-07, -6.464195e-07, -6.462126e-07, -6.462786e-07, 
    -6.457852e-07, -6.4605e-07, -6.452946e-07, -6.450188e-07, -6.442227e-07, 
    -6.437367e-07, -6.432232e-07, -6.430006e-07, -6.429318e-07, -6.429037e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.71156, 84.71111, 84.7112, 84.71084, 84.71104, 84.7108, 84.71146, 
    84.71109, 84.71133, 84.71152, 84.71021, 84.71082, 84.70963, 84.70997, 
    84.70869, 84.70968, 84.70859, 84.70871, 84.70834, 84.70845, 84.708, 
    84.7083, 84.70778, 84.70807, 84.70802, 84.70831, 84.71069, 84.71028, 
    84.71072, 84.71066, 84.71069, 84.71103, 84.71121, 84.71159, 84.71152, 
    84.71124, 84.71063, 84.71083, 84.71033, 84.71034, 84.70984, 84.71005, 
    84.70884, 84.70949, 84.70844, 84.7086, 84.70845, 84.7085, 84.70845, 
    84.70867, 84.70857, 84.70877, 84.71001, 84.70977, 84.71055, 84.71109, 
    84.71145, 84.71172, 84.71168, 84.71161, 84.71124, 84.7109, 84.71066, 
    84.71049, 84.71034, 84.70992, 84.70969, 84.70879, 84.70888, 84.70874, 
    84.70861, 84.7084, 84.70843, 84.70834, 84.70874, 84.70847, 84.70936, 
    84.70879, 84.71031, 84.71077, 84.71099, 84.71117, 84.71165, 84.71132, 
    84.71145, 84.71114, 84.71095, 84.71104, 84.71049, 84.7107, 84.70969, 
    84.71009, 84.70863, 84.70885, 84.70856, 84.70872, 84.70847, 84.70869, 
    84.70831, 84.70822, 84.70827, 84.70806, 84.7087, 84.70845, 84.71105, 
    84.71104, 84.71096, 84.71128, 84.7113, 84.71159, 84.71133, 84.71122, 
    84.71095, 84.71078, 84.71064, 84.71032, 84.70999, 84.70957, 84.70884, 
    84.70866, 84.70877, 84.70866, 84.70878, 84.70883, 84.70825, 84.70857, 
    84.70809, 84.70811, 84.70834, 84.70811, 84.71103, 84.71111, 84.71143, 
    84.71118, 84.71162, 84.71138, 84.71124, 84.7107, 84.71059, 84.71049, 
    84.71028, 84.71004, 84.70966, 84.70889, 84.7086, 84.70862, 84.70861, 
    84.70855, 84.70871, 84.70853, 84.7085, 84.70857, 84.70812, 84.70825, 
    84.70811, 84.7082, 84.71108, 84.71094, 84.71101, 84.71087, 84.71098, 
    84.71053, 84.7104, 84.70983, 84.71004, 84.7097, 84.71001, 84.70995, 
    84.70969, 84.70999, 84.70935, 84.70979, 84.70855, 84.70941, 84.70853, 
    84.7086, 84.70847, 84.70836, 84.70821, 84.70795, 84.70802, 84.7078, 
    84.71072, 84.71055, 84.71056, 84.71037, 84.71024, 84.70996, 84.70956, 
    84.70971, 84.70943, 84.70938, 84.7098, 84.70954, 84.71043, 84.71027, 
    84.71036, 84.71071, 84.70968, 84.71017, 84.70884, 84.70953, 84.70837, 
    84.70872, 84.70805, 84.70777, 84.70752, 84.70724, 84.71045, 84.71056, 
    84.71035, 84.71007, 84.70982, 84.70951, 84.70948, 84.70943, 84.70884, 
    84.70872, 84.70941, 84.70869, 84.71024, 84.70963, 84.71062, 84.7103, 
    84.71008, 84.71017, 84.70972, 84.70963, 84.70879, 84.70943, 84.70784, 
    84.70834, 84.70702, 84.70737, 84.71061, 84.71044, 84.70992, 84.71015, 
    84.7095, 84.70934, 84.70878, 84.70862, 84.7086, 84.70851, 84.70866, 
    84.70852, 84.70951, 84.70882, 84.70997, 84.70979, 84.70988, 84.70996, 
    84.70969, 84.7094, 84.7094, 84.70887, 84.70863, 84.70949, 84.70779, 
    84.70856, 84.71027, 84.70998, 84.70995, 84.71004, 84.70936, 84.7096, 
    84.70851, 84.70869, 84.7084, 84.70854, 84.70856, 84.70874, 84.70885, 
    84.70959, 84.70983, 84.71003, 84.70998, 84.70977, 84.70939, 84.7086, 
    84.70868, 84.70843, 84.70954, 84.70882, 84.70937, 84.70864, 84.70972, 
    84.70874, 84.70985, 84.70979, 84.7096, 84.70879, 84.70871, 84.70863, 
    84.70868, 84.70938, 84.70942, 84.70961, 84.70966, 84.70981, 84.70993, 
    84.70982, 84.7097, 84.70938, 84.70866, 84.70835, 84.70828, 84.70795, 
    84.70822, 84.70778, 84.70816, 84.70751, 84.7087, 84.70817, 84.70959, 
    84.70948, 84.70885, 84.7084, 84.70864, 84.70837, 84.70943, 84.70976, 
    84.70985, 84.71002, 84.70985, 84.70986, 84.70969, 84.70975, 84.70937, 
    84.70957, 84.70856, 84.70837, 84.70782, 84.7075, 84.70719, 84.70706, 
    84.70702, 84.707 ;

 RH2M_R =
  84.71156, 84.71111, 84.7112, 84.71084, 84.71104, 84.7108, 84.71146, 
    84.71109, 84.71133, 84.71152, 84.71021, 84.71082, 84.70963, 84.70997, 
    84.70869, 84.70968, 84.70859, 84.70871, 84.70834, 84.70845, 84.708, 
    84.7083, 84.70778, 84.70807, 84.70802, 84.70831, 84.71069, 84.71028, 
    84.71072, 84.71066, 84.71069, 84.71103, 84.71121, 84.71159, 84.71152, 
    84.71124, 84.71063, 84.71083, 84.71033, 84.71034, 84.70984, 84.71005, 
    84.70884, 84.70949, 84.70844, 84.7086, 84.70845, 84.7085, 84.70845, 
    84.70867, 84.70857, 84.70877, 84.71001, 84.70977, 84.71055, 84.71109, 
    84.71145, 84.71172, 84.71168, 84.71161, 84.71124, 84.7109, 84.71066, 
    84.71049, 84.71034, 84.70992, 84.70969, 84.70879, 84.70888, 84.70874, 
    84.70861, 84.7084, 84.70843, 84.70834, 84.70874, 84.70847, 84.70936, 
    84.70879, 84.71031, 84.71077, 84.71099, 84.71117, 84.71165, 84.71132, 
    84.71145, 84.71114, 84.71095, 84.71104, 84.71049, 84.7107, 84.70969, 
    84.71009, 84.70863, 84.70885, 84.70856, 84.70872, 84.70847, 84.70869, 
    84.70831, 84.70822, 84.70827, 84.70806, 84.7087, 84.70845, 84.71105, 
    84.71104, 84.71096, 84.71128, 84.7113, 84.71159, 84.71133, 84.71122, 
    84.71095, 84.71078, 84.71064, 84.71032, 84.70999, 84.70957, 84.70884, 
    84.70866, 84.70877, 84.70866, 84.70878, 84.70883, 84.70825, 84.70857, 
    84.70809, 84.70811, 84.70834, 84.70811, 84.71103, 84.71111, 84.71143, 
    84.71118, 84.71162, 84.71138, 84.71124, 84.7107, 84.71059, 84.71049, 
    84.71028, 84.71004, 84.70966, 84.70889, 84.7086, 84.70862, 84.70861, 
    84.70855, 84.70871, 84.70853, 84.7085, 84.70857, 84.70812, 84.70825, 
    84.70811, 84.7082, 84.71108, 84.71094, 84.71101, 84.71087, 84.71098, 
    84.71053, 84.7104, 84.70983, 84.71004, 84.7097, 84.71001, 84.70995, 
    84.70969, 84.70999, 84.70935, 84.70979, 84.70855, 84.70941, 84.70853, 
    84.7086, 84.70847, 84.70836, 84.70821, 84.70795, 84.70802, 84.7078, 
    84.71072, 84.71055, 84.71056, 84.71037, 84.71024, 84.70996, 84.70956, 
    84.70971, 84.70943, 84.70938, 84.7098, 84.70954, 84.71043, 84.71027, 
    84.71036, 84.71071, 84.70968, 84.71017, 84.70884, 84.70953, 84.70837, 
    84.70872, 84.70805, 84.70777, 84.70752, 84.70724, 84.71045, 84.71056, 
    84.71035, 84.71007, 84.70982, 84.70951, 84.70948, 84.70943, 84.70884, 
    84.70872, 84.70941, 84.70869, 84.71024, 84.70963, 84.71062, 84.7103, 
    84.71008, 84.71017, 84.70972, 84.70963, 84.70879, 84.70943, 84.70784, 
    84.70834, 84.70702, 84.70737, 84.71061, 84.71044, 84.70992, 84.71015, 
    84.7095, 84.70934, 84.70878, 84.70862, 84.7086, 84.70851, 84.70866, 
    84.70852, 84.70951, 84.70882, 84.70997, 84.70979, 84.70988, 84.70996, 
    84.70969, 84.7094, 84.7094, 84.70887, 84.70863, 84.70949, 84.70779, 
    84.70856, 84.71027, 84.70998, 84.70995, 84.71004, 84.70936, 84.7096, 
    84.70851, 84.70869, 84.7084, 84.70854, 84.70856, 84.70874, 84.70885, 
    84.70959, 84.70983, 84.71003, 84.70998, 84.70977, 84.70939, 84.7086, 
    84.70868, 84.70843, 84.70954, 84.70882, 84.70937, 84.70864, 84.70972, 
    84.70874, 84.70985, 84.70979, 84.7096, 84.70879, 84.70871, 84.70863, 
    84.70868, 84.70938, 84.70942, 84.70961, 84.70966, 84.70981, 84.70993, 
    84.70982, 84.7097, 84.70938, 84.70866, 84.70835, 84.70828, 84.70795, 
    84.70822, 84.70778, 84.70816, 84.70751, 84.7087, 84.70817, 84.70959, 
    84.70948, 84.70885, 84.7084, 84.70864, 84.70837, 84.70943, 84.70976, 
    84.70985, 84.71002, 84.70985, 84.70986, 84.70969, 84.70975, 84.70937, 
    84.70957, 84.70856, 84.70837, 84.70782, 84.7075, 84.70719, 84.70706, 
    84.70702, 84.707 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004631331, 0.0004650735, 0.0004646961, 0.0004662612, 0.0004653929, 
    0.0004664176, 0.0004635262, 0.0004651503, 0.0004641133, 0.0004633072, 
    0.0004692978, 0.0004663305, 0.0004723785, 0.0004704865, 0.0004752382, 
    0.000472084, 0.000475874, 0.0004751468, 0.0004773345, 0.0004767077, 
    0.000479506, 0.0004776236, 0.000480956, 0.0004790563, 0.0004793535, 
    0.0004775613, 0.0004669279, 0.0004689289, 0.0004668093, 0.0004670946, 
    0.0004669664, 0.0004654107, 0.0004646268, 0.0004629842, 0.0004632823, 
    0.0004644885, 0.0004672225, 0.0004662942, 0.0004686329, 0.0004685801, 
    0.0004711834, 0.0004700096, 0.0004743846, 0.0004731411, 0.0004767338, 
    0.0004758303, 0.0004766913, 0.0004764301, 0.0004766945, 0.0004753695, 
    0.0004759372, 0.0004747711, 0.0004702302, 0.0004715652, 0.0004675831, 
    0.0004651885, 0.0004635972, 0.0004624682, 0.0004626277, 0.000462932, 
    0.0004644955, 0.0004659652, 0.0004670851, 0.0004678343, 0.0004685723, 
    0.000470807, 0.0004719891, 0.0004746361, 0.0004741582, 0.0004749675, 
    0.0004757403, 0.0004770381, 0.0004768244, 0.0004773962, 0.0004749456, 
    0.0004765744, 0.0004738855, 0.000474621, 0.0004687743, 0.0004665449, 
    0.0004655978, 0.0004647682, 0.0004627504, 0.0004641439, 0.0004635945, 
    0.000464901, 0.0004657313, 0.0004653205, 0.0004678547, 0.0004668694, 
    0.0004720591, 0.0004698239, 0.0004756503, 0.0004742561, 0.0004759842, 
    0.0004751023, 0.0004766133, 0.0004752534, 0.0004776088, 0.0004781218, 
    0.0004777711, 0.0004791173, 0.0004751777, 0.0004766908, 0.0004653094, 
    0.0004653764, 0.0004656883, 0.0004643168, 0.0004642329, 0.0004629757, 
    0.0004640941, 0.0004645705, 0.0004657792, 0.0004664943, 0.0004671739, 
    0.0004686684, 0.0004703373, 0.0004726705, 0.0004743464, 0.0004754697, 
    0.0004747808, 0.0004753889, 0.000474709, 0.0004743902, 0.0004779295, 
    0.0004759423, 0.0004789236, 0.0004787586, 0.0004774094, 0.000478777, 
    0.0004654233, 0.0004650378, 0.0004636997, 0.0004647468, 0.0004628387, 
    0.0004639068, 0.000464521, 0.0004668902, 0.0004674104, 0.0004678931, 
    0.0004688462, 0.0004700693, 0.0004722149, 0.0004740814, 0.0004757851, 
    0.0004756601, 0.0004757041, 0.0004760846, 0.0004751418, 0.0004762393, 
    0.0004764235, 0.0004759418, 0.0004787363, 0.000477938, 0.0004787548, 
    0.0004782349, 0.000465163, 0.0004658114, 0.0004654609, 0.0004661199, 
    0.0004656556, 0.0004677198, 0.0004683386, 0.0004712337, 0.0004700453, 
    0.0004719362, 0.0004702372, 0.0004705383, 0.0004719981, 0.0004703288, 
    0.0004739785, 0.0004715044, 0.0004760993, 0.0004736294, 0.000476254, 
    0.0004757772, 0.0004765663, 0.0004772732, 0.0004781622, 0.0004798028, 
    0.0004794228, 0.0004807946, 0.000466778, 0.0004676191, 0.0004675449, 
    0.0004684249, 0.0004690758, 0.0004704863, 0.0004727485, 0.0004718977, 
    0.0004734592, 0.0004737727, 0.0004714001, 0.000472857, 0.0004681814, 
    0.0004689369, 0.0004684869, 0.0004668436, 0.0004720935, 0.0004693994, 
    0.0004743735, 0.0004729142, 0.0004771723, 0.000475055, 0.0004792136, 
    0.0004809916, 0.0004826639, 0.0004846189, 0.000468078, 0.0004675064, 
    0.0004685294, 0.0004699452, 0.0004712582, 0.0004730039, 0.0004731824, 
    0.0004735094, 0.0004743563, 0.0004750685, 0.0004736128, 0.0004752468, 
    0.0004691124, 0.0004723272, 0.0004672897, 0.0004688069, 0.0004698609, 
    0.0004693984, 0.0004717997, 0.0004723656, 0.0004746653, 0.0004734764, 
    0.0004805528, 0.0004774223, 0.0004861067, 0.0004836803, 0.0004673066, 
    0.0004680757, 0.0004707524, 0.0004694788, 0.0004731202, 0.0004740165, 
    0.0004747449, 0.0004756763, 0.0004757766, 0.0004763284, 0.0004754241, 
    0.0004762925, 0.000473007, 0.0004744753, 0.0004704456, 0.0004714265, 
    0.0004709752, 0.0004704801, 0.0004720076, 0.0004736351, 0.0004736696, 
    0.0004741914, 0.0004756623, 0.000473134, 0.000480957, 0.0004761264, 
    0.0004689143, 0.0004703958, 0.000470607, 0.0004700332, 0.0004739265, 
    0.0004725159, 0.0004763149, 0.0004752881, 0.0004769702, 0.0004761344, 
    0.0004760113, 0.0004749376, 0.0004742691, 0.0004725802, 0.0004712058, 
    0.0004701157, 0.0004703691, 0.0004715664, 0.0004737345, 0.0004757851, 
    0.0004753359, 0.0004768417, 0.0004728551, 0.000474527, 0.0004738808, 
    0.0004755653, 0.0004718749, 0.0004750193, 0.0004710711, 0.0004714172, 
    0.0004724878, 0.0004746414, 0.0004751173, 0.0004756261, 0.000475312, 
    0.0004737899, 0.0004735403, 0.0004724613, 0.0004721635, 0.0004713413, 
    0.0004706605, 0.0004712825, 0.0004719355, 0.00047379, 0.000475461, 
    0.0004772827, 0.0004777283, 0.0004798571, 0.0004781244, 0.0004809837, 
    0.0004785533, 0.0004827599, 0.000475201, 0.0004784824, 0.0004725364, 
    0.0004731769, 0.0004743358, 0.0004769929, 0.0004755581, 0.0004772359, 
    0.0004735305, 0.000471608, 0.0004711101, 0.000470182, 0.0004711313, 
    0.0004710541, 0.0004719624, 0.0004716704, 0.0004738514, 0.0004726799, 
    0.0004760076, 0.0004772219, 0.0004806503, 0.0004827518, 0.0004848903, 
    0.0004858344, 0.0004861217, 0.0004862418 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.113387e-14, 3.121816e-14, 3.120179e-14, 3.126972e-14, 3.123206e-14, 
    3.127652e-14, 3.115098e-14, 3.12215e-14, 3.117649e-14, 3.114148e-14, 
    3.140134e-14, 3.127275e-14, 3.153481e-14, 3.145295e-14, 3.165846e-14, 
    3.152206e-14, 3.168595e-14, 3.165456e-14, 3.174906e-14, 3.1722e-14, 
    3.184269e-14, 3.176155e-14, 3.190522e-14, 3.182333e-14, 3.183614e-14, 
    3.175886e-14, 3.129867e-14, 3.138533e-14, 3.129353e-14, 3.130589e-14, 
    3.130035e-14, 3.123282e-14, 3.119875e-14, 3.112744e-14, 3.11404e-14, 
    3.119278e-14, 3.131145e-14, 3.127121e-14, 3.137266e-14, 3.137037e-14, 
    3.148314e-14, 3.143231e-14, 3.162162e-14, 3.156788e-14, 3.172313e-14, 
    3.168411e-14, 3.17213e-14, 3.171002e-14, 3.172144e-14, 3.16642e-14, 
    3.168873e-14, 3.163835e-14, 3.144183e-14, 3.149963e-14, 3.132709e-14, 
    3.122313e-14, 3.115407e-14, 3.110501e-14, 3.111195e-14, 3.112516e-14, 
    3.119309e-14, 3.125693e-14, 3.130553e-14, 3.133803e-14, 3.137004e-14, 
    3.146677e-14, 3.151798e-14, 3.163247e-14, 3.161185e-14, 3.164681e-14, 
    3.168023e-14, 3.173627e-14, 3.172705e-14, 3.175173e-14, 3.16459e-14, 
    3.171624e-14, 3.160011e-14, 3.163187e-14, 3.137864e-14, 3.128207e-14, 
    3.124091e-14, 3.120493e-14, 3.111728e-14, 3.117782e-14, 3.115396e-14, 
    3.121073e-14, 3.124678e-14, 3.122896e-14, 3.133892e-14, 3.129618e-14, 
    3.152102e-14, 3.142425e-14, 3.167633e-14, 3.161608e-14, 3.169077e-14, 
    3.165267e-14, 3.171793e-14, 3.16592e-14, 3.176092e-14, 3.178304e-14, 
    3.176792e-14, 3.182601e-14, 3.165594e-14, 3.172129e-14, 3.122845e-14, 
    3.123136e-14, 3.124491e-14, 3.118533e-14, 3.118169e-14, 3.112708e-14, 
    3.117568e-14, 3.119636e-14, 3.124888e-14, 3.12799e-14, 3.130939e-14, 
    3.13742e-14, 3.144649e-14, 3.15475e-14, 3.161999e-14, 3.166855e-14, 
    3.163878e-14, 3.166506e-14, 3.163568e-14, 3.162191e-14, 3.177474e-14, 
    3.168895e-14, 3.181766e-14, 3.181055e-14, 3.175231e-14, 3.181135e-14, 
    3.12334e-14, 3.121667e-14, 3.115854e-14, 3.120404e-14, 3.112114e-14, 
    3.116754e-14, 3.11942e-14, 3.129705e-14, 3.131966e-14, 3.134058e-14, 
    3.138191e-14, 3.143491e-14, 3.15278e-14, 3.160852e-14, 3.168218e-14, 
    3.167678e-14, 3.167868e-14, 3.169512e-14, 3.165439e-14, 3.17018e-14, 
    3.170975e-14, 3.168896e-14, 3.180959e-14, 3.177515e-14, 3.181039e-14, 
    3.178797e-14, 3.122212e-14, 3.125026e-14, 3.123505e-14, 3.126365e-14, 
    3.124349e-14, 3.133303e-14, 3.135986e-14, 3.14853e-14, 3.143387e-14, 
    3.151573e-14, 3.144219e-14, 3.145522e-14, 3.151835e-14, 3.144618e-14, 
    3.160407e-14, 3.149702e-14, 3.169575e-14, 3.158895e-14, 3.170244e-14, 
    3.168186e-14, 3.171594e-14, 3.174645e-14, 3.178483e-14, 3.185556e-14, 
    3.183919e-14, 3.189833e-14, 3.129222e-14, 3.132868e-14, 3.132549e-14, 
    3.136365e-14, 3.139186e-14, 3.145298e-14, 3.155089e-14, 3.151409e-14, 
    3.158166e-14, 3.159521e-14, 3.149257e-14, 3.155559e-14, 3.135309e-14, 
    3.138582e-14, 3.136635e-14, 3.129508e-14, 3.152255e-14, 3.140588e-14, 
    3.162118e-14, 3.15581e-14, 3.17421e-14, 3.165062e-14, 3.183018e-14, 
    3.190676e-14, 3.197885e-14, 3.206291e-14, 3.13486e-14, 3.132382e-14, 
    3.136819e-14, 3.14295e-14, 3.14864e-14, 3.156195e-14, 3.156968e-14, 
    3.158382e-14, 3.162044e-14, 3.165122e-14, 3.158827e-14, 3.165893e-14, 
    3.139338e-14, 3.153268e-14, 3.131444e-14, 3.13802e-14, 3.14259e-14, 
    3.140587e-14, 3.150989e-14, 3.153438e-14, 3.16338e-14, 3.158244e-14, 
    3.188785e-14, 3.175286e-14, 3.212692e-14, 3.202256e-14, 3.131516e-14, 
    3.134852e-14, 3.146448e-14, 3.140933e-14, 3.1567e-14, 3.160575e-14, 
    3.163724e-14, 3.167746e-14, 3.168182e-14, 3.170564e-14, 3.16666e-14, 
    3.170411e-14, 3.156211e-14, 3.162559e-14, 3.145126e-14, 3.149372e-14, 
    3.14742e-14, 3.145276e-14, 3.151889e-14, 3.158926e-14, 3.15908e-14, 
    3.161332e-14, 3.167676e-14, 3.156764e-14, 3.19052e-14, 3.169684e-14, 
    3.138488e-14, 3.144902e-14, 3.145822e-14, 3.143337e-14, 3.160187e-14, 
    3.154085e-14, 3.170507e-14, 3.166072e-14, 3.173338e-14, 3.169728e-14, 
    3.169196e-14, 3.164558e-14, 3.161668e-14, 3.154365e-14, 3.148416e-14, 
    3.143698e-14, 3.144795e-14, 3.149978e-14, 3.159357e-14, 3.16822e-14, 
    3.166279e-14, 3.172786e-14, 3.155558e-14, 3.162784e-14, 3.159992e-14, 
    3.167273e-14, 3.151311e-14, 3.164896e-14, 3.147833e-14, 3.149331e-14, 
    3.153964e-14, 3.163272e-14, 3.165334e-14, 3.167531e-14, 3.166176e-14, 
    3.159596e-14, 3.158518e-14, 3.153852e-14, 3.152562e-14, 3.149005e-14, 
    3.146058e-14, 3.14875e-14, 3.151576e-14, 3.1596e-14, 3.16682e-14, 
    3.174688e-14, 3.176613e-14, 3.185786e-14, 3.178316e-14, 3.190635e-14, 
    3.180156e-14, 3.19829e-14, 3.165687e-14, 3.179854e-14, 3.154176e-14, 
    3.156947e-14, 3.161952e-14, 3.17343e-14, 3.167239e-14, 3.174481e-14, 
    3.158476e-14, 3.150155e-14, 3.148004e-14, 3.143984e-14, 3.148096e-14, 
    3.147762e-14, 3.151695e-14, 3.150431e-14, 3.159866e-14, 3.1548e-14, 
    3.169182e-14, 3.174424e-14, 3.189212e-14, 3.198262e-14, 3.207467e-14, 
    3.211526e-14, 3.212761e-14, 3.213277e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.035197e-14, 1.038003e-14, 1.037458e-14, 1.039719e-14, 1.038465e-14, 
    1.039945e-14, 1.035767e-14, 1.038114e-14, 1.036616e-14, 1.035451e-14, 
    1.044099e-14, 1.03982e-14, 1.048542e-14, 1.045817e-14, 1.052657e-14, 
    1.048117e-14, 1.053572e-14, 1.052527e-14, 1.055673e-14, 1.054772e-14, 
    1.058789e-14, 1.056088e-14, 1.06087e-14, 1.058145e-14, 1.058571e-14, 
    1.055999e-14, 1.040682e-14, 1.043567e-14, 1.040511e-14, 1.040923e-14, 
    1.040738e-14, 1.038491e-14, 1.037357e-14, 1.034984e-14, 1.035415e-14, 
    1.037158e-14, 1.041108e-14, 1.039768e-14, 1.043145e-14, 1.043069e-14, 
    1.046822e-14, 1.04513e-14, 1.051431e-14, 1.049642e-14, 1.05481e-14, 
    1.053511e-14, 1.054748e-14, 1.054373e-14, 1.054753e-14, 1.052848e-14, 
    1.053665e-14, 1.051988e-14, 1.045447e-14, 1.047371e-14, 1.041628e-14, 
    1.038168e-14, 1.03587e-14, 1.034237e-14, 1.034468e-14, 1.034908e-14, 
    1.037168e-14, 1.039293e-14, 1.040911e-14, 1.041992e-14, 1.043058e-14, 
    1.046277e-14, 1.047982e-14, 1.051792e-14, 1.051106e-14, 1.052269e-14, 
    1.053382e-14, 1.055247e-14, 1.05494e-14, 1.055761e-14, 1.052239e-14, 
    1.05458e-14, 1.050715e-14, 1.051772e-14, 1.043344e-14, 1.04013e-14, 
    1.03876e-14, 1.037563e-14, 1.034645e-14, 1.03666e-14, 1.035866e-14, 
    1.037756e-14, 1.038955e-14, 1.038362e-14, 1.042022e-14, 1.0406e-14, 
    1.048083e-14, 1.044862e-14, 1.053252e-14, 1.051247e-14, 1.053732e-14, 
    1.052464e-14, 1.054636e-14, 1.052682e-14, 1.056067e-14, 1.056803e-14, 
    1.0563e-14, 1.058234e-14, 1.052573e-14, 1.054748e-14, 1.038345e-14, 
    1.038442e-14, 1.038893e-14, 1.03691e-14, 1.036789e-14, 1.034972e-14, 
    1.036589e-14, 1.037277e-14, 1.039025e-14, 1.040058e-14, 1.041039e-14, 
    1.043196e-14, 1.045602e-14, 1.048964e-14, 1.051377e-14, 1.052993e-14, 
    1.052002e-14, 1.052877e-14, 1.051899e-14, 1.051441e-14, 1.056527e-14, 
    1.053672e-14, 1.057956e-14, 1.057719e-14, 1.055781e-14, 1.057746e-14, 
    1.03851e-14, 1.037953e-14, 1.036018e-14, 1.037533e-14, 1.034774e-14, 
    1.036318e-14, 1.037205e-14, 1.040629e-14, 1.041381e-14, 1.042077e-14, 
    1.043453e-14, 1.045217e-14, 1.048308e-14, 1.050995e-14, 1.053446e-14, 
    1.053267e-14, 1.05333e-14, 1.053877e-14, 1.052522e-14, 1.0541e-14, 
    1.054364e-14, 1.053672e-14, 1.057687e-14, 1.056541e-14, 1.057714e-14, 
    1.056968e-14, 1.038134e-14, 1.039071e-14, 1.038565e-14, 1.039517e-14, 
    1.038846e-14, 1.041826e-14, 1.042719e-14, 1.046894e-14, 1.045182e-14, 
    1.047907e-14, 1.045459e-14, 1.045893e-14, 1.047994e-14, 1.045592e-14, 
    1.050847e-14, 1.047284e-14, 1.053898e-14, 1.050344e-14, 1.054121e-14, 
    1.053436e-14, 1.05457e-14, 1.055586e-14, 1.056863e-14, 1.059217e-14, 
    1.058673e-14, 1.060641e-14, 1.040467e-14, 1.041681e-14, 1.041575e-14, 
    1.042845e-14, 1.043784e-14, 1.045818e-14, 1.049077e-14, 1.047852e-14, 
    1.050101e-14, 1.050552e-14, 1.047136e-14, 1.049233e-14, 1.042494e-14, 
    1.043583e-14, 1.042935e-14, 1.040563e-14, 1.048134e-14, 1.044251e-14, 
    1.051416e-14, 1.049317e-14, 1.055441e-14, 1.052396e-14, 1.058372e-14, 
    1.060921e-14, 1.063321e-14, 1.066119e-14, 1.042344e-14, 1.04152e-14, 
    1.042996e-14, 1.045037e-14, 1.04693e-14, 1.049445e-14, 1.049702e-14, 
    1.050173e-14, 1.051392e-14, 1.052416e-14, 1.050321e-14, 1.052673e-14, 
    1.043834e-14, 1.048471e-14, 1.041207e-14, 1.043396e-14, 1.044917e-14, 
    1.04425e-14, 1.047712e-14, 1.048527e-14, 1.051836e-14, 1.050127e-14, 
    1.060292e-14, 1.055799e-14, 1.068249e-14, 1.064776e-14, 1.041231e-14, 
    1.042341e-14, 1.046201e-14, 1.044365e-14, 1.049613e-14, 1.050903e-14, 
    1.051951e-14, 1.05329e-14, 1.053435e-14, 1.054228e-14, 1.052928e-14, 
    1.054176e-14, 1.04945e-14, 1.051563e-14, 1.045761e-14, 1.047174e-14, 
    1.046524e-14, 1.045811e-14, 1.048012e-14, 1.050354e-14, 1.050405e-14, 
    1.051155e-14, 1.053266e-14, 1.049634e-14, 1.060869e-14, 1.053934e-14, 
    1.043552e-14, 1.045686e-14, 1.045992e-14, 1.045166e-14, 1.050774e-14, 
    1.048743e-14, 1.054208e-14, 1.052732e-14, 1.055151e-14, 1.053949e-14, 
    1.053772e-14, 1.052228e-14, 1.051267e-14, 1.048836e-14, 1.046856e-14, 
    1.045286e-14, 1.045651e-14, 1.047376e-14, 1.050497e-14, 1.053447e-14, 
    1.052801e-14, 1.054967e-14, 1.049233e-14, 1.051638e-14, 1.050709e-14, 
    1.053132e-14, 1.047819e-14, 1.052341e-14, 1.046662e-14, 1.047161e-14, 
    1.048702e-14, 1.0518e-14, 1.052487e-14, 1.053218e-14, 1.052767e-14, 
    1.050577e-14, 1.050218e-14, 1.048665e-14, 1.048236e-14, 1.047052e-14, 
    1.046071e-14, 1.046967e-14, 1.047907e-14, 1.050578e-14, 1.052981e-14, 
    1.0556e-14, 1.056241e-14, 1.059294e-14, 1.056807e-14, 1.060908e-14, 
    1.05742e-14, 1.063455e-14, 1.052604e-14, 1.057319e-14, 1.048773e-14, 
    1.049695e-14, 1.051361e-14, 1.055181e-14, 1.053121e-14, 1.055531e-14, 
    1.050204e-14, 1.047435e-14, 1.046719e-14, 1.045381e-14, 1.04675e-14, 
    1.046638e-14, 1.047947e-14, 1.047527e-14, 1.050667e-14, 1.048981e-14, 
    1.053768e-14, 1.055512e-14, 1.060434e-14, 1.063446e-14, 1.06651e-14, 
    1.067861e-14, 1.068272e-14, 1.068444e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.364721e-11, -8.401534e-11, -8.394378e-11, -8.42407e-11, -8.407599e-11, 
    -8.427042e-11, -8.372185e-11, -8.402996e-11, -8.383327e-11, 
    -8.368035e-11, -8.481693e-11, -8.425394e-11, -8.540167e-11, 
    -8.504263e-11, -8.594454e-11, -8.534581e-11, -8.606527e-11, 
    -8.592726e-11, -8.63426e-11, -8.622361e-11, -8.675488e-11, -8.639752e-11, 
    -8.703026e-11, -8.666953e-11, -8.672597e-11, -8.638573e-11, 
    -8.436724e-11, -8.474684e-11, -8.434475e-11, -8.439888e-11, 
    -8.437458e-11, -8.407939e-11, -8.393064e-11, -8.361907e-11, 
    -8.367564e-11, -8.390447e-11, -8.442322e-11, -8.424712e-11, 
    -8.469091e-11, -8.468089e-11, -8.517495e-11, -8.495219e-11, 
    -8.578258e-11, -8.554657e-11, -8.622858e-11, -8.605706e-11, 
    -8.622052e-11, -8.617096e-11, -8.622117e-11, -8.596962e-11, -8.60774e-11, 
    -8.585604e-11, -8.499391e-11, -8.52473e-11, -8.449159e-11, -8.403719e-11, 
    -8.373537e-11, -8.352118e-11, -8.355146e-11, -8.360918e-11, 
    -8.390581e-11, -8.418468e-11, -8.43972e-11, -8.453937e-11, -8.467944e-11, 
    -8.510346e-11, -8.532786e-11, -8.583032e-11, -8.573963e-11, 
    -8.589325e-11, -8.604e-11, -8.628639e-11, -8.624583e-11, -8.635439e-11, 
    -8.588919e-11, -8.619837e-11, -8.568798e-11, -8.582757e-11, 
    -8.471756e-11, -8.429463e-11, -8.411489e-11, -8.395754e-11, 
    -8.357474e-11, -8.38391e-11, -8.373489e-11, -8.398279e-11, -8.414033e-11, 
    -8.406241e-11, -8.454326e-11, -8.435632e-11, -8.534116e-11, 
    -8.491696e-11, -8.602288e-11, -8.575824e-11, -8.608631e-11, -8.59189e-11, 
    -8.620575e-11, -8.594759e-11, -8.639479e-11, -8.649217e-11, 
    -8.642562e-11, -8.668123e-11, -8.593328e-11, -8.622052e-11, 
    -8.406023e-11, -8.407294e-11, -8.413214e-11, -8.387192e-11, -8.3856e-11, 
    -8.361752e-11, -8.382971e-11, -8.392008e-11, -8.414945e-11, 
    -8.428513e-11, -8.441411e-11, -8.469769e-11, -8.50144e-11, -8.545725e-11, 
    -8.577539e-11, -8.598866e-11, -8.585788e-11, -8.597334e-11, 
    -8.584428e-11, -8.578378e-11, -8.645568e-11, -8.60784e-11, -8.664447e-11, 
    -8.661314e-11, -8.635697e-11, -8.661667e-11, -8.408186e-11, 
    -8.400874e-11, -8.375486e-11, -8.395354e-11, -8.359155e-11, 
    -8.379418e-11, -8.391069e-11, -8.436023e-11, -8.4459e-11, -8.455058e-11, 
    -8.473146e-11, -8.496359e-11, -8.537081e-11, -8.572511e-11, 
    -8.604854e-11, -8.602484e-11, -8.603318e-11, -8.610544e-11, 
    -8.592646e-11, -8.613482e-11, -8.616979e-11, -8.607835e-11, 
    -8.660895e-11, -8.645736e-11, -8.661247e-11, -8.651378e-11, -8.40325e-11, 
    -8.415554e-11, -8.408906e-11, -8.421409e-11, -8.4126e-11, -8.451766e-11, 
    -8.463508e-11, -8.518453e-11, -8.495903e-11, -8.53179e-11, -8.499548e-11, 
    -8.505261e-11, -8.532962e-11, -8.50129e-11, -8.570558e-11, -8.523598e-11, 
    -8.610825e-11, -8.563932e-11, -8.613763e-11, -8.604713e-11, 
    -8.619696e-11, -8.633115e-11, -8.649996e-11, -8.681145e-11, 
    -8.673932e-11, -8.699982e-11, -8.433897e-11, -8.449856e-11, -8.44845e-11, 
    -8.465151e-11, -8.477503e-11, -8.504272e-11, -8.547207e-11, 
    -8.531062e-11, -8.560702e-11, -8.566653e-11, -8.521622e-11, 
    -8.549271e-11, -8.460536e-11, -8.474874e-11, -8.466337e-11, 
    -8.435156e-11, -8.534783e-11, -8.483655e-11, -8.578065e-11, 
    -8.550368e-11, -8.631202e-11, -8.591002e-11, -8.669962e-11, 
    -8.703718e-11, -8.735484e-11, -8.772611e-11, -8.458565e-11, 
    -8.447721e-11, -8.467137e-11, -8.494001e-11, -8.518923e-11, 
    -8.552058e-11, -8.555447e-11, -8.561656e-11, -8.577734e-11, 
    -8.591253e-11, -8.563619e-11, -8.594642e-11, -8.4782e-11, -8.539221e-11, 
    -8.443622e-11, -8.47241e-11, -8.492416e-11, -8.48364e-11, -8.529216e-11, 
    -8.539958e-11, -8.58361e-11, -8.561044e-11, -8.695387e-11, -8.63595e-11, 
    -8.800877e-11, -8.754788e-11, -8.443933e-11, -8.458528e-11, 
    -8.509322e-11, -8.485154e-11, -8.55427e-11, -8.571282e-11, -8.585111e-11, 
    -8.602791e-11, -8.604699e-11, -8.615174e-11, -8.598009e-11, 
    -8.614495e-11, -8.552128e-11, -8.579999e-11, -8.503516e-11, 
    -8.522132e-11, -8.513568e-11, -8.504174e-11, -8.533166e-11, 
    -8.564054e-11, -8.564713e-11, -8.574617e-11, -8.602529e-11, 
    -8.554549e-11, -8.70306e-11, -8.611346e-11, -8.474442e-11, -8.502556e-11, 
    -8.506569e-11, -8.495679e-11, -8.569576e-11, -8.542801e-11, 
    -8.614919e-11, -8.595427e-11, -8.627363e-11, -8.611493e-11, 
    -8.609159e-11, -8.588777e-11, -8.576088e-11, -8.544029e-11, 
    -8.517944e-11, -8.497258e-11, -8.502068e-11, -8.524791e-11, 
    -8.565943e-11, -8.604872e-11, -8.596344e-11, -8.624935e-11, 
    -8.549258e-11, -8.580991e-11, -8.568727e-11, -8.600706e-11, 
    -8.530633e-11, -8.590308e-11, -8.51538e-11, -8.521949e-11, -8.54227e-11, 
    -8.583145e-11, -8.592186e-11, -8.601842e-11, -8.595884e-11, 
    -8.566987e-11, -8.562253e-11, -8.541776e-11, -8.536123e-11, 
    -8.520519e-11, -8.507601e-11, -8.519404e-11, -8.531799e-11, 
    -8.566999e-11, -8.598721e-11, -8.633307e-11, -8.64177e-11, -8.682181e-11, 
    -8.649286e-11, -8.703572e-11, -8.657421e-11, -8.737309e-11, 
    -8.593765e-11, -8.656062e-11, -8.543194e-11, -8.555354e-11, 
    -8.577347e-11, -8.627789e-11, -8.600556e-11, -8.632405e-11, 
    -8.562067e-11, -8.525575e-11, -8.516132e-11, -8.498516e-11, 
    -8.516535e-11, -8.51507e-11, -8.532312e-11, -8.526771e-11, -8.568168e-11, 
    -8.545931e-11, -8.6091e-11, -8.632153e-11, -8.697252e-11, -8.73716e-11, 
    -8.777782e-11, -8.795716e-11, -8.801175e-11, -8.803457e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.016046e-12, -2.024917e-12, -2.023193e-12, -2.030347e-12, -2.026378e-12, 
    -2.031063e-12, -2.017845e-12, -2.025269e-12, -2.02053e-12, -2.016845e-12, 
    -2.044232e-12, -2.030666e-12, -2.058323e-12, -2.049671e-12, 
    -2.071404e-12, -2.056977e-12, -2.074313e-12, -2.070987e-12, 
    -2.080995e-12, -2.078128e-12, -2.09093e-12, -2.082319e-12, -2.097565e-12, 
    -2.088873e-12, -2.090233e-12, -2.082035e-12, -2.033396e-12, 
    -2.042544e-12, -2.032854e-12, -2.034159e-12, -2.033573e-12, -2.02646e-12, 
    -2.022876e-12, -2.015368e-12, -2.016731e-12, -2.022245e-12, 
    -2.034745e-12, -2.030502e-12, -2.041196e-12, -2.040954e-12, 
    -2.052859e-12, -2.047492e-12, -2.067501e-12, -2.061814e-12, 
    -2.078248e-12, -2.074115e-12, -2.078054e-12, -2.07686e-12, -2.078069e-12, 
    -2.072008e-12, -2.074605e-12, -2.069271e-12, -2.048497e-12, 
    -2.054603e-12, -2.036393e-12, -2.025444e-12, -2.018171e-12, -2.01301e-12, 
    -2.013739e-12, -2.01513e-12, -2.022278e-12, -2.028998e-12, -2.034119e-12, 
    -2.037544e-12, -2.04092e-12, -2.051137e-12, -2.056544e-12, -2.068651e-12, 
    -2.066466e-12, -2.070168e-12, -2.073704e-12, -2.079641e-12, 
    -2.078664e-12, -2.081279e-12, -2.07007e-12, -2.07752e-12, -2.065221e-12, 
    -2.068585e-12, -2.041838e-12, -2.031647e-12, -2.027316e-12, 
    -2.023524e-12, -2.0143e-12, -2.02067e-12, -2.018159e-12, -2.024133e-12, 
    -2.027929e-12, -2.026051e-12, -2.037638e-12, -2.033133e-12, 
    -2.056864e-12, -2.046643e-12, -2.073291e-12, -2.066915e-12, -2.07482e-12, 
    -2.070786e-12, -2.077698e-12, -2.071477e-12, -2.082253e-12, 
    -2.084599e-12, -2.082996e-12, -2.089155e-12, -2.071132e-12, 
    -2.078054e-12, -2.025999e-12, -2.026305e-12, -2.027731e-12, 
    -2.021461e-12, -2.021078e-12, -2.015331e-12, -2.020444e-12, 
    -2.022621e-12, -2.028149e-12, -2.031418e-12, -2.034526e-12, 
    -2.041359e-12, -2.048991e-12, -2.059662e-12, -2.067328e-12, 
    -2.072467e-12, -2.069316e-12, -2.072098e-12, -2.068988e-12, -2.06753e-12, 
    -2.08372e-12, -2.074629e-12, -2.088269e-12, -2.087514e-12, -2.081342e-12, 
    -2.087599e-12, -2.02652e-12, -2.024758e-12, -2.01864e-12, -2.023428e-12, 
    -2.014705e-12, -2.019588e-12, -2.022395e-12, -2.033228e-12, 
    -2.035607e-12, -2.037814e-12, -2.042173e-12, -2.047766e-12, 
    -2.057579e-12, -2.066116e-12, -2.07391e-12, -2.073338e-12, -2.073539e-12, 
    -2.075281e-12, -2.070968e-12, -2.075989e-12, -2.076831e-12, 
    -2.074628e-12, -2.087413e-12, -2.083761e-12, -2.087498e-12, -2.08512e-12, 
    -2.025331e-12, -2.028296e-12, -2.026693e-12, -2.029706e-12, 
    -2.027584e-12, -2.037021e-12, -2.03985e-12, -2.05309e-12, -2.047656e-12, 
    -2.056304e-12, -2.048535e-12, -2.049911e-12, -2.056586e-12, 
    -2.048955e-12, -2.065646e-12, -2.05433e-12, -2.075348e-12, -2.064049e-12, 
    -2.076056e-12, -2.073876e-12, -2.077486e-12, -2.080719e-12, 
    -2.084787e-12, -2.092293e-12, -2.090555e-12, -2.096832e-12, 
    -2.032715e-12, -2.036561e-12, -2.036222e-12, -2.040246e-12, 
    -2.043223e-12, -2.049673e-12, -2.060019e-12, -2.056128e-12, 
    -2.063271e-12, -2.064705e-12, -2.053854e-12, -2.060516e-12, 
    -2.039134e-12, -2.042589e-12, -2.040532e-12, -2.033019e-12, 
    -2.057025e-12, -2.044705e-12, -2.067455e-12, -2.060781e-12, 
    -2.080258e-12, -2.070572e-12, -2.089598e-12, -2.097732e-12, 
    -2.105387e-12, -2.114333e-12, -2.038659e-12, -2.036046e-12, 
    -2.040725e-12, -2.047198e-12, -2.053204e-12, -2.061188e-12, 
    -2.062005e-12, -2.0635e-12, -2.067375e-12, -2.070632e-12, -2.063974e-12, 
    -2.071449e-12, -2.043391e-12, -2.058095e-12, -2.035059e-12, 
    -2.041996e-12, -2.046816e-12, -2.044702e-12, -2.055684e-12, 
    -2.058272e-12, -2.068791e-12, -2.063353e-12, -2.095725e-12, 
    -2.081403e-12, -2.121144e-12, -2.110038e-12, -2.035134e-12, -2.03865e-12, 
    -2.05089e-12, -2.045067e-12, -2.061721e-12, -2.06582e-12, -2.069152e-12, 
    -2.073412e-12, -2.073872e-12, -2.076396e-12, -2.07226e-12, -2.076233e-12, 
    -2.061205e-12, -2.06792e-12, -2.049491e-12, -2.053977e-12, -2.051913e-12, 
    -2.04965e-12, -2.056635e-12, -2.064079e-12, -2.064237e-12, -2.066624e-12, 
    -2.07335e-12, -2.061788e-12, -2.097574e-12, -2.075474e-12, -2.042485e-12, 
    -2.049259e-12, -2.050227e-12, -2.047603e-12, -2.065409e-12, 
    -2.058957e-12, -2.076335e-12, -2.071638e-12, -2.079333e-12, 
    -2.075509e-12, -2.074947e-12, -2.070036e-12, -2.066978e-12, 
    -2.059253e-12, -2.052968e-12, -2.047983e-12, -2.049142e-12, 
    -2.054618e-12, -2.064534e-12, -2.073914e-12, -2.071859e-12, 
    -2.078749e-12, -2.060513e-12, -2.06816e-12, -2.065205e-12, -2.07291e-12, 
    -2.056025e-12, -2.070405e-12, -2.05235e-12, -2.053933e-12, -2.058829e-12, 
    -2.068679e-12, -2.070857e-12, -2.073184e-12, -2.071748e-12, 
    -2.064785e-12, -2.063644e-12, -2.05871e-12, -2.057348e-12, -2.053588e-12, 
    -2.050475e-12, -2.053319e-12, -2.056306e-12, -2.064788e-12, 
    -2.072432e-12, -2.080766e-12, -2.082805e-12, -2.092543e-12, 
    -2.084616e-12, -2.097697e-12, -2.086576e-12, -2.105826e-12, 
    -2.071237e-12, -2.086249e-12, -2.059052e-12, -2.061982e-12, 
    -2.067281e-12, -2.079436e-12, -2.072874e-12, -2.080548e-12, -2.0636e-12, 
    -2.054806e-12, -2.052531e-12, -2.048286e-12, -2.052628e-12, 
    -2.052275e-12, -2.05643e-12, -2.055095e-12, -2.06507e-12, -2.059712e-12, 
    -2.074933e-12, -2.080488e-12, -2.096174e-12, -2.10579e-12, -2.115579e-12, 
    -2.1199e-12, -2.121215e-12, -2.121765e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.36288e-15, 3.371994e-15, 3.370224e-15, 3.377568e-15, 3.373496e-15, 
    3.378303e-15, 3.36473e-15, 3.372355e-15, 3.367489e-15, 3.363703e-15, 
    3.391799e-15, 3.377896e-15, 3.40623e-15, 3.397378e-15, 3.419599e-15, 
    3.404851e-15, 3.422571e-15, 3.419177e-15, 3.429395e-15, 3.426469e-15, 
    3.439517e-15, 3.430745e-15, 3.446279e-15, 3.437425e-15, 3.43881e-15, 
    3.430455e-15, 3.380698e-15, 3.390068e-15, 3.380142e-15, 3.381479e-15, 
    3.38088e-15, 3.373579e-15, 3.369895e-15, 3.362185e-15, 3.363586e-15, 
    3.36925e-15, 3.38208e-15, 3.377729e-15, 3.388697e-15, 3.38845e-15, 
    3.400643e-15, 3.395148e-15, 3.415616e-15, 3.409805e-15, 3.426591e-15, 
    3.422372e-15, 3.426392e-15, 3.425174e-15, 3.426408e-15, 3.42022e-15, 
    3.422872e-15, 3.417425e-15, 3.396176e-15, 3.402426e-15, 3.383771e-15, 
    3.37253e-15, 3.365064e-15, 3.35976e-15, 3.36051e-15, 3.361939e-15, 
    3.369283e-15, 3.376185e-15, 3.38144e-15, 3.384954e-15, 3.388414e-15, 
    3.398873e-15, 3.40441e-15, 3.416789e-15, 3.414559e-15, 3.418339e-15, 
    3.421952e-15, 3.428012e-15, 3.427015e-15, 3.429683e-15, 3.418241e-15, 
    3.425846e-15, 3.413289e-15, 3.416724e-15, 3.389344e-15, 3.378904e-15, 
    3.374453e-15, 3.370564e-15, 3.361086e-15, 3.367632e-15, 3.365052e-15, 
    3.371191e-15, 3.375088e-15, 3.373161e-15, 3.38505e-15, 3.380429e-15, 
    3.404738e-15, 3.394276e-15, 3.421531e-15, 3.415017e-15, 3.423092e-15, 
    3.418973e-15, 3.426028e-15, 3.419679e-15, 3.430677e-15, 3.433068e-15, 
    3.431434e-15, 3.437715e-15, 3.419326e-15, 3.426391e-15, 3.373106e-15, 
    3.373421e-15, 3.374886e-15, 3.368444e-15, 3.368051e-15, 3.362147e-15, 
    3.367401e-15, 3.369637e-15, 3.375314e-15, 3.378669e-15, 3.381857e-15, 
    3.388864e-15, 3.39668e-15, 3.407601e-15, 3.415439e-15, 3.420689e-15, 
    3.417471e-15, 3.420312e-15, 3.417135e-15, 3.415647e-15, 3.432172e-15, 
    3.422896e-15, 3.436811e-15, 3.436043e-15, 3.429746e-15, 3.436129e-15, 
    3.373641e-15, 3.371833e-15, 3.365547e-15, 3.370467e-15, 3.361503e-15, 
    3.36652e-15, 3.369403e-15, 3.380523e-15, 3.382967e-15, 3.38523e-15, 
    3.389698e-15, 3.395429e-15, 3.405471e-15, 3.414199e-15, 3.422163e-15, 
    3.42158e-15, 3.421785e-15, 3.423562e-15, 3.419158e-15, 3.424285e-15, 
    3.425144e-15, 3.422896e-15, 3.435939e-15, 3.432215e-15, 3.436026e-15, 
    3.433602e-15, 3.372421e-15, 3.375464e-15, 3.37382e-15, 3.376911e-15, 
    3.374733e-15, 3.384414e-15, 3.387314e-15, 3.400876e-15, 3.395315e-15, 
    3.404166e-15, 3.396216e-15, 3.397624e-15, 3.40445e-15, 3.396646e-15, 
    3.413718e-15, 3.402143e-15, 3.423631e-15, 3.412083e-15, 3.424354e-15, 
    3.422128e-15, 3.425814e-15, 3.429112e-15, 3.433262e-15, 3.44091e-15, 
    3.43914e-15, 3.445534e-15, 3.38e-15, 3.383943e-15, 3.383598e-15, 
    3.387724e-15, 3.390773e-15, 3.397382e-15, 3.407968e-15, 3.40399e-15, 
    3.411295e-15, 3.41276e-15, 3.401662e-15, 3.408476e-15, 3.386582e-15, 
    3.390121e-15, 3.388016e-15, 3.38031e-15, 3.404904e-15, 3.39229e-15, 
    3.415568e-15, 3.408748e-15, 3.428642e-15, 3.418751e-15, 3.438165e-15, 
    3.446445e-15, 3.45424e-15, 3.463329e-15, 3.386096e-15, 3.383418e-15, 
    3.388215e-15, 3.394844e-15, 3.400995e-15, 3.409164e-15, 3.41e-15, 
    3.411529e-15, 3.415488e-15, 3.418816e-15, 3.41201e-15, 3.41965e-15, 
    3.390938e-15, 3.405999e-15, 3.382403e-15, 3.389512e-15, 3.394454e-15, 
    3.392289e-15, 3.403535e-15, 3.406183e-15, 3.416932e-15, 3.411379e-15, 
    3.444401e-15, 3.429806e-15, 3.47025e-15, 3.458966e-15, 3.382481e-15, 
    3.386088e-15, 3.398626e-15, 3.392663e-15, 3.40971e-15, 3.4139e-15, 
    3.417304e-15, 3.421653e-15, 3.422124e-15, 3.4247e-15, 3.420478e-15, 
    3.424534e-15, 3.409181e-15, 3.416045e-15, 3.397196e-15, 3.401787e-15, 
    3.399676e-15, 3.397358e-15, 3.404509e-15, 3.412117e-15, 3.412282e-15, 
    3.414718e-15, 3.421577e-15, 3.409779e-15, 3.446276e-15, 3.423748e-15, 
    3.390019e-15, 3.396954e-15, 3.397948e-15, 3.395262e-15, 3.41348e-15, 
    3.406883e-15, 3.424638e-15, 3.419843e-15, 3.427699e-15, 3.423796e-15, 
    3.423221e-15, 3.418206e-15, 3.415082e-15, 3.407185e-15, 3.400753e-15, 
    3.395652e-15, 3.396839e-15, 3.402442e-15, 3.412583e-15, 3.422166e-15, 
    3.420066e-15, 3.427102e-15, 3.408475e-15, 3.416288e-15, 3.413269e-15, 
    3.421142e-15, 3.403883e-15, 3.418572e-15, 3.400123e-15, 3.401743e-15, 
    3.406752e-15, 3.416815e-15, 3.419045e-15, 3.42142e-15, 3.419955e-15, 
    3.412841e-15, 3.411675e-15, 3.406631e-15, 3.405236e-15, 3.40139e-15, 
    3.398204e-15, 3.401114e-15, 3.40417e-15, 3.412845e-15, 3.420652e-15, 
    3.429159e-15, 3.43124e-15, 3.441158e-15, 3.433081e-15, 3.446401e-15, 
    3.435071e-15, 3.454677e-15, 3.419427e-15, 3.434744e-15, 3.406981e-15, 
    3.409977e-15, 3.415388e-15, 3.427799e-15, 3.421105e-15, 3.428934e-15, 
    3.41163e-15, 3.402633e-15, 3.400308e-15, 3.395962e-15, 3.400408e-15, 
    3.400046e-15, 3.404298e-15, 3.402932e-15, 3.413133e-15, 3.407655e-15, 
    3.423206e-15, 3.428873e-15, 3.444863e-15, 3.454647e-15, 3.4646e-15, 
    3.468989e-15, 3.470325e-15, 3.470883e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.757414e-09, -8.795924e-09, -8.788438e-09, -8.819499e-09, -8.802268e-09, 
    -8.822607e-09, -8.765221e-09, -8.797453e-09, -8.776877e-09, 
    -8.760881e-09, -8.879777e-09, -8.820884e-09, -8.940946e-09, 
    -8.903387e-09, -8.997732e-09, -8.935102e-09, -9.010361e-09, 
    -8.995925e-09, -9.039372e-09, -9.026925e-09, -9.082499e-09, 
    -9.045117e-09, -9.111305e-09, -9.073571e-09, -9.079475e-09, 
    -9.043884e-09, -8.832735e-09, -8.872445e-09, -8.830383e-09, 
    -8.836045e-09, -8.833504e-09, -8.802624e-09, -8.787064e-09, 
    -8.754471e-09, -8.760388e-09, -8.784326e-09, -8.838591e-09, -8.82017e-09, 
    -8.866594e-09, -8.865546e-09, -8.917229e-09, -8.893926e-09, 
    -8.980791e-09, -8.956103e-09, -9.027445e-09, -9.009503e-09, 
    -9.026603e-09, -9.021417e-09, -9.02667e-09, -9.000356e-09, -9.011631e-09, 
    -8.988476e-09, -8.89829e-09, -8.924796e-09, -8.845744e-09, -8.79821e-09, 
    -8.766635e-09, -8.74423e-09, -8.747398e-09, -8.753436e-09, -8.784466e-09, 
    -8.813639e-09, -8.835871e-09, -8.850742e-09, -8.865395e-09, -8.90975e-09, 
    -8.933224e-09, -8.985784e-09, -8.976298e-09, -8.992368e-09, 
    -9.007718e-09, -9.033492e-09, -9.029249e-09, -9.040606e-09, 
    -8.991943e-09, -9.024284e-09, -8.970894e-09, -8.985497e-09, 
    -8.869382e-09, -8.82514e-09, -8.806338e-09, -8.789877e-09, -8.749834e-09, 
    -8.777487e-09, -8.766586e-09, -8.79252e-09, -8.808999e-09, -8.800848e-09, 
    -8.851148e-09, -8.831593e-09, -8.934615e-09, -8.890241e-09, 
    -9.005928e-09, -8.978245e-09, -9.012563e-09, -8.995051e-09, 
    -9.025057e-09, -8.998052e-09, -9.044831e-09, -9.055017e-09, 
    -9.048057e-09, -9.074795e-09, -8.996555e-09, -9.026603e-09, -8.80062e-09, 
    -8.801949e-09, -8.808142e-09, -8.780921e-09, -8.779256e-09, 
    -8.754308e-09, -8.776506e-09, -8.785959e-09, -8.809954e-09, 
    -8.824147e-09, -8.837639e-09, -8.867303e-09, -8.900433e-09, 
    -8.946759e-09, -8.980039e-09, -9.002348e-09, -8.988668e-09, 
    -9.000745e-09, -8.987245e-09, -8.980916e-09, -9.051201e-09, 
    -9.011735e-09, -9.070949e-09, -9.067673e-09, -9.040876e-09, 
    -9.068041e-09, -8.802883e-09, -8.795233e-09, -8.768676e-09, 
    -8.789459e-09, -8.751592e-09, -8.772789e-09, -8.784977e-09, 
    -8.832003e-09, -8.842334e-09, -8.851915e-09, -8.870836e-09, 
    -8.895118e-09, -8.937716e-09, -8.974778e-09, -9.008612e-09, 
    -9.006132e-09, -9.007005e-09, -9.014563e-09, -8.995841e-09, 
    -9.017637e-09, -9.021296e-09, -9.011731e-09, -9.067234e-09, 
    -9.051377e-09, -9.067603e-09, -9.057278e-09, -8.79772e-09, -8.81059e-09, 
    -8.803636e-09, -8.816714e-09, -8.807501e-09, -8.84847e-09, -8.860754e-09, 
    -8.91823e-09, -8.894641e-09, -8.932182e-09, -8.898454e-09, -8.904431e-09, 
    -8.933408e-09, -8.900276e-09, -8.972736e-09, -8.923612e-09, 
    -9.014857e-09, -8.965804e-09, -9.017931e-09, -9.008465e-09, 
    -9.024138e-09, -9.038175e-09, -9.055833e-09, -9.088417e-09, 
    -9.080871e-09, -9.10812e-09, -8.829778e-09, -8.846473e-09, -8.845002e-09, 
    -8.862473e-09, -8.875393e-09, -8.903396e-09, -8.94831e-09, -8.93142e-09, 
    -8.962426e-09, -8.968651e-09, -8.921545e-09, -8.950468e-09, 
    -8.857645e-09, -8.872643e-09, -8.863712e-09, -8.831096e-09, 
    -8.935314e-09, -8.881829e-09, -8.98059e-09, -8.951616e-09, -9.036174e-09, 
    -8.994122e-09, -9.076718e-09, -9.112028e-09, -9.145258e-09, 
    -9.184094e-09, -8.855583e-09, -8.84424e-09, -8.86455e-09, -8.892651e-09, 
    -8.918723e-09, -8.953384e-09, -8.956929e-09, -8.963423e-09, 
    -8.980242e-09, -8.994384e-09, -8.965477e-09, -8.997929e-09, 
    -8.876123e-09, -8.939955e-09, -8.839952e-09, -8.870066e-09, 
    -8.890995e-09, -8.881814e-09, -8.92949e-09, -8.940726e-09, -8.986389e-09, 
    -8.962784e-09, -9.103315e-09, -9.04114e-09, -9.213662e-09, -9.165451e-09, 
    -8.840277e-09, -8.855544e-09, -8.908679e-09, -8.883398e-09, 
    -8.955698e-09, -8.973494e-09, -8.98796e-09, -9.006453e-09, -9.008449e-09, 
    -9.019407e-09, -9.001451e-09, -9.018698e-09, -8.953458e-09, 
    -8.982612e-09, -8.902605e-09, -8.922079e-09, -8.91312e-09, -8.903293e-09, 
    -8.933621e-09, -8.965932e-09, -8.966621e-09, -8.976982e-09, -9.00618e-09, 
    -8.95599e-09, -9.111341e-09, -9.015403e-09, -8.872192e-09, -8.9016e-09, 
    -8.9058e-09, -8.894408e-09, -8.97171e-09, -8.943701e-09, -9.019139e-09, 
    -8.998751e-09, -9.032157e-09, -9.015557e-09, -9.013115e-09, 
    -8.991794e-09, -8.97852e-09, -8.944985e-09, -8.917699e-09, -8.89606e-09, 
    -8.901091e-09, -8.924861e-09, -8.967908e-09, -9.008631e-09, -8.99971e-09, 
    -9.029618e-09, -8.950455e-09, -8.98365e-09, -8.970821e-09, -9.004273e-09, 
    -8.930972e-09, -8.993395e-09, -8.915016e-09, -8.921888e-09, 
    -8.943145e-09, -8.985903e-09, -8.995361e-09, -9.005461e-09, 
    -8.999228e-09, -8.969001e-09, -8.964048e-09, -8.942628e-09, 
    -8.936714e-09, -8.920392e-09, -8.906879e-09, -8.919225e-09, 
    -8.932191e-09, -8.969013e-09, -9.002196e-09, -9.038374e-09, 
    -9.047228e-09, -9.089501e-09, -9.05509e-09, -9.111876e-09, -9.063601e-09, 
    -9.147167e-09, -8.997011e-09, -9.062178e-09, -8.944111e-09, 
    -8.956831e-09, -8.979838e-09, -9.032603e-09, -9.004116e-09, 
    -9.037431e-09, -8.963855e-09, -8.925682e-09, -8.915803e-09, 
    -8.897375e-09, -8.916224e-09, -8.914691e-09, -8.932727e-09, 
    -8.926931e-09, -8.970236e-09, -8.946975e-09, -9.013053e-09, 
    -9.037167e-09, -9.105265e-09, -9.147011e-09, -9.189503e-09, 
    -9.208263e-09, -9.213973e-09, -9.21636e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039165e-10, -1.043737e-10, -1.042848e-10, -1.046535e-10, -1.04449e-10, 
    -1.046904e-10, -1.040092e-10, -1.043918e-10, -1.041476e-10, 
    -1.039577e-10, -1.053691e-10, -1.046699e-10, -1.060952e-10, 
    -1.056493e-10, -1.067693e-10, -1.060258e-10, -1.069192e-10, 
    -1.067479e-10, -1.072636e-10, -1.071159e-10, -1.077756e-10, 
    -1.073318e-10, -1.081176e-10, -1.076696e-10, -1.077397e-10, 
    -1.073172e-10, -1.048106e-10, -1.05282e-10, -1.047827e-10, -1.048499e-10, 
    -1.048198e-10, -1.044532e-10, -1.042685e-10, -1.038816e-10, 
    -1.039518e-10, -1.04236e-10, -1.048801e-10, -1.046615e-10, -1.052126e-10, 
    -1.052001e-10, -1.058136e-10, -1.05537e-10, -1.065682e-10, -1.062751e-10, 
    -1.07122e-10, -1.069091e-10, -1.07112e-10, -1.070505e-10, -1.071128e-10, 
    -1.068005e-10, -1.069343e-10, -1.066594e-10, -1.055888e-10, 
    -1.059035e-10, -1.04965e-10, -1.044008e-10, -1.04026e-10, -1.0376e-10, 
    -1.037976e-10, -1.038693e-10, -1.042376e-10, -1.045839e-10, 
    -1.048478e-10, -1.050244e-10, -1.051983e-10, -1.057249e-10, 
    -1.060035e-10, -1.066275e-10, -1.065149e-10, -1.067056e-10, 
    -1.068879e-10, -1.071938e-10, -1.071435e-10, -1.072783e-10, 
    -1.067006e-10, -1.070845e-10, -1.064507e-10, -1.066241e-10, 
    -1.052457e-10, -1.047205e-10, -1.044973e-10, -1.043019e-10, 
    -1.038265e-10, -1.041548e-10, -1.040254e-10, -1.043332e-10, 
    -1.045289e-10, -1.044321e-10, -1.050292e-10, -1.047971e-10, -1.0602e-10, 
    -1.054933e-10, -1.068666e-10, -1.06538e-10, -1.069454e-10, -1.067375e-10, 
    -1.070937e-10, -1.067731e-10, -1.073285e-10, -1.074494e-10, 
    -1.073667e-10, -1.076842e-10, -1.067553e-10, -1.07112e-10, -1.044294e-10, 
    -1.044452e-10, -1.045187e-10, -1.041956e-10, -1.041758e-10, 
    -1.038797e-10, -1.041432e-10, -1.042554e-10, -1.045402e-10, 
    -1.047087e-10, -1.048688e-10, -1.05221e-10, -1.056143e-10, -1.061642e-10, 
    -1.065593e-10, -1.068241e-10, -1.066617e-10, -1.068051e-10, 
    -1.066448e-10, -1.065697e-10, -1.074041e-10, -1.069356e-10, 
    -1.076385e-10, -1.075996e-10, -1.072815e-10, -1.07604e-10, -1.044563e-10, 
    -1.043655e-10, -1.040502e-10, -1.042969e-10, -1.038474e-10, -1.04099e-10, 
    -1.042437e-10, -1.048019e-10, -1.049246e-10, -1.050383e-10, 
    -1.052629e-10, -1.055512e-10, -1.060569e-10, -1.064968e-10, 
    -1.068985e-10, -1.06869e-10, -1.068794e-10, -1.069691e-10, -1.067469e-10, 
    -1.070056e-10, -1.070491e-10, -1.069355e-10, -1.075944e-10, 
    -1.074062e-10, -1.075988e-10, -1.074762e-10, -1.04395e-10, -1.045478e-10, 
    -1.044652e-10, -1.046204e-10, -1.045111e-10, -1.049974e-10, 
    -1.051432e-10, -1.058255e-10, -1.055455e-10, -1.059912e-10, 
    -1.055908e-10, -1.056617e-10, -1.060057e-10, -1.056124e-10, 
    -1.064726e-10, -1.058894e-10, -1.069726e-10, -1.063903e-10, 
    -1.070091e-10, -1.068967e-10, -1.070828e-10, -1.072494e-10, 
    -1.074591e-10, -1.078459e-10, -1.077563e-10, -1.080798e-10, 
    -1.047755e-10, -1.049737e-10, -1.049562e-10, -1.051636e-10, -1.05317e-10, 
    -1.056494e-10, -1.061826e-10, -1.059821e-10, -1.063502e-10, 
    -1.064241e-10, -1.058649e-10, -1.062082e-10, -1.051063e-10, 
    -1.052844e-10, -1.051784e-10, -1.047912e-10, -1.060283e-10, 
    -1.053934e-10, -1.065658e-10, -1.062219e-10, -1.072257e-10, 
    -1.067265e-10, -1.07707e-10, -1.081262e-10, -1.085207e-10, -1.089817e-10, 
    -1.050819e-10, -1.049472e-10, -1.051883e-10, -1.055219e-10, 
    -1.058314e-10, -1.062428e-10, -1.062849e-10, -1.06362e-10, -1.065617e-10, 
    -1.067296e-10, -1.063864e-10, -1.067717e-10, -1.053257e-10, 
    -1.060834e-10, -1.048963e-10, -1.052538e-10, -1.055022e-10, 
    -1.053932e-10, -1.059592e-10, -1.060926e-10, -1.066347e-10, 
    -1.063544e-10, -1.080227e-10, -1.072846e-10, -1.093328e-10, 
    -1.087604e-10, -1.049002e-10, -1.050814e-10, -1.057122e-10, -1.05412e-10, 
    -1.062703e-10, -1.064816e-10, -1.066533e-10, -1.068729e-10, 
    -1.068965e-10, -1.070266e-10, -1.068135e-10, -1.070182e-10, 
    -1.062437e-10, -1.065898e-10, -1.0564e-10, -1.058712e-10, -1.057649e-10, 
    -1.056482e-10, -1.060082e-10, -1.063918e-10, -1.064e-10, -1.06523e-10, 
    -1.068696e-10, -1.062738e-10, -1.08118e-10, -1.069791e-10, -1.05279e-10, 
    -1.056281e-10, -1.05678e-10, -1.055427e-10, -1.064604e-10, -1.061279e-10, 
    -1.070235e-10, -1.067814e-10, -1.07178e-10, -1.069809e-10, -1.069519e-10, 
    -1.066988e-10, -1.065412e-10, -1.061431e-10, -1.058192e-10, 
    -1.055624e-10, -1.056221e-10, -1.059042e-10, -1.064153e-10, 
    -1.068987e-10, -1.067928e-10, -1.071479e-10, -1.062081e-10, 
    -1.066022e-10, -1.064498e-10, -1.06847e-10, -1.059768e-10, -1.067178e-10, 
    -1.057874e-10, -1.05869e-10, -1.061213e-10, -1.066289e-10, -1.067412e-10, 
    -1.068611e-10, -1.067871e-10, -1.064282e-10, -1.063694e-10, 
    -1.061152e-10, -1.06045e-10, -1.058512e-10, -1.056908e-10, -1.058373e-10, 
    -1.059913e-10, -1.064284e-10, -1.068223e-10, -1.072518e-10, 
    -1.073569e-10, -1.078588e-10, -1.074502e-10, -1.081244e-10, 
    -1.075513e-10, -1.085433e-10, -1.067608e-10, -1.075344e-10, 
    -1.061328e-10, -1.062838e-10, -1.065569e-10, -1.071833e-10, 
    -1.068451e-10, -1.072406e-10, -1.063671e-10, -1.05914e-10, -1.057967e-10, 
    -1.05578e-10, -1.058017e-10, -1.057835e-10, -1.059976e-10, -1.059288e-10, 
    -1.064429e-10, -1.061668e-10, -1.069512e-10, -1.072375e-10, 
    -1.080459e-10, -1.085415e-10, -1.09046e-10, -1.092687e-10, -1.093365e-10, 
    -1.093648e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.619386e-12, -8.657319e-12, -8.649944e-12, -8.680541e-12, -8.663568e-12, 
    -8.683602e-12, -8.627076e-12, -8.658825e-12, -8.638557e-12, -8.6228e-12, 
    -8.739918e-12, -8.681905e-12, -8.800172e-12, -8.763176e-12, 
    -8.856112e-12, -8.794416e-12, -8.868552e-12, -8.854331e-12, -8.89713e-12, 
    -8.884869e-12, -8.939613e-12, -8.902789e-12, -8.96799e-12, -8.930819e-12, 
    -8.936634e-12, -8.901574e-12, -8.693579e-12, -8.732696e-12, 
    -8.691262e-12, -8.696839e-12, -8.694337e-12, -8.663919e-12, 
    -8.648591e-12, -8.616485e-12, -8.622314e-12, -8.645894e-12, 
    -8.699348e-12, -8.681202e-12, -8.726932e-12, -8.725899e-12, -8.77681e-12, 
    -8.753855e-12, -8.839423e-12, -8.815103e-12, -8.88538e-12, -8.867707e-12, 
    -8.88455e-12, -8.879443e-12, -8.884617e-12, -8.858696e-12, -8.869802e-12, 
    -8.846993e-12, -8.758155e-12, -8.784264e-12, -8.706393e-12, -8.65957e-12, 
    -8.628469e-12, -8.606399e-12, -8.609518e-12, -8.615467e-12, 
    -8.646032e-12, -8.674768e-12, -8.696668e-12, -8.711317e-12, 
    -8.725751e-12, -8.769443e-12, -8.792566e-12, -8.844342e-12, 
    -8.834997e-12, -8.850827e-12, -8.865949e-12, -8.891337e-12, 
    -8.887158e-12, -8.898345e-12, -8.850408e-12, -8.882267e-12, 
    -8.829675e-12, -8.844059e-12, -8.729678e-12, -8.686097e-12, 
    -8.667576e-12, -8.651362e-12, -8.611918e-12, -8.639157e-12, 
    -8.628419e-12, -8.653965e-12, -8.670197e-12, -8.662169e-12, 
    -8.711717e-12, -8.692455e-12, -8.793937e-12, -8.750225e-12, 
    -8.864185e-12, -8.836915e-12, -8.870721e-12, -8.85347e-12, -8.883028e-12, 
    -8.856426e-12, -8.902507e-12, -8.912542e-12, -8.905684e-12, 
    -8.932024e-12, -8.854951e-12, -8.884551e-12, -8.661944e-12, 
    -8.663253e-12, -8.669353e-12, -8.64254e-12, -8.6409e-12, -8.616326e-12, 
    -8.638191e-12, -8.647502e-12, -8.671138e-12, -8.685119e-12, -8.69841e-12, 
    -8.727631e-12, -8.760266e-12, -8.8059e-12, -8.838682e-12, -8.860658e-12, 
    -8.847183e-12, -8.859079e-12, -8.84578e-12, -8.839547e-12, -8.908782e-12, 
    -8.869906e-12, -8.928236e-12, -8.925007e-12, -8.89861e-12, -8.925372e-12, 
    -8.664173e-12, -8.656638e-12, -8.630477e-12, -8.650951e-12, -8.61365e-12, 
    -8.63453e-12, -8.646535e-12, -8.692858e-12, -8.703035e-12, -8.712472e-12, 
    -8.73111e-12, -8.755031e-12, -8.796992e-12, -8.8335e-12, -8.866828e-12, 
    -8.864386e-12, -8.865245e-12, -8.872692e-12, -8.854249e-12, 
    -8.875719e-12, -8.879323e-12, -8.8699e-12, -8.924575e-12, -8.908955e-12, 
    -8.924939e-12, -8.914768e-12, -8.659087e-12, -8.671766e-12, 
    -8.664915e-12, -8.677798e-12, -8.668722e-12, -8.709079e-12, 
    -8.721179e-12, -8.777796e-12, -8.75456e-12, -8.79154e-12, -8.758316e-12, 
    -8.764203e-12, -8.792748e-12, -8.760112e-12, -8.831488e-12, 
    -8.783098e-12, -8.87298e-12, -8.82466e-12, -8.876008e-12, -8.866683e-12, 
    -8.882122e-12, -8.89595e-12, -8.913345e-12, -8.945442e-12, -8.93801e-12, 
    -8.964852e-12, -8.690666e-12, -8.707111e-12, -8.705663e-12, 
    -8.722872e-12, -8.7356e-12, -8.763185e-12, -8.807427e-12, -8.79079e-12, 
    -8.821333e-12, -8.827464e-12, -8.781062e-12, -8.809553e-12, 
    -8.718117e-12, -8.73289e-12, -8.724093e-12, -8.691964e-12, -8.794625e-12, 
    -8.741939e-12, -8.839224e-12, -8.810684e-12, -8.893978e-12, 
    -8.852555e-12, -8.933919e-12, -8.968703e-12, -9.001436e-12, 
    -9.039693e-12, -8.716086e-12, -8.704912e-12, -8.724918e-12, -8.7526e-12, 
    -8.778282e-12, -8.812425e-12, -8.815918e-12, -8.822314e-12, 
    -8.838882e-12, -8.852813e-12, -8.824338e-12, -8.856305e-12, 
    -8.736318e-12, -8.799197e-12, -8.700688e-12, -8.730352e-12, 
    -8.750968e-12, -8.741924e-12, -8.788888e-12, -8.799957e-12, 
    -8.844938e-12, -8.821686e-12, -8.960118e-12, -8.898872e-12, 
    -9.068819e-12, -9.021327e-12, -8.701008e-12, -8.716047e-12, 
    -8.768389e-12, -8.743484e-12, -8.814704e-12, -8.832234e-12, 
    -8.846484e-12, -8.864702e-12, -8.866669e-12, -8.877462e-12, 
    -8.859775e-12, -8.876764e-12, -8.812498e-12, -8.841217e-12, 
    -8.762405e-12, -8.781587e-12, -8.772763e-12, -8.763083e-12, 
    -8.792958e-12, -8.824786e-12, -8.825466e-12, -8.835671e-12, 
    -8.864433e-12, -8.814992e-12, -8.968025e-12, -8.873518e-12, 
    -8.732446e-12, -8.761415e-12, -8.765552e-12, -8.75433e-12, -8.830477e-12, 
    -8.802886e-12, -8.877199e-12, -8.857115e-12, -8.890022e-12, -8.87367e-12, 
    -8.871264e-12, -8.850262e-12, -8.837186e-12, -8.804152e-12, 
    -8.777272e-12, -8.755958e-12, -8.760914e-12, -8.784328e-12, 
    -8.826733e-12, -8.866847e-12, -8.85806e-12, -8.887522e-12, -8.80954e-12, 
    -8.842239e-12, -8.829602e-12, -8.862555e-12, -8.790348e-12, 
    -8.851839e-12, -8.77463e-12, -8.781399e-12, -8.802339e-12, -8.844458e-12, 
    -8.853775e-12, -8.863725e-12, -8.857585e-12, -8.827809e-12, -8.82293e-12, 
    -8.80183e-12, -8.796004e-12, -8.779926e-12, -8.766615e-12, -8.778777e-12, 
    -8.791549e-12, -8.827821e-12, -8.860509e-12, -8.896147e-12, 
    -8.904868e-12, -8.94651e-12, -8.912614e-12, -8.968552e-12, -8.920996e-12, 
    -9.003316e-12, -8.855401e-12, -8.919595e-12, -8.803291e-12, -8.81582e-12, 
    -8.838484e-12, -8.890462e-12, -8.8624e-12, -8.895218e-12, -8.822739e-12, 
    -8.785137e-12, -8.775406e-12, -8.757254e-12, -8.775821e-12, -8.77431e-12, 
    -8.792077e-12, -8.786368e-12, -8.829025e-12, -8.806112e-12, 
    -8.871204e-12, -8.894959e-12, -8.962039e-12, -9.003163e-12, 
    -9.045022e-12, -9.063502e-12, -9.069127e-12, -9.071478e-12 ;

 SMIN_NH4 =
  0.0004617845, 0.0004637133, 0.0004633381, 0.0004648938, 0.0004640307, 
    0.0004650494, 0.0004621751, 0.0004637896, 0.0004627588, 0.0004619575, 
    0.0004679122, 0.0004649628, 0.0004709742, 0.0004690938, 0.0004738166, 
    0.0004706816, 0.0004744485, 0.0004737258, 0.0004759001, 0.0004752771, 
    0.0004780583, 0.0004761874, 0.0004794993, 0.0004776113, 0.0004779067, 
    0.0004761255, 0.0004655565, 0.0004675456, 0.0004654386, 0.0004657223, 
    0.0004655949, 0.0004640484, 0.0004632692, 0.0004616363, 0.0004619327, 
    0.0004631318, 0.0004658494, 0.0004649267, 0.0004672513, 0.0004671988, 
    0.0004697865, 0.0004686198, 0.0004729683, 0.0004717323, 0.0004753031, 
    0.0004744051, 0.0004752608, 0.0004750012, 0.000475264, 0.0004739472, 
    0.0004745113, 0.0004733524, 0.000468839, 0.0004701659, 0.0004662078, 
    0.0004638275, 0.0004622457, 0.0004611234, 0.000461282, 0.0004615845, 
    0.0004631387, 0.0004645996, 0.0004657129, 0.0004664575, 0.0004671911, 
    0.0004694124, 0.0004705873, 0.0004732182, 0.0004727432, 0.0004735475, 
    0.0004743157, 0.0004756055, 0.0004753931, 0.0004759614, 0.0004735259, 
    0.0004751446, 0.0004724722, 0.0004732032, 0.0004673919, 0.0004651758, 
    0.0004642345, 0.0004634098, 0.0004614039, 0.0004627892, 0.0004622431, 
    0.0004635418, 0.0004643671, 0.0004639588, 0.0004664778, 0.0004654985, 
    0.0004706568, 0.0004684352, 0.0004742262, 0.0004728405, 0.0004745581, 
    0.0004736816, 0.0004751833, 0.0004738317, 0.0004761727, 0.0004766826, 
    0.000476334, 0.000477672, 0.0004737564, 0.0004752603, 0.0004639477, 
    0.0004640144, 0.0004643244, 0.0004629611, 0.0004628777, 0.0004616279, 
    0.0004627397, 0.0004632132, 0.0004644148, 0.0004651255, 0.0004658011, 
    0.0004672866, 0.0004689455, 0.0004712645, 0.0004729303, 0.0004740467, 
    0.000473362, 0.0004739664, 0.0004732907, 0.0004729738, 0.0004764914, 
    0.0004745164, 0.0004774794, 0.0004773154, 0.0004759745, 0.0004773338, 
    0.000464061, 0.0004636777, 0.0004623476, 0.0004633885, 0.0004614917, 
    0.0004625536, 0.000463164, 0.0004655191, 0.0004660362, 0.000466516, 
    0.0004674633, 0.0004686791, 0.0004708118, 0.0004726669, 0.0004743601, 
    0.000474236, 0.0004742796, 0.0004746579, 0.0004737208, 0.0004748116, 
    0.0004749947, 0.0004745159, 0.0004772933, 0.0004764998, 0.0004773117, 
    0.000476795, 0.0004638022, 0.0004644468, 0.0004640984, 0.0004647534, 
    0.0004642919, 0.0004663437, 0.0004669588, 0.0004698364, 0.0004686552, 
    0.0004705348, 0.000468846, 0.0004691453, 0.0004705962, 0.000468937, 
    0.0004725646, 0.0004701055, 0.0004746725, 0.0004722176, 0.0004748262, 
    0.0004743524, 0.0004751367, 0.0004758392, 0.0004767227, 0.0004783532, 
    0.0004779755, 0.0004793389, 0.0004654076, 0.0004662437, 0.0004661698, 
    0.0004670446, 0.0004676915, 0.0004690936, 0.0004713421, 0.0004704964, 
    0.0004720484, 0.0004723601, 0.0004700018, 0.0004714499, 0.0004668025, 
    0.0004675535, 0.0004671062, 0.0004654728, 0.000470691, 0.0004680133, 
    0.0004729572, 0.0004715068, 0.0004757389, 0.0004736345, 0.0004777677, 
    0.0004795346, 0.0004811966, 0.0004831394, 0.0004666997, 0.0004661315, 
    0.0004671485, 0.0004685558, 0.0004698608, 0.000471596, 0.0004717733, 
    0.0004720983, 0.0004729401, 0.0004736479, 0.0004722011, 0.0004738252, 
    0.000467728, 0.0004709233, 0.0004659162, 0.0004674243, 0.000468472, 
    0.0004680122, 0.000470399, 0.0004709615, 0.0004732472, 0.0004720656, 
    0.0004790986, 0.0004759874, 0.000484618, 0.0004822067, 0.000465933, 
    0.0004666975, 0.000469358, 0.0004680922, 0.0004717115, 0.0004726024, 
    0.0004733263, 0.000474252, 0.0004743517, 0.0004749002, 0.0004740014, 
    0.0004748645, 0.0004715991, 0.0004730583, 0.0004690531, 0.0004700281, 
    0.0004695795, 0.0004690874, 0.0004706056, 0.0004722233, 0.0004722576, 
    0.0004727762, 0.0004742382, 0.0004717252, 0.0004795003, 0.0004746995, 
    0.000467531, 0.0004690036, 0.0004692136, 0.0004686432, 0.0004725129, 
    0.0004711109, 0.0004748868, 0.0004738662, 0.0004755381, 0.0004747073, 
    0.000474585, 0.0004735179, 0.0004728534, 0.0004711748, 0.0004698087, 
    0.0004687253, 0.000468977, 0.0004701672, 0.000472322, 0.0004743602, 
    0.0004739137, 0.0004754103, 0.000471448, 0.0004731097, 0.0004724675, 
    0.0004741417, 0.0004704738, 0.0004735991, 0.0004696749, 0.0004700188, 
    0.0004710829, 0.0004732235, 0.0004736964, 0.0004742021, 0.0004738899, 
    0.0004723771, 0.0004721291, 0.0004710566, 0.0004707606, 0.0004699434, 
    0.0004692668, 0.000469885, 0.000470534, 0.0004723772, 0.0004740381, 
    0.0004758486, 0.0004762915, 0.0004784071, 0.0004766852, 0.0004795268, 
    0.0004771114, 0.000481292, 0.0004737796, 0.0004770409, 0.0004711313, 
    0.0004717679, 0.0004729197, 0.0004755605, 0.0004741345, 0.0004758021, 
    0.0004721193, 0.0004702084, 0.0004697136, 0.0004687911, 0.0004697346, 
    0.0004696579, 0.0004705607, 0.0004702705, 0.0004724382, 0.0004712738, 
    0.0004745813, 0.0004757882, 0.0004791955, 0.0004812839, 0.0004834092, 
    0.0004843474, 0.0004846329, 0.0004847522 ;

 SMIN_NH4_vr =
  0.003023126, 0.003028289, 0.003027279, 0.003031441, 0.003029128, 
    0.003031848, 0.003024156, 0.003028473, 0.003025713, 0.003023563, 
    0.003039481, 0.003031601, 0.003047637, 0.003042621, 0.003055192, 
    0.003046851, 0.003056868, 0.003054941, 0.003060716, 0.003059057, 
    0.003066436, 0.003061471, 0.003070248, 0.003065244, 0.003066024, 
    0.003061292, 0.003033208, 0.003038524, 0.003032887, 0.003033646, 
    0.003033301, 0.003029163, 0.003027078, 0.003022701, 0.003023491, 
    0.003026702, 0.003033965, 0.003031493, 0.003037699, 0.003037559, 
    0.003044455, 0.003041345, 0.003052923, 0.00304963, 0.003059123, 
    0.003056733, 0.003059005, 0.003058311, 0.003059005, 0.003055507, 
    0.003057, 0.003053919, 0.003041965, 0.003045498, 0.003034937, 
    0.003028572, 0.003024333, 0.003021328, 0.003021746, 0.003022557, 
    0.003026715, 0.003030617, 0.003033591, 0.003035575, 0.00303753, 
    0.003043459, 0.003046585, 0.003053582, 0.003052316, 0.003054452, 
    0.003056492, 0.003059914, 0.003059348, 0.003060853, 0.003054378, 
    0.003058681, 0.003051569, 0.003053515, 0.003038101, 0.003032173, 
    0.003029657, 0.003027445, 0.003022071, 0.003025781, 0.003024315, 
    0.003027786, 0.003029992, 0.003028895, 0.003035626, 0.003033005, 
    0.003046765, 0.003040843, 0.003056258, 0.003052569, 0.003057131, 
    0.003054802, 0.003058787, 0.003055195, 0.003061408, 0.003062762, 
    0.003061831, 0.003065381, 0.003054977, 0.003058975, 0.003028883, 
    0.003029062, 0.003029887, 0.003026236, 0.003026012, 0.003022661, 
    0.003025633, 0.003026902, 0.003030111, 0.003032007, 0.003033808, 
    0.003037776, 0.003042198, 0.003048373, 0.003052804, 0.003055768, 
    0.003053946, 0.003055549, 0.003053751, 0.003052903, 0.003062247, 
    0.003057002, 0.003064861, 0.003064427, 0.003060865, 0.003064467, 
    0.003029181, 0.003028151, 0.00302459, 0.003027371, 0.00302229, 
    0.003025134, 0.003026765, 0.003033057, 0.003034434, 0.003035716, 
    0.003038241, 0.00304148, 0.003047164, 0.003052097, 0.003056597, 
    0.003056263, 0.003056378, 0.003057379, 0.003054887, 0.003057781, 
    0.003058264, 0.003056992, 0.00306436, 0.003062255, 0.003064405, 
    0.003063029, 0.00302848, 0.0030302, 0.003029264, 0.003031017, 
    0.003029776, 0.003035261, 0.0030369, 0.003044571, 0.003041417, 
    0.003046428, 0.00304192, 0.003042719, 0.003046584, 0.003042154, 
    0.003051817, 0.003045265, 0.003057414, 0.003050884, 0.003057817, 
    0.003056552, 0.003058632, 0.003060499, 0.003062838, 0.003067164, 
    0.003066156, 0.00306977, 0.003032765, 0.003034994, 0.003034795, 
    0.003037127, 0.00303885, 0.00304259, 0.003048577, 0.00304632, 
    0.003050449, 0.003051279, 0.003044992, 0.003048851, 0.003036456, 
    0.003038457, 0.003037261, 0.003032894, 0.003046815, 0.003039672, 
    0.00305284, 0.003048976, 0.003060224, 0.003054634, 0.003065602, 
    0.003070288, 0.003074682, 0.003079817, 0.003036208, 0.003034686, 
    0.003037398, 0.003041155, 0.003044627, 0.003049249, 0.003049717, 
    0.003050578, 0.003052813, 0.003054696, 0.003050845, 0.003055159, 
    0.003038921, 0.003047433, 0.003034072, 0.003038102, 0.003040889, 
    0.003039663, 0.003046022, 0.003047516, 0.003053596, 0.003050452, 
    0.003069124, 0.003060872, 0.003083715, 0.003077345, 0.003034153, 
    0.00303619, 0.003043285, 0.003039909, 0.003049548, 0.00305192, 
    0.003053838, 0.003056301, 0.003056559, 0.003058017, 0.003055621, 
    0.003057916, 0.003049225, 0.003053109, 0.003042439, 0.003045033, 
    0.003043836, 0.00304252, 0.003046562, 0.003050871, 0.003050957, 
    0.003052333, 0.003056224, 0.003049529, 0.003070181, 0.003057438, 
    0.003038411, 0.003042337, 0.003042891, 0.003041371, 0.003051673, 
    0.003047942, 0.003057981, 0.003055264, 0.003059702, 0.003057496, 
    0.003057165, 0.003054329, 0.003052555, 0.003048089, 0.003044443, 
    0.003041554, 0.003042219, 0.003045393, 0.003051125, 0.003056545, 
    0.003055355, 0.003059326, 0.003048785, 0.003053209, 0.003051494, 
    0.003055946, 0.003046248, 0.003054571, 0.003044115, 0.003045027, 
    0.003047859, 0.003053557, 0.003054806, 0.003056152, 0.003055315, 
    0.003051293, 0.003050629, 0.003047769, 0.003046977, 0.0030448, 
    0.00304299, 0.003044638, 0.003046362, 0.003051269, 0.003055683, 
    0.003060488, 0.003061662, 0.003067273, 0.003062704, 0.003070236, 
    0.003063832, 0.003074902, 0.00305504, 0.003063703, 0.003047987, 
    0.003049678, 0.003052743, 0.003059758, 0.003055963, 0.003060395, 
    0.0030506, 0.003045509, 0.003044185, 0.003041726, 0.003044235, 
    0.003044031, 0.003046433, 0.003045655, 0.003051423, 0.003048324, 
    0.003057116, 0.003060323, 0.003069356, 0.003074882, 0.003080498, 
    0.003082972, 0.003083724, 0.003084036,
  0.001810043, 0.001816795, 0.001815482, 0.001820924, 0.001817906, 
    0.001821468, 0.001811412, 0.001817063, 0.001813456, 0.001810651, 
    0.001831472, 0.001821166, 0.001842153, 0.001835595, 0.001852053, 
    0.001841133, 0.001854252, 0.001851737, 0.001859301, 0.001857135, 
    0.0018668, 0.0018603, 0.001871802, 0.001865248, 0.001866274, 0.001860086, 
    0.001823241, 0.00183019, 0.001822829, 0.00182382, 0.001823375, 
    0.001817968, 0.001815242, 0.001809526, 0.001810564, 0.001814762, 
    0.001824266, 0.001821041, 0.001829164, 0.001828981, 0.001838012, 
    0.001833942, 0.0018491, 0.001844796, 0.001857225, 0.001854102, 
    0.001857079, 0.001856176, 0.00185709, 0.001852509, 0.001854473, 
    0.001850439, 0.001834704, 0.001839334, 0.001825517, 0.001817196, 
    0.00181166, 0.00180773, 0.001808286, 0.001809345, 0.001814787, 
    0.001819897, 0.001823789, 0.001826391, 0.001828954, 0.001836708, 
    0.001840805, 0.001849971, 0.001848317, 0.001851118, 0.001853791, 
    0.001858278, 0.001857539, 0.001859515, 0.001851043, 0.001856676, 
    0.001847375, 0.00184992, 0.001829654, 0.001821911, 0.00181862, 
    0.001815735, 0.001808713, 0.001813563, 0.001811652, 0.001816197, 
    0.001819085, 0.001817657, 0.001826463, 0.001823041, 0.001841048, 
    0.001833298, 0.001853479, 0.001848656, 0.001854635, 0.001851585, 
    0.00185681, 0.001852107, 0.00186025, 0.001862022, 0.001860812, 
    0.00186546, 0.001851847, 0.001857079, 0.001817617, 0.00181785, 
    0.001818934, 0.001814165, 0.001813873, 0.001809498, 0.001813391, 
    0.001815048, 0.001819252, 0.001821737, 0.001824099, 0.001829288, 
    0.001835079, 0.001843167, 0.001848969, 0.001852856, 0.001850473, 
    0.001852577, 0.001850225, 0.001849122, 0.001861359, 0.001854491, 
    0.001864792, 0.001864222, 0.001859563, 0.001864286, 0.001818013, 
    0.001816673, 0.001812018, 0.001815661, 0.001809021, 0.001812739, 
    0.001814876, 0.001823113, 0.00182492, 0.001826597, 0.001829906, 
    0.00183415, 0.001841589, 0.001848052, 0.001853946, 0.001853515, 
    0.001853667, 0.001854983, 0.001851722, 0.001855518, 0.001856155, 
    0.00185449, 0.001864146, 0.001861389, 0.00186421, 0.001862415, 
    0.001817108, 0.001819363, 0.001818145, 0.001820436, 0.001818822, 
    0.001825995, 0.001828144, 0.001838188, 0.001834067, 0.001840623, 
    0.001834733, 0.001835777, 0.001840838, 0.001835051, 0.001847697, 
    0.001839128, 0.001855034, 0.001846489, 0.001855569, 0.001853921, 
    0.00185665, 0.001859093, 0.001862164, 0.001867828, 0.001866516, 
    0.001871249, 0.001822723, 0.001825645, 0.001825387, 0.001828443, 
    0.001830703, 0.001835596, 0.001843437, 0.001840489, 0.001845898, 
    0.001846984, 0.001838765, 0.001843813, 0.001827599, 0.001830223, 
    0.00182866, 0.001822954, 0.00184117, 0.001831829, 0.001849065, 
    0.001844013, 0.001858744, 0.001851424, 0.001865795, 0.001871929, 
    0.001877693, 0.001884425, 0.001827239, 0.001825254, 0.001828807, 
    0.00183372, 0.001838273, 0.001844322, 0.00184494, 0.001846072, 
    0.001849004, 0.001851468, 0.001846431, 0.001852086, 0.001830832, 
    0.001841979, 0.001824504, 0.001829772, 0.00183343, 0.001831825, 
    0.001840152, 0.001842113, 0.001850076, 0.001845961, 0.001870416, 
    0.001859609, 0.001889542, 0.001881194, 0.00182456, 0.001827231, 
    0.001836519, 0.001832102, 0.001844725, 0.001847828, 0.001850349, 
    0.001853571, 0.001853918, 0.001855826, 0.0018527, 0.001855703, 
    0.001844335, 0.001849417, 0.001835458, 0.001838859, 0.001837294, 
    0.001835578, 0.001840873, 0.001846511, 0.00184663, 0.001848437, 
    0.001853527, 0.001844776, 0.001871812, 0.001855132, 0.001830143, 
    0.001835283, 0.001836016, 0.001834026, 0.001847517, 0.001842632, 
    0.00185578, 0.001852229, 0.001858045, 0.001855156, 0.001854731, 
    0.001851017, 0.001848704, 0.001842857, 0.001838094, 0.001834314, 
    0.001835193, 0.001839345, 0.001846855, 0.00185395, 0.001852397, 
    0.001857603, 0.001843811, 0.001849599, 0.001847363, 0.001853191, 
    0.001840411, 0.001851299, 0.001837625, 0.001838825, 0.001842535, 
    0.001849992, 0.001851639, 0.001853398, 0.001852312, 0.001847045, 
    0.001846182, 0.001842445, 0.001841413, 0.001838564, 0.001836204, 
    0.00183836, 0.001840624, 0.001847047, 0.00185283, 0.001859128, 
    0.001860667, 0.001868017, 0.001862036, 0.001871904, 0.001863518, 
    0.001878026, 0.001851928, 0.001863269, 0.001842704, 0.001844923, 
    0.001848935, 0.001858124, 0.001853164, 0.001858964, 0.001846148, 
    0.001839488, 0.001837763, 0.001834544, 0.001837836, 0.001837569, 
    0.001840717, 0.001839706, 0.00184726, 0.001843203, 0.00185472, 
    0.001858918, 0.001870754, 0.001877998, 0.00188536, 0.001888608, 
    0.001889596, 0.001890009,
  0.001646087, 0.001653291, 0.001651891, 0.001657698, 0.001654477, 
    0.001658279, 0.001647547, 0.001653577, 0.001649728, 0.001646735, 
    0.00166896, 0.001657957, 0.001680371, 0.001673365, 0.001690952, 
    0.001679281, 0.001693303, 0.001690615, 0.001698702, 0.001696386, 
    0.001706724, 0.001699771, 0.001712076, 0.001705063, 0.001706161, 
    0.001699542, 0.001660172, 0.001667591, 0.001659732, 0.001660791, 
    0.001660316, 0.001654544, 0.001651634, 0.001645535, 0.001646643, 
    0.001651122, 0.001661266, 0.001657823, 0.001666497, 0.001666301, 
    0.001675947, 0.001671599, 0.001687796, 0.001683195, 0.001696483, 
    0.001693143, 0.001696326, 0.001695361, 0.001696339, 0.00169144, 
    0.001693539, 0.001689228, 0.001672414, 0.001677359, 0.001662602, 
    0.001653719, 0.001647812, 0.001643619, 0.001644212, 0.001645342, 
    0.001651148, 0.001656603, 0.001660758, 0.001663536, 0.001666273, 
    0.001674553, 0.001678931, 0.001688727, 0.001686959, 0.001689953, 
    0.001692811, 0.001697608, 0.001696819, 0.001698932, 0.001689873, 
    0.001695895, 0.001685952, 0.001688673, 0.001667019, 0.001658752, 
    0.001655239, 0.00165216, 0.001644668, 0.001649842, 0.001647803, 
    0.001652654, 0.001655735, 0.001654211, 0.001663612, 0.001659958, 
    0.00167919, 0.001670911, 0.001692478, 0.001687322, 0.001693713, 
    0.001690452, 0.001696039, 0.001691011, 0.001699718, 0.001701613, 
    0.001700318, 0.001705291, 0.001690732, 0.001696326, 0.001654169, 
    0.001654417, 0.001655575, 0.001650485, 0.001650173, 0.001645505, 
    0.001649659, 0.001651427, 0.001655914, 0.001658567, 0.001661088, 
    0.001666629, 0.001672814, 0.001681454, 0.001687656, 0.001691811, 
    0.001689263, 0.001691513, 0.001688998, 0.001687819, 0.001700903, 
    0.001693559, 0.001704575, 0.001703966, 0.001698982, 0.001704035, 
    0.001654592, 0.001653161, 0.001648194, 0.001652081, 0.001644997, 
    0.001648963, 0.001651244, 0.001660035, 0.001661965, 0.001663755, 
    0.001667289, 0.001671822, 0.001679768, 0.001686676, 0.001692977, 
    0.001692516, 0.001692678, 0.001694085, 0.001690599, 0.001694657, 
    0.001695339, 0.001693558, 0.001703885, 0.001700936, 0.001703953, 
    0.001702033, 0.001653626, 0.001656033, 0.001654733, 0.001657178, 
    0.001655455, 0.001663112, 0.001665407, 0.001676134, 0.001671733, 
    0.001678736, 0.001672444, 0.001673559, 0.001678966, 0.001672784, 
    0.001686296, 0.001677138, 0.00169414, 0.001685005, 0.001694712, 
    0.00169295, 0.001695867, 0.00169848, 0.001701765, 0.001707823, 
    0.00170642, 0.001711484, 0.001659619, 0.001662739, 0.001662464, 
    0.001665727, 0.00166814, 0.001673366, 0.001681743, 0.001678594, 
    0.001684374, 0.001685534, 0.001676752, 0.001682146, 0.001664826, 
    0.001667627, 0.001665959, 0.001659866, 0.00167932, 0.001669342, 
    0.001687759, 0.001682359, 0.001698107, 0.00169028, 0.001705648, 
    0.001712211, 0.00171838, 0.001725587, 0.00166444, 0.001662321, 
    0.001666115, 0.001671362, 0.001676226, 0.001682689, 0.00168335, 
    0.00168456, 0.001687694, 0.001690328, 0.001684943, 0.001690988, 
    0.001668277, 0.001680186, 0.00166152, 0.001667146, 0.001671052, 
    0.001669338, 0.001678234, 0.001680329, 0.001688839, 0.001684441, 
    0.001710592, 0.001699032, 0.001731069, 0.001722129, 0.001661581, 
    0.001664433, 0.001674352, 0.001669634, 0.00168312, 0.001686436, 
    0.001689131, 0.001692576, 0.001692947, 0.001694987, 0.001691644, 
    0.001694855, 0.001682703, 0.001688135, 0.001673219, 0.001676852, 
    0.00167518, 0.001673347, 0.001679004, 0.001685028, 0.001685156, 
    0.001687087, 0.001692527, 0.001683174, 0.001712085, 0.001694243, 
    0.001667542, 0.001673032, 0.001673815, 0.001671689, 0.001686104, 
    0.001680884, 0.001694937, 0.001691141, 0.00169736, 0.00169427, 
    0.001693816, 0.001689845, 0.001687373, 0.001681123, 0.001676035, 
    0.001671997, 0.001672936, 0.001677371, 0.001685396, 0.001692981, 
    0.00169132, 0.001696887, 0.001682143, 0.001688329, 0.001685939, 
    0.001692169, 0.00167851, 0.001690146, 0.001675534, 0.001676816, 
    0.00168078, 0.001688749, 0.00169051, 0.001692391, 0.00169123, 0.0016856, 
    0.001684677, 0.001680684, 0.001679581, 0.001676537, 0.001674016, 
    0.001676319, 0.001678738, 0.001685602, 0.001691783, 0.001698517, 
    0.001700164, 0.001708025, 0.001701627, 0.001712184, 0.001703211, 
    0.001718736, 0.001690818, 0.001702946, 0.00168096, 0.001683331, 
    0.001687619, 0.001697444, 0.00169214, 0.001698342, 0.00168464, 
    0.001677524, 0.001675681, 0.001672243, 0.001675759, 0.001675474, 
    0.001678837, 0.001677757, 0.001685829, 0.001681494, 0.001693804, 
    0.001698293, 0.001710954, 0.001718707, 0.00172659, 0.001730068, 
    0.001731126, 0.001731568,
  0.001514891, 0.001522022, 0.001520636, 0.001526387, 0.001523197, 
    0.001526962, 0.001516337, 0.001522306, 0.001518495, 0.001515533, 
    0.001537544, 0.001526643, 0.001548859, 0.001541911, 0.00155936, 
    0.001547779, 0.001561694, 0.001559025, 0.001567056, 0.001564756, 
    0.001575026, 0.001568118, 0.001580347, 0.001573376, 0.001574467, 
    0.00156789, 0.001528837, 0.001536188, 0.001528401, 0.00152945, 
    0.001528979, 0.001523263, 0.001520382, 0.001514346, 0.001515442, 
    0.001519875, 0.001529921, 0.001526511, 0.001535103, 0.001534909, 
    0.001544472, 0.001540161, 0.001556227, 0.001551662, 0.001564852, 
    0.001561535, 0.001564696, 0.001563738, 0.001564708, 0.001559845, 
    0.001561929, 0.001557648, 0.001540968, 0.001545872, 0.001531245, 
    0.001522446, 0.001516599, 0.001512449, 0.001513036, 0.001514154, 
    0.001519901, 0.001525302, 0.001529417, 0.00153217, 0.001534881, 
    0.001543089, 0.001547431, 0.001557151, 0.001555396, 0.001558368, 
    0.001561205, 0.001565969, 0.001565185, 0.001567284, 0.001558289, 
    0.001564268, 0.001554397, 0.001557097, 0.001535621, 0.001527431, 
    0.001523951, 0.001520903, 0.001513487, 0.001518609, 0.00151659, 
    0.001521392, 0.001524443, 0.001522934, 0.001532245, 0.001528625, 
    0.001547688, 0.001539479, 0.001560874, 0.001555756, 0.001562101, 
    0.001558864, 0.001564411, 0.001559418, 0.001568065, 0.001569948, 
    0.001568661, 0.001573602, 0.001559142, 0.001564696, 0.001522891, 
    0.001523138, 0.001524284, 0.001519244, 0.001518936, 0.001514316, 
    0.001518427, 0.001520177, 0.001524619, 0.001527247, 0.001529744, 
    0.001535235, 0.001541365, 0.001549934, 0.001556088, 0.001560212, 
    0.001557683, 0.001559916, 0.00155742, 0.00155625, 0.001569242, 
    0.001561948, 0.001572891, 0.001572286, 0.001567334, 0.001572354, 
    0.00152331, 0.001521894, 0.001516977, 0.001520825, 0.001513813, 
    0.001517738, 0.001519996, 0.001528702, 0.001530613, 0.001532387, 
    0.001535888, 0.001540381, 0.001548262, 0.001555116, 0.00156137, 
    0.001560912, 0.001561073, 0.001562471, 0.00155901, 0.001563039, 
    0.001563715, 0.001561947, 0.001572205, 0.001569275, 0.001572273, 
    0.001570365, 0.001522354, 0.001524737, 0.00152345, 0.001525871, 
    0.001524166, 0.00153175, 0.001534023, 0.001544658, 0.001540293, 
    0.001547238, 0.001540999, 0.001542104, 0.001547466, 0.001541336, 
    0.001554738, 0.001545653, 0.001562525, 0.001553457, 0.001563093, 
    0.001561343, 0.00156424, 0.001566835, 0.001570098, 0.001576119, 
    0.001574725, 0.001579758, 0.001528289, 0.00153138, 0.001531107, 
    0.001534341, 0.001536732, 0.001541913, 0.001550221, 0.001547097, 
    0.001552831, 0.001553982, 0.00154527, 0.00155062, 0.001533447, 
    0.001536223, 0.00153457, 0.001528533, 0.001547817, 0.001537923, 
    0.00155619, 0.001550832, 0.001566465, 0.001558692, 0.001573957, 
    0.001580481, 0.001586617, 0.001593787, 0.001533066, 0.001530966, 
    0.001534725, 0.001539925, 0.001544748, 0.001551159, 0.001551815, 
    0.001553016, 0.001556126, 0.00155874, 0.001553396, 0.001559396, 
    0.001536868, 0.001548676, 0.001530173, 0.001535747, 0.001539619, 
    0.00153792, 0.00154674, 0.001548818, 0.001557262, 0.001552897, 
    0.001578871, 0.001567384, 0.001599244, 0.001590346, 0.001530233, 
    0.001533058, 0.001542891, 0.001538213, 0.001551587, 0.001554878, 
    0.001557552, 0.001560972, 0.001561341, 0.001563366, 0.001560047, 
    0.001563235, 0.001551173, 0.001556564, 0.001541766, 0.001545369, 
    0.001543712, 0.001541894, 0.001547504, 0.00155348, 0.001553607, 
    0.001555523, 0.001560923, 0.001551641, 0.001580355, 0.001562627, 
    0.001536139, 0.001541581, 0.001542357, 0.00154025, 0.001554548, 
    0.001549368, 0.001563317, 0.001559547, 0.001565723, 0.001562654, 
    0.001562203, 0.001558261, 0.001555807, 0.001549606, 0.001544559, 
    0.001540555, 0.001541486, 0.001545884, 0.001553845, 0.001561374, 
    0.001559725, 0.001565253, 0.001550617, 0.001556756, 0.001554384, 
    0.001560569, 0.001547014, 0.001558559, 0.001544062, 0.001545334, 
    0.001549265, 0.001557173, 0.001558921, 0.001560788, 0.001559636, 
    0.001554047, 0.001553131, 0.00154917, 0.001548076, 0.001545057, 
    0.001542557, 0.001544841, 0.00154724, 0.001554049, 0.001560185, 
    0.001566872, 0.001568508, 0.00157632, 0.001569962, 0.001580454, 
    0.001571535, 0.001586971, 0.001559227, 0.001571272, 0.001549444, 
    0.001551796, 0.001556051, 0.001565806, 0.001560539, 0.001566698, 
    0.001553095, 0.001546036, 0.001544208, 0.001540799, 0.001544286, 
    0.001544002, 0.001547339, 0.001546266, 0.001554275, 0.001549974, 
    0.001562192, 0.001566649, 0.001579231, 0.001586941, 0.001594785, 
    0.001598248, 0.001599301, 0.001599742,
  0.0013795, 0.001385892, 0.001384649, 0.001389807, 0.001386945, 0.001390324, 
    0.001380796, 0.001386147, 0.00138273, 0.001380075, 0.001399825, 
    0.001390037, 0.001409999, 0.00140375, 0.001419454, 0.001409027, 
    0.001421558, 0.001419152, 0.001426392, 0.001424317, 0.001433584, 
    0.001427349, 0.00143839, 0.001432094, 0.001433079, 0.001427144, 
    0.001392006, 0.001398606, 0.001391615, 0.001392556, 0.001392134, 
    0.001387005, 0.001384422, 0.001379012, 0.001379993, 0.001383967, 
    0.001392979, 0.001389918, 0.001397632, 0.001397458, 0.001406052, 
    0.001402176, 0.001416632, 0.001412521, 0.001424404, 0.001421414, 
    0.001424263, 0.001423399, 0.001424275, 0.001419891, 0.001421769, 
    0.001417912, 0.001402902, 0.001407311, 0.001394167, 0.001386273, 
    0.00138103, 0.001377313, 0.001377838, 0.00137884, 0.00138399, 
    0.001388834, 0.001392527, 0.001394998, 0.001397433, 0.001404809, 
    0.001408714, 0.001417464, 0.001415883, 0.00141856, 0.001421117, 
    0.001425412, 0.001424705, 0.001426598, 0.001418489, 0.001423877, 
    0.001414984, 0.001417415, 0.001398097, 0.001390744, 0.001387622, 
    0.001384888, 0.001378242, 0.001382832, 0.001381022, 0.001385327, 
    0.001388063, 0.00138671, 0.001395065, 0.001391816, 0.001408946, 
    0.001401564, 0.001420819, 0.001416208, 0.001421924, 0.001419007, 
    0.001424006, 0.001419507, 0.001427302, 0.001429, 0.00142784, 0.001432298, 
    0.001419257, 0.001424264, 0.001386672, 0.001386893, 0.001387921, 
    0.001383402, 0.001383125, 0.001378985, 0.001382669, 0.001384238, 
    0.001388222, 0.001390579, 0.001392821, 0.00139775, 0.001403259, 
    0.001410966, 0.001416507, 0.001420222, 0.001417944, 0.001419955, 
    0.001417706, 0.001416653, 0.001428364, 0.001421786, 0.001431657, 
    0.00143111, 0.001426643, 0.001431172, 0.001387047, 0.001385777, 
    0.001381369, 0.001384819, 0.001378534, 0.001382052, 0.001384075, 
    0.001391885, 0.0013936, 0.001395193, 0.001398337, 0.001402375, 
    0.001409461, 0.001415631, 0.001421266, 0.001420853, 0.001420998, 
    0.001422257, 0.001419138, 0.00142277, 0.001423379, 0.001421785, 
    0.001431037, 0.001428393, 0.001431099, 0.001429377, 0.00138619, 
    0.001388327, 0.001387172, 0.001389345, 0.001387815, 0.001394621, 
    0.001396662, 0.001406219, 0.001402295, 0.00140854, 0.001402929, 
    0.001403924, 0.001408745, 0.001403232, 0.001415291, 0.001407115, 
    0.001422306, 0.001414137, 0.001422819, 0.001421241, 0.001423853, 
    0.001426192, 0.001429136, 0.001434571, 0.001433312, 0.001437858, 
    0.001391515, 0.001394288, 0.001394044, 0.001396947, 0.001399095, 
    0.001403751, 0.001411224, 0.001408413, 0.001413574, 0.00141461, 
    0.00140677, 0.001411584, 0.001396145, 0.001398638, 0.001397153, 
    0.001391734, 0.001409062, 0.001400165, 0.001416598, 0.001411774, 
    0.001425859, 0.001418852, 0.001432619, 0.001438511, 0.001444058, 
    0.001450546, 0.001395802, 0.001393917, 0.001397292, 0.001401965, 
    0.001406301, 0.001412069, 0.001412659, 0.00141374, 0.00141654, 
    0.001418896, 0.001414082, 0.001419486, 0.001399218, 0.001409834, 
    0.001393205, 0.00139821, 0.001401689, 0.001400162, 0.001408092, 
    0.001409962, 0.001417564, 0.001413633, 0.001437057, 0.001426687, 
    0.001455488, 0.001447431, 0.001393259, 0.001395796, 0.00140463, 
    0.001400426, 0.001412454, 0.001415417, 0.001417825, 0.001420906, 
    0.001421239, 0.001423065, 0.001420073, 0.001422946, 0.001412081, 
    0.001416935, 0.00140362, 0.001406859, 0.001405369, 0.001403734, 
    0.001408779, 0.001414158, 0.001414272, 0.001415998, 0.001420863, 
    0.001412502, 0.001438398, 0.001422399, 0.001398563, 0.001403453, 
    0.001404151, 0.001402256, 0.00141512, 0.001410457, 0.00142302, 
    0.001419623, 0.001425189, 0.001422423, 0.001422016, 0.001418464, 
    0.001416254, 0.001410671, 0.00140613, 0.001402531, 0.001403368, 
    0.001407322, 0.001414487, 0.001421269, 0.001419783, 0.001424766, 
    0.001411581, 0.001417108, 0.001414972, 0.001420543, 0.001408339, 
    0.001418733, 0.001405684, 0.001406827, 0.001410364, 0.001417484, 
    0.001419058, 0.001420741, 0.001419702, 0.001414669, 0.001413844, 
    0.001410278, 0.001409294, 0.001406578, 0.00140433, 0.001406384, 
    0.001408542, 0.001414671, 0.001420197, 0.001426226, 0.001427701, 
    0.001434753, 0.001429013, 0.001438487, 0.001430434, 0.001444378, 
    0.001419334, 0.001430195, 0.001410525, 0.001412642, 0.001416474, 
    0.001425264, 0.001420517, 0.001426069, 0.001413812, 0.001407459, 
    0.001405815, 0.00140275, 0.001405885, 0.00140563, 0.001408631, 
    0.001407666, 0.001414874, 0.001411002, 0.001422006, 0.001426025, 
    0.001437382, 0.001444351, 0.001451449, 0.001454585, 0.00145554, 
    0.001455939,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.34869e-06, 1.360238e-06, 1.357989e-06, 1.367333e-06, 1.362145e-06, 
    1.368269e-06, 1.351026e-06, 1.360697e-06, 1.354519e-06, 1.349726e-06, 
    1.385558e-06, 1.367749e-06, 1.404176e-06, 1.392728e-06, 1.421575e-06, 
    1.402392e-06, 1.425458e-06, 1.421018e-06, 1.4344e-06, 1.43056e-06, 
    1.447748e-06, 1.436174e-06, 1.456697e-06, 1.444979e-06, 1.446809e-06, 
    1.435792e-06, 1.371323e-06, 1.383336e-06, 1.370613e-06, 1.372323e-06, 
    1.371555e-06, 1.362252e-06, 1.357576e-06, 1.347807e-06, 1.349578e-06, 
    1.356754e-06, 1.373091e-06, 1.367533e-06, 1.381559e-06, 1.381241e-06, 
    1.39694e-06, 1.389851e-06, 1.416371e-06, 1.408807e-06, 1.43072e-06, 
    1.425193e-06, 1.43046e-06, 1.428861e-06, 1.43048e-06, 1.422379e-06, 
    1.425847e-06, 1.418728e-06, 1.391179e-06, 1.399248e-06, 1.375252e-06, 
    1.360925e-06, 1.351449e-06, 1.344746e-06, 1.345692e-06, 1.347498e-06, 
    1.356795e-06, 1.365565e-06, 1.372268e-06, 1.376761e-06, 1.381195e-06, 
    1.394665e-06, 1.401818e-06, 1.417904e-06, 1.414993e-06, 1.419925e-06, 
    1.424643e-06, 1.432585e-06, 1.431276e-06, 1.43478e-06, 1.419793e-06, 
    1.429745e-06, 1.413335e-06, 1.417814e-06, 1.382407e-06, 1.369031e-06, 
    1.363369e-06, 1.35842e-06, 1.34642e-06, 1.354701e-06, 1.351434e-06, 
    1.359213e-06, 1.364168e-06, 1.361716e-06, 1.376884e-06, 1.370977e-06, 
    1.402242e-06, 1.388731e-06, 1.424093e-06, 1.415589e-06, 1.426134e-06, 
    1.420748e-06, 1.429983e-06, 1.42167e-06, 1.436085e-06, 1.439234e-06, 
    1.437081e-06, 1.445356e-06, 1.421209e-06, 1.430459e-06, 1.361648e-06, 
    1.362048e-06, 1.36391e-06, 1.355731e-06, 1.355232e-06, 1.347758e-06, 
    1.354406e-06, 1.357243e-06, 1.364455e-06, 1.368731e-06, 1.372801e-06, 
    1.381773e-06, 1.391829e-06, 1.40595e-06, 1.41614e-06, 1.422991e-06, 
    1.418787e-06, 1.422498e-06, 1.41835e-06, 1.416408e-06, 1.438053e-06, 
    1.425879e-06, 1.444164e-06, 1.443149e-06, 1.434862e-06, 1.443263e-06, 
    1.362328e-06, 1.360028e-06, 1.352059e-06, 1.358293e-06, 1.346945e-06, 
    1.353292e-06, 1.356948e-06, 1.371101e-06, 1.374219e-06, 1.377115e-06, 
    1.382843e-06, 1.390212e-06, 1.403188e-06, 1.414526e-06, 1.424917e-06, 
    1.424154e-06, 1.424423e-06, 1.426749e-06, 1.42099e-06, 1.427695e-06, 
    1.428823e-06, 1.425876e-06, 1.443013e-06, 1.438106e-06, 1.443127e-06, 
    1.439931e-06, 1.360775e-06, 1.364647e-06, 1.362554e-06, 1.366491e-06, 
    1.363717e-06, 1.376075e-06, 1.37979e-06, 1.397245e-06, 1.390067e-06, 
    1.401499e-06, 1.391225e-06, 1.393043e-06, 1.401874e-06, 1.391779e-06, 
    1.4139e-06, 1.398885e-06, 1.42684e-06, 1.411777e-06, 1.427786e-06, 
    1.424871e-06, 1.429698e-06, 1.434028e-06, 1.439484e-06, 1.449581e-06, 
    1.447239e-06, 1.455703e-06, 1.370429e-06, 1.37547e-06, 1.375025e-06, 
    1.38031e-06, 1.384225e-06, 1.392729e-06, 1.406424e-06, 1.401265e-06, 
    1.410741e-06, 1.412648e-06, 1.398253e-06, 1.407083e-06, 1.378848e-06, 
    1.38339e-06, 1.380684e-06, 1.370825e-06, 1.402453e-06, 1.386176e-06, 
    1.416307e-06, 1.407433e-06, 1.43341e-06, 1.420462e-06, 1.445951e-06, 
    1.45692e-06, 1.467278e-06, 1.479434e-06, 1.378225e-06, 1.374794e-06, 
    1.380938e-06, 1.389463e-06, 1.397394e-06, 1.407975e-06, 1.409059e-06, 
    1.411047e-06, 1.416201e-06, 1.420542e-06, 1.411676e-06, 1.421631e-06, 
    1.384446e-06, 1.40387e-06, 1.373498e-06, 1.382609e-06, 1.388958e-06, 
    1.38617e-06, 1.400674e-06, 1.404104e-06, 1.418086e-06, 1.410849e-06, 
    1.454209e-06, 1.434944e-06, 1.488721e-06, 1.473592e-06, 1.373597e-06, 
    1.378212e-06, 1.394336e-06, 1.386652e-06, 1.408682e-06, 1.414132e-06, 
    1.418569e-06, 1.424253e-06, 1.424867e-06, 1.428241e-06, 1.422714e-06, 
    1.428022e-06, 1.407996e-06, 1.416927e-06, 1.392486e-06, 1.398415e-06, 
    1.395685e-06, 1.392695e-06, 1.401934e-06, 1.411814e-06, 1.412024e-06, 
    1.415199e-06, 1.42417e-06, 1.408769e-06, 1.456707e-06, 1.427008e-06, 
    1.383253e-06, 1.392183e-06, 1.393459e-06, 1.389995e-06, 1.413585e-06, 
    1.405014e-06, 1.428158e-06, 1.421884e-06, 1.432171e-06, 1.427054e-06, 
    1.426302e-06, 1.419746e-06, 1.415672e-06, 1.405406e-06, 1.39708e-06, 
    1.390495e-06, 1.392025e-06, 1.399263e-06, 1.412419e-06, 1.424921e-06, 
    1.422178e-06, 1.431386e-06, 1.407076e-06, 1.417244e-06, 1.41331e-06, 
    1.42358e-06, 1.401128e-06, 1.420242e-06, 1.396264e-06, 1.398357e-06, 
    1.404844e-06, 1.417939e-06, 1.420842e-06, 1.423947e-06, 1.42203e-06, 
    1.412754e-06, 1.411237e-06, 1.404685e-06, 1.402879e-06, 1.3979e-06, 
    1.393785e-06, 1.397545e-06, 1.401498e-06, 1.412756e-06, 1.422942e-06, 
    1.434088e-06, 1.436822e-06, 1.449917e-06, 1.439254e-06, 1.456873e-06, 
    1.441889e-06, 1.467875e-06, 1.421351e-06, 1.44145e-06, 1.405139e-06, 
    1.409028e-06, 1.416077e-06, 1.432309e-06, 1.423533e-06, 1.433799e-06, 
    1.411177e-06, 1.399514e-06, 1.396502e-06, 1.390895e-06, 1.39663e-06, 
    1.396163e-06, 1.401661e-06, 1.399893e-06, 1.413131e-06, 1.406012e-06, 
    1.426282e-06, 1.433716e-06, 1.454814e-06, 1.467825e-06, 1.481128e-06, 
    1.487021e-06, 1.488817e-06, 1.489568e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.295124e-06, 8.33173e-06, 8.32459e-06, 8.35414e-06, 8.337733e-06, 
    8.357074e-06, 8.302497e-06, 8.333132e-06, 8.313559e-06, 8.298343e-06, 
    8.411485e-06, 8.355393e-06, 8.469779e-06, 8.433943e-06, 8.523965e-06, 
    8.464186e-06, 8.536018e-06, 8.522208e-06, 8.563719e-06, 8.551809e-06, 
    8.604957e-06, 8.569189e-06, 8.632504e-06, 8.596393e-06, 8.602034e-06, 
    8.567971e-06, 8.366723e-06, 8.404561e-06, 8.364469e-06, 8.369863e-06, 
    8.367431e-06, 8.33804e-06, 8.323246e-06, 8.292246e-06, 8.297858e-06, 
    8.320617e-06, 8.372229e-06, 8.354679e-06, 8.398863e-06, 8.397866e-06, 
    8.447106e-06, 8.424891e-06, 8.507747e-06, 8.484165e-06, 8.552296e-06, 
    8.53514e-06, 8.551476e-06, 8.546507e-06, 8.551517e-06, 8.526378e-06, 
    8.53713e-06, 8.515013e-06, 8.42915e-06, 8.45441e-06, 8.379078e-06, 
    8.333848e-06, 8.303808e-06, 8.282522e-06, 8.285513e-06, 8.291253e-06, 
    8.320733e-06, 8.34846e-06, 8.36961e-06, 8.383756e-06, 8.397698e-06, 
    8.439987e-06, 8.462353e-06, 8.5125e-06, 8.503433e-06, 8.51877e-06, 
    8.533425e-06, 8.558044e-06, 8.553984e-06, 8.564828e-06, 8.518316e-06, 
    8.549221e-06, 8.4982e-06, 8.512147e-06, 8.401606e-06, 8.359445e-06, 
    8.341567e-06, 8.32589e-06, 8.287821e-06, 8.314104e-06, 8.303732e-06, 
    8.328367e-06, 8.344036e-06, 8.33627e-06, 8.384134e-06, 8.365507e-06, 
    8.463667e-06, 8.421356e-06, 8.531726e-06, 8.505273e-06, 8.538041e-06, 
    8.521312e-06, 8.549966e-06, 8.524163e-06, 8.56885e-06, 8.578596e-06, 
    8.571919e-06, 8.597493e-06, 8.522682e-06, 8.551397e-06, 8.336102e-06, 
    8.337369e-06, 8.343247e-06, 8.317355e-06, 8.315767e-06, 8.292045e-06, 
    8.313128e-06, 8.322118e-06, 8.344921e-06, 8.358415e-06, 8.371245e-06, 
    8.399494e-06, 8.431056e-06, 8.475222e-06, 8.506978e-06, 8.528269e-06, 
    8.515199e-06, 8.526722e-06, 8.513824e-06, 8.507768e-06, 8.574923e-06, 
    8.537201e-06, 8.593789e-06, 8.590656e-06, 8.565024e-06, 8.590986e-06, 
    8.33824e-06, 8.330951e-06, 8.305704e-06, 8.325445e-06, 8.289447e-06, 
    8.309593e-06, 8.321172e-06, 8.365892e-06, 8.375707e-06, 8.384833e-06, 
    8.402841e-06, 8.425966e-06, 8.466583e-06, 8.50194e-06, 8.534244e-06, 
    8.531862e-06, 8.532693e-06, 8.539903e-06, 8.522014e-06, 8.542824e-06, 
    8.546312e-06, 8.537171e-06, 8.590213e-06, 8.575049e-06, 8.590557e-06, 
    8.580668e-06, 8.333306e-06, 8.345537e-06, 8.33891e-06, 8.351356e-06, 
    8.342573e-06, 8.38157e-06, 8.393258e-06, 8.448018e-06, 8.425513e-06, 
    8.461311e-06, 8.429129e-06, 8.434829e-06, 8.462465e-06, 8.430842e-06, 
    8.49997e-06, 8.453088e-06, 8.540175e-06, 8.493331e-06, 8.543096e-06, 
    8.534036e-06, 8.549001e-06, 8.562423e-06, 8.579287e-06, 8.610465e-06, 
    8.603224e-06, 8.629304e-06, 8.363784e-06, 8.379668e-06, 8.378259e-06, 
    8.394883e-06, 8.407182e-06, 8.433867e-06, 8.476693e-06, 8.460565e-06, 
    8.490138e-06, 8.496083e-06, 8.451118e-06, 8.478717e-06, 8.390221e-06, 
    8.404499e-06, 8.395982e-06, 8.364917e-06, 8.464219e-06, 8.413218e-06, 
    8.507406e-06, 8.479738e-06, 8.560486e-06, 8.520313e-06, 8.599244e-06, 
    8.633052e-06, 8.66485e-06, 8.702066e-06, 8.38833e-06, 8.377514e-06, 
    8.396843e-06, 8.423628e-06, 8.448457e-06, 8.481524e-06, 8.484893e-06, 
    8.49108e-06, 8.507123e-06, 8.52063e-06, 8.493026e-06, 8.523993e-06, 
    8.407816e-06, 8.468643e-06, 8.373328e-06, 8.402016e-06, 8.421932e-06, 
    8.413182e-06, 8.458616e-06, 8.469323e-06, 8.512901e-06, 8.490362e-06, 
    8.624687e-06, 8.565206e-06, 8.730394e-06, 8.684178e-06, 8.373732e-06, 
    8.388255e-06, 8.438879e-06, 8.414781e-06, 8.483705e-06, 8.500695e-06, 
    8.514487e-06, 8.532158e-06, 8.534043e-06, 8.544517e-06, 8.52734e-06, 
    8.543821e-06, 8.481506e-06, 8.509335e-06, 8.432992e-06, 8.45155e-06, 
    8.443e-06, 8.43362e-06, 8.462528e-06, 8.493371e-06, 8.494008e-06, 
    8.503891e-06, 8.531801e-06, 8.483832e-06, 8.632357e-06, 8.540578e-06, 
    8.404103e-06, 8.432125e-06, 8.436108e-06, 8.425249e-06, 8.498968e-06, 
    8.47224e-06, 8.54426e-06, 8.524767e-06, 8.556676e-06, 8.540814e-06, 
    8.538463e-06, 8.518096e-06, 8.505405e-06, 8.473402e-06, 8.447357e-06, 
    8.426726e-06, 8.431504e-06, 8.454173e-06, 8.495231e-06, 8.534119e-06, 
    8.525588e-06, 8.554146e-06, 8.478534e-06, 8.510227e-06, 8.497961e-06, 
    8.529904e-06, 8.460105e-06, 8.519713e-06, 8.444877e-06, 8.451418e-06, 
    8.471685e-06, 8.512508e-06, 8.521512e-06, 8.531166e-06, 8.52519e-06, 
    8.496333e-06, 8.491593e-06, 8.471136e-06, 8.465488e-06, 8.449917e-06, 
    8.437015e-06, 8.44879e-06, 8.461142e-06, 8.496278e-06, 8.527955e-06, 
    8.562514e-06, 8.570971e-06, 8.611415e-06, 8.578489e-06, 8.632829e-06, 
    8.586631e-06, 8.6666e-06, 8.523131e-06, 8.585423e-06, 8.472606e-06, 
    8.484731e-06, 8.506699e-06, 8.557097e-06, 8.529854e-06, 8.561701e-06, 
    8.491401e-06, 8.454974e-06, 8.445534e-06, 8.42797e-06, 8.44592e-06, 
    8.44446e-06, 8.461649e-06, 8.456108e-06, 8.49742e-06, 8.47522e-06, 
    8.538298e-06, 8.561349e-06, 8.626479e-06, 8.666447e-06, 8.707158e-06, 
    8.725135e-06, 8.730607e-06, 8.732887e-06,
  4.945751e-06, 4.982884e-06, 4.975656e-06, 5.005666e-06, 4.98901e-06, 
    5.008672e-06, 4.95327e-06, 4.984362e-06, 4.964504e-06, 4.949087e-06, 
    5.064093e-06, 5.007006e-06, 5.123616e-06, 5.087033e-06, 5.179099e-06, 
    5.117919e-06, 5.191465e-06, 5.177326e-06, 5.219911e-06, 5.207698e-06, 
    5.262306e-06, 5.22555e-06, 5.290683e-06, 5.253517e-06, 5.259328e-06, 
    5.224339e-06, 5.018472e-06, 5.056974e-06, 5.016195e-06, 5.021678e-06, 
    5.019217e-06, 4.989355e-06, 4.974333e-06, 4.942914e-06, 4.948612e-06, 
    4.97169e-06, 5.024144e-06, 5.006313e-06, 5.051286e-06, 5.050269e-06, 
    5.100503e-06, 5.077832e-06, 5.162522e-06, 5.1384e-06, 5.208208e-06, 
    5.190622e-06, 5.207382e-06, 5.202297e-06, 5.207448e-06, 5.181665e-06, 
    5.192706e-06, 5.170037e-06, 5.082076e-06, 5.107874e-06, 5.031071e-06, 
    4.985096e-06, 4.954632e-06, 4.933059e-06, 4.936107e-06, 4.94192e-06, 
    4.971825e-06, 4.999998e-06, 5.021507e-06, 5.035914e-06, 5.050123e-06, 
    5.093229e-06, 5.116087e-06, 5.167406e-06, 5.158128e-06, 5.173847e-06, 
    5.188873e-06, 5.214141e-06, 5.209979e-06, 5.221122e-06, 5.173429e-06, 
    5.20511e-06, 5.152846e-06, 5.167123e-06, 5.054002e-06, 5.011121e-06, 
    4.992946e-06, 4.977046e-06, 4.938451e-06, 4.965093e-06, 4.954585e-06, 
    4.979595e-06, 4.995512e-06, 4.987637e-06, 5.036308e-06, 5.017366e-06, 
    5.117443e-06, 5.074251e-06, 5.18712e-06, 5.160031e-06, 5.193619e-06, 
    5.17647e-06, 5.205868e-06, 5.179407e-06, 5.22527e-06, 5.235277e-06, 
    5.228438e-06, 5.25472e-06, 5.177942e-06, 5.207383e-06, 4.987417e-06, 
    4.988701e-06, 4.994684e-06, 4.968405e-06, 4.966799e-06, 4.942759e-06, 
    4.964146e-06, 4.973265e-06, 4.996435e-06, 5.01016e-06, 5.02322e-06, 
    5.051976e-06, 5.084161e-06, 5.129285e-06, 5.161786e-06, 5.183613e-06, 
    5.170224e-06, 5.182044e-06, 5.168832e-06, 5.162643e-06, 5.231528e-06, 
    5.19281e-06, 5.250937e-06, 5.247714e-06, 5.221387e-06, 5.248077e-06, 
    4.989603e-06, 4.982215e-06, 4.956598e-06, 4.976641e-06, 4.940143e-06, 
    4.960563e-06, 4.972318e-06, 5.017765e-06, 5.027766e-06, 5.037051e-06, 
    5.055403e-06, 5.078991e-06, 5.120465e-06, 5.156644e-06, 5.189747e-06, 
    5.187319e-06, 5.188174e-06, 5.19558e-06, 5.177244e-06, 5.198592e-06, 
    5.202179e-06, 5.192804e-06, 5.247283e-06, 5.231698e-06, 5.247646e-06, 
    5.237496e-06, 4.984615e-06, 4.997051e-06, 4.99033e-06, 5.002972e-06, 
    4.994065e-06, 5.033715e-06, 5.045625e-06, 5.10148e-06, 5.078527e-06, 
    5.115071e-06, 5.082234e-06, 5.088048e-06, 5.11627e-06, 5.084006e-06, 
    5.15465e-06, 5.106723e-06, 5.195868e-06, 5.14788e-06, 5.19888e-06, 
    5.189604e-06, 5.204964e-06, 5.218736e-06, 5.236077e-06, 5.268129e-06, 
    5.2607e-06, 5.287541e-06, 5.015609e-06, 5.031778e-06, 5.030351e-06, 
    5.047288e-06, 5.059828e-06, 5.087041e-06, 5.130797e-06, 5.114326e-06, 
    5.144575e-06, 5.150655e-06, 5.104705e-06, 5.132903e-06, 5.042607e-06, 
    5.057161e-06, 5.048492e-06, 5.016886e-06, 5.118124e-06, 5.06608e-06, 
    5.162324e-06, 5.134022e-06, 5.216772e-06, 5.175564e-06, 5.256613e-06, 
    5.291399e-06, 5.324197e-06, 5.362626e-06, 5.040607e-06, 5.029613e-06, 
    5.049303e-06, 5.076596e-06, 5.101957e-06, 5.135747e-06, 5.139208e-06, 
    5.145549e-06, 5.161984e-06, 5.175817e-06, 5.147557e-06, 5.179287e-06, 
    5.060543e-06, 5.122648e-06, 5.02546e-06, 5.05466e-06, 5.074984e-06, 
    5.066062e-06, 5.112444e-06, 5.123398e-06, 5.167997e-06, 5.144924e-06, 
    5.282809e-06, 5.22165e-06, 5.39194e-06, 5.344168e-06, 5.025774e-06, 
    5.040568e-06, 5.092183e-06, 5.067601e-06, 5.138004e-06, 5.155387e-06, 
    5.169531e-06, 5.187635e-06, 5.189589e-06, 5.200327e-06, 5.182736e-06, 
    5.199631e-06, 5.135819e-06, 5.164301e-06, 5.08627e-06, 5.105226e-06, 
    5.096502e-06, 5.08694e-06, 5.116471e-06, 5.148002e-06, 5.148672e-06, 
    5.158798e-06, 5.187378e-06, 5.13829e-06, 5.290728e-06, 5.196412e-06, 
    5.056719e-06, 5.085297e-06, 5.089379e-06, 5.0783e-06, 5.153644e-06, 
    5.1263e-06, 5.200065e-06, 5.180092e-06, 5.21283e-06, 5.196554e-06, 
    5.19416e-06, 5.173283e-06, 5.160301e-06, 5.127553e-06, 5.10096e-06, 
    5.079905e-06, 5.084798e-06, 5.107936e-06, 5.149932e-06, 5.189768e-06, 
    5.181033e-06, 5.21034e-06, 5.132888e-06, 5.165318e-06, 5.152777e-06, 
    5.185499e-06, 5.11389e-06, 5.174861e-06, 5.098347e-06, 5.105039e-06, 
    5.125757e-06, 5.167523e-06, 5.176773e-06, 5.186664e-06, 5.180559e-06, 
    5.150999e-06, 5.14616e-06, 5.125252e-06, 5.119487e-06, 5.103581e-06, 
    5.090428e-06, 5.102446e-06, 5.115079e-06, 5.15101e-06, 5.183467e-06, 
    5.218933e-06, 5.227623e-06, 5.269202e-06, 5.235352e-06, 5.291256e-06, 
    5.243723e-06, 5.326092e-06, 5.178395e-06, 5.242319e-06, 5.126699e-06, 
    5.139111e-06, 5.161592e-06, 5.213273e-06, 5.185345e-06, 5.218009e-06, 
    5.14597e-06, 5.108737e-06, 5.099114e-06, 5.081185e-06, 5.099524e-06, 
    5.098031e-06, 5.1156e-06, 5.109951e-06, 5.152204e-06, 5.129492e-06, 
    5.194101e-06, 5.21775e-06, 5.284727e-06, 5.325933e-06, 5.367981e-06, 
    5.386582e-06, 5.392248e-06, 5.394617e-06,
  4.461286e-06, 4.50057e-06, 4.492922e-06, 4.52469e-06, 4.507055e-06, 
    4.527874e-06, 4.469238e-06, 4.502134e-06, 4.481122e-06, 4.464815e-06, 
    4.586609e-06, 4.526109e-06, 4.64979e-06, 4.610951e-06, 4.708768e-06, 
    4.643739e-06, 4.721924e-06, 4.706884e-06, 4.752203e-06, 4.739202e-06, 
    4.797367e-06, 4.758209e-06, 4.827627e-06, 4.788002e-06, 4.794194e-06, 
    4.75692e-06, 4.538255e-06, 4.579059e-06, 4.535842e-06, 4.54165e-06, 
    4.539043e-06, 4.507419e-06, 4.49152e-06, 4.458288e-06, 4.464313e-06, 
    4.488723e-06, 4.544263e-06, 4.525376e-06, 4.573033e-06, 4.571954e-06, 
    4.625248e-06, 4.601188e-06, 4.69114e-06, 4.6655e-06, 4.739744e-06, 
    4.721028e-06, 4.738865e-06, 4.733453e-06, 4.738936e-06, 4.711498e-06, 
    4.723246e-06, 4.699131e-06, 4.60569e-06, 4.633073e-06, 4.551604e-06, 
    4.502909e-06, 4.470679e-06, 4.447869e-06, 4.451091e-06, 4.457236e-06, 
    4.488867e-06, 4.518688e-06, 4.54147e-06, 4.556737e-06, 4.571799e-06, 
    4.617524e-06, 4.641794e-06, 4.696332e-06, 4.686468e-06, 4.703182e-06, 
    4.719168e-06, 4.74606e-06, 4.741629e-06, 4.753493e-06, 4.702739e-06, 
    4.736446e-06, 4.680854e-06, 4.696033e-06, 4.575907e-06, 4.530468e-06, 
    4.511219e-06, 4.494392e-06, 4.453569e-06, 4.481744e-06, 4.470628e-06, 
    4.49709e-06, 4.513939e-06, 4.505602e-06, 4.557155e-06, 4.537084e-06, 
    4.643235e-06, 4.597388e-06, 4.717302e-06, 4.688492e-06, 4.724218e-06, 
    4.705973e-06, 4.737253e-06, 4.709098e-06, 4.757911e-06, 4.768568e-06, 
    4.761284e-06, 4.789285e-06, 4.707539e-06, 4.738866e-06, 4.505369e-06, 
    4.506729e-06, 4.513062e-06, 4.485248e-06, 4.483548e-06, 4.458123e-06, 
    4.480743e-06, 4.49039e-06, 4.514916e-06, 4.529451e-06, 4.543285e-06, 
    4.573763e-06, 4.607903e-06, 4.655813e-06, 4.690357e-06, 4.713572e-06, 
    4.699331e-06, 4.711903e-06, 4.69785e-06, 4.691269e-06, 4.764574e-06, 
    4.723356e-06, 4.785253e-06, 4.781819e-06, 4.753776e-06, 4.782206e-06, 
    4.507683e-06, 4.499863e-06, 4.472758e-06, 4.493964e-06, 4.455358e-06, 
    4.476952e-06, 4.489389e-06, 4.537505e-06, 4.548103e-06, 4.557942e-06, 
    4.577398e-06, 4.602418e-06, 4.646445e-06, 4.68489e-06, 4.720098e-06, 
    4.717515e-06, 4.718424e-06, 4.726304e-06, 4.706797e-06, 4.72951e-06, 
    4.733327e-06, 4.72335e-06, 4.781359e-06, 4.764757e-06, 4.781746e-06, 
    4.770933e-06, 4.502404e-06, 4.515568e-06, 4.508453e-06, 4.521838e-06, 
    4.512407e-06, 4.554405e-06, 4.567029e-06, 4.626284e-06, 4.601925e-06, 
    4.640715e-06, 4.605859e-06, 4.612028e-06, 4.641987e-06, 4.607739e-06, 
    4.682769e-06, 4.63185e-06, 4.72661e-06, 4.675571e-06, 4.729816e-06, 
    4.719946e-06, 4.736292e-06, 4.750952e-06, 4.769421e-06, 4.803576e-06, 
    4.795658e-06, 4.824276e-06, 4.535223e-06, 4.552353e-06, 4.550842e-06, 
    4.568794e-06, 4.582089e-06, 4.610959e-06, 4.657421e-06, 4.639926e-06, 
    4.672062e-06, 4.678524e-06, 4.62971e-06, 4.659658e-06, 4.563831e-06, 
    4.57926e-06, 4.57007e-06, 4.536574e-06, 4.643957e-06, 4.58872e-06, 
    4.690929e-06, 4.660847e-06, 4.748862e-06, 4.705008e-06, 4.791301e-06, 
    4.82839e-06, 4.863392e-06, 4.904435e-06, 4.561712e-06, 4.550059e-06, 
    4.57093e-06, 4.599875e-06, 4.626792e-06, 4.662681e-06, 4.666358e-06, 
    4.673097e-06, 4.690568e-06, 4.705279e-06, 4.67523e-06, 4.70897e-06, 
    4.582844e-06, 4.648764e-06, 4.545659e-06, 4.576608e-06, 4.598166e-06, 
    4.588702e-06, 4.637928e-06, 4.649562e-06, 4.696961e-06, 4.672433e-06, 
    4.819227e-06, 4.754054e-06, 4.935772e-06, 4.884715e-06, 4.545991e-06, 
    4.56167e-06, 4.616415e-06, 4.590334e-06, 4.665079e-06, 4.683554e-06, 
    4.698594e-06, 4.71785e-06, 4.71993e-06, 4.731356e-06, 4.712638e-06, 
    4.730616e-06, 4.662757e-06, 4.693032e-06, 4.610142e-06, 4.630263e-06, 
    4.621002e-06, 4.610853e-06, 4.642204e-06, 4.675703e-06, 4.676417e-06, 
    4.68718e-06, 4.717571e-06, 4.665383e-06, 4.82767e-06, 4.727184e-06, 
    4.578793e-06, 4.609108e-06, 4.613441e-06, 4.601684e-06, 4.681701e-06, 
    4.652643e-06, 4.731077e-06, 4.709826e-06, 4.744665e-06, 4.72734e-06, 
    4.724794e-06, 4.702584e-06, 4.688779e-06, 4.653974e-06, 4.625734e-06, 
    4.603388e-06, 4.60858e-06, 4.633139e-06, 4.677755e-06, 4.72012e-06, 
    4.710826e-06, 4.742014e-06, 4.659643e-06, 4.694113e-06, 4.680779e-06, 
    4.715578e-06, 4.639462e-06, 4.704256e-06, 4.62296e-06, 4.630064e-06, 
    4.652067e-06, 4.696456e-06, 4.706296e-06, 4.716816e-06, 4.710323e-06, 
    4.678889e-06, 4.673746e-06, 4.651531e-06, 4.645407e-06, 4.628517e-06, 
    4.614555e-06, 4.627312e-06, 4.640725e-06, 4.678901e-06, 4.713415e-06, 
    4.751162e-06, 4.760417e-06, 4.804717e-06, 4.768646e-06, 4.828233e-06, 
    4.77756e-06, 4.865411e-06, 4.708018e-06, 4.776067e-06, 4.653068e-06, 
    4.666255e-06, 4.69015e-06, 4.745134e-06, 4.715414e-06, 4.750177e-06, 
    4.673544e-06, 4.633989e-06, 4.623774e-06, 4.604746e-06, 4.624209e-06, 
    4.622625e-06, 4.641279e-06, 4.635281e-06, 4.680171e-06, 4.656035e-06, 
    4.72473e-06, 4.749902e-06, 4.821275e-06, 4.865243e-06, 4.91016e-06, 
    4.930043e-06, 4.936102e-06, 4.938635e-06,
  4.331469e-06, 4.372469e-06, 4.364484e-06, 4.397659e-06, 4.37924e-06, 
    4.400985e-06, 4.339765e-06, 4.374102e-06, 4.352167e-06, 4.335151e-06, 
    4.462383e-06, 4.399141e-06, 4.528512e-06, 4.48785e-06, 4.59032e-06, 
    4.522175e-06, 4.604118e-06, 4.588344e-06, 4.635889e-06, 4.622244e-06, 
    4.683315e-06, 4.642192e-06, 4.715116e-06, 4.673477e-06, 4.679981e-06, 
    4.640839e-06, 4.411831e-06, 4.454487e-06, 4.40931e-06, 4.415379e-06, 
    4.412655e-06, 4.379621e-06, 4.363021e-06, 4.328341e-06, 4.334627e-06, 
    4.360102e-06, 4.41811e-06, 4.398375e-06, 4.448184e-06, 4.447056e-06, 
    4.502814e-06, 4.477633e-06, 4.571838e-06, 4.544968e-06, 4.622813e-06, 
    4.603178e-06, 4.621891e-06, 4.616212e-06, 4.621965e-06, 4.593183e-06, 
    4.605504e-06, 4.580215e-06, 4.482345e-06, 4.511006e-06, 4.425782e-06, 
    4.374911e-06, 4.341269e-06, 4.317473e-06, 4.320834e-06, 4.327244e-06, 
    4.360251e-06, 4.39139e-06, 4.415191e-06, 4.431146e-06, 4.446894e-06, 
    4.49473e-06, 4.520138e-06, 4.577281e-06, 4.566941e-06, 4.584463e-06, 
    4.601226e-06, 4.629441e-06, 4.624791e-06, 4.637242e-06, 4.583997e-06, 
    4.619353e-06, 4.561056e-06, 4.576967e-06, 4.451191e-06, 4.403695e-06, 
    4.383589e-06, 4.366018e-06, 4.323419e-06, 4.352817e-06, 4.341216e-06, 
    4.368836e-06, 4.386429e-06, 4.377723e-06, 4.431583e-06, 4.410607e-06, 
    4.521647e-06, 4.473658e-06, 4.59927e-06, 4.569062e-06, 4.606524e-06, 
    4.587389e-06, 4.620199e-06, 4.590665e-06, 4.641879e-06, 4.653068e-06, 
    4.645421e-06, 4.674823e-06, 4.589032e-06, 4.621892e-06, 4.37748e-06, 
    4.378899e-06, 4.385514e-06, 4.356474e-06, 4.3547e-06, 4.328169e-06, 
    4.351771e-06, 4.361841e-06, 4.387449e-06, 4.402632e-06, 4.417087e-06, 
    4.448948e-06, 4.48466e-06, 4.534821e-06, 4.571018e-06, 4.595357e-06, 
    4.580425e-06, 4.593607e-06, 4.578872e-06, 4.571973e-06, 4.648874e-06, 
    4.60562e-06, 4.670589e-06, 4.666982e-06, 4.637539e-06, 4.667389e-06, 
    4.379896e-06, 4.37173e-06, 4.343439e-06, 4.365572e-06, 4.325285e-06, 
    4.347815e-06, 4.360796e-06, 4.411047e-06, 4.422122e-06, 4.432407e-06, 
    4.452749e-06, 4.478921e-06, 4.525008e-06, 4.565287e-06, 4.602202e-06, 
    4.599493e-06, 4.600447e-06, 4.608712e-06, 4.588253e-06, 4.612075e-06, 
    4.61608e-06, 4.605613e-06, 4.6665e-06, 4.649066e-06, 4.666906e-06, 
    4.655551e-06, 4.374383e-06, 4.388131e-06, 4.3807e-06, 4.394679e-06, 
    4.384829e-06, 4.42871e-06, 4.441907e-06, 4.503899e-06, 4.478406e-06, 
    4.519008e-06, 4.482521e-06, 4.488977e-06, 4.520341e-06, 4.484489e-06, 
    4.563065e-06, 4.509726e-06, 4.609034e-06, 4.555522e-06, 4.612397e-06, 
    4.602042e-06, 4.619191e-06, 4.634576e-06, 4.653963e-06, 4.689838e-06, 
    4.681518e-06, 4.711593e-06, 4.408662e-06, 4.426565e-06, 4.424985e-06, 
    4.443752e-06, 4.457655e-06, 4.487858e-06, 4.536504e-06, 4.518181e-06, 
    4.551843e-06, 4.558615e-06, 4.507484e-06, 4.538848e-06, 4.438563e-06, 
    4.454696e-06, 4.445086e-06, 4.410075e-06, 4.522403e-06, 4.464591e-06, 
    4.571617e-06, 4.540094e-06, 4.632381e-06, 4.586378e-06, 4.676942e-06, 
    4.715918e-06, 4.752727e-06, 4.795926e-06, 4.436347e-06, 4.424167e-06, 
    4.445985e-06, 4.47626e-06, 4.50443e-06, 4.542014e-06, 4.545866e-06, 
    4.552927e-06, 4.571238e-06, 4.586661e-06, 4.555163e-06, 4.590531e-06, 
    4.458446e-06, 4.527437e-06, 4.419568e-06, 4.451923e-06, 4.474472e-06, 
    4.464572e-06, 4.516089e-06, 4.528272e-06, 4.577941e-06, 4.552232e-06, 
    4.706286e-06, 4.637831e-06, 4.828933e-06, 4.775166e-06, 4.419915e-06, 
    4.436304e-06, 4.493569e-06, 4.466279e-06, 4.544527e-06, 4.563887e-06, 
    4.579652e-06, 4.599845e-06, 4.602026e-06, 4.614012e-06, 4.594378e-06, 
    4.613235e-06, 4.542094e-06, 4.573821e-06, 4.487003e-06, 4.508063e-06, 
    4.498369e-06, 4.487747e-06, 4.520566e-06, 4.555659e-06, 4.556407e-06, 
    4.567687e-06, 4.599554e-06, 4.544846e-06, 4.715163e-06, 4.609637e-06, 
    4.454208e-06, 4.485921e-06, 4.490455e-06, 4.478153e-06, 4.561944e-06, 
    4.5315e-06, 4.613719e-06, 4.591429e-06, 4.627977e-06, 4.609799e-06, 
    4.607128e-06, 4.583835e-06, 4.569363e-06, 4.532894e-06, 4.503322e-06, 
    4.479936e-06, 4.485368e-06, 4.511076e-06, 4.557809e-06, 4.602225e-06, 
    4.592478e-06, 4.625195e-06, 4.538832e-06, 4.574954e-06, 4.560978e-06, 
    4.597462e-06, 4.517696e-06, 4.58559e-06, 4.500419e-06, 4.507856e-06, 
    4.530896e-06, 4.577412e-06, 4.587727e-06, 4.598761e-06, 4.591951e-06, 
    4.558997e-06, 4.553608e-06, 4.530335e-06, 4.523921e-06, 4.506236e-06, 
    4.491621e-06, 4.504974e-06, 4.519018e-06, 4.55901e-06, 4.595193e-06, 
    4.634795e-06, 4.64451e-06, 4.691038e-06, 4.65315e-06, 4.715754e-06, 
    4.662512e-06, 4.754852e-06, 4.589534e-06, 4.660943e-06, 4.531945e-06, 
    4.545759e-06, 4.5708e-06, 4.628469e-06, 4.59729e-06, 4.633762e-06, 
    4.553396e-06, 4.511965e-06, 4.501271e-06, 4.481356e-06, 4.501726e-06, 
    4.500068e-06, 4.519597e-06, 4.513317e-06, 4.56034e-06, 4.535053e-06, 
    4.607061e-06, 4.633473e-06, 4.708438e-06, 4.754676e-06, 4.801953e-06, 
    4.822897e-06, 4.82928e-06, 4.831949e-06,
  4.36444e-06, 4.405082e-06, 4.397164e-06, 4.430068e-06, 4.411796e-06, 
    4.433368e-06, 4.372661e-06, 4.406701e-06, 4.384953e-06, 4.368088e-06, 
    4.494327e-06, 4.431539e-06, 4.560063e-06, 4.51963e-06, 4.621586e-06, 
    4.55376e-06, 4.635331e-06, 4.619616e-06, 4.666993e-06, 4.653392e-06, 
    4.714303e-06, 4.673278e-06, 4.746049e-06, 4.704484e-06, 4.710975e-06, 
    4.67193e-06, 4.44413e-06, 4.486484e-06, 4.441629e-06, 4.447652e-06, 
    4.444948e-06, 4.412175e-06, 4.395714e-06, 4.36134e-06, 4.367569e-06, 
    4.392819e-06, 4.450362e-06, 4.430779e-06, 4.48022e-06, 4.4791e-06, 
    4.534505e-06, 4.509477e-06, 4.603179e-06, 4.576434e-06, 4.653959e-06, 
    4.634393e-06, 4.65304e-06, 4.647381e-06, 4.653114e-06, 4.624437e-06, 
    4.636711e-06, 4.611521e-06, 4.514159e-06, 4.542651e-06, 4.457977e-06, 
    4.407505e-06, 4.374152e-06, 4.350573e-06, 4.353903e-06, 4.360253e-06, 
    4.392967e-06, 4.423848e-06, 4.447465e-06, 4.463303e-06, 4.478939e-06, 
    4.526471e-06, 4.551734e-06, 4.6086e-06, 4.598304e-06, 4.615752e-06, 
    4.632449e-06, 4.660566e-06, 4.655931e-06, 4.668344e-06, 4.615288e-06, 
    4.650512e-06, 4.592446e-06, 4.608286e-06, 4.48321e-06, 4.436056e-06, 
    4.416112e-06, 4.398686e-06, 4.356463e-06, 4.385598e-06, 4.3741e-06, 
    4.401478e-06, 4.418927e-06, 4.410292e-06, 4.463736e-06, 4.442916e-06, 
    4.553234e-06, 4.505527e-06, 4.6305e-06, 4.600416e-06, 4.637727e-06, 
    4.618666e-06, 4.651354e-06, 4.621929e-06, 4.672966e-06, 4.684124e-06, 
    4.676498e-06, 4.705827e-06, 4.620301e-06, 4.653041e-06, 4.410051e-06, 
    4.411459e-06, 4.418019e-06, 4.389223e-06, 4.387464e-06, 4.36117e-06, 
    4.384561e-06, 4.394544e-06, 4.419939e-06, 4.435002e-06, 4.449347e-06, 
    4.480979e-06, 4.51646e-06, 4.566338e-06, 4.602363e-06, 4.626602e-06, 
    4.611729e-06, 4.624859e-06, 4.610184e-06, 4.603314e-06, 4.679943e-06, 
    4.636826e-06, 4.701602e-06, 4.698004e-06, 4.668639e-06, 4.698409e-06, 
    4.412447e-06, 4.404349e-06, 4.376302e-06, 4.398242e-06, 4.358312e-06, 
    4.380639e-06, 4.393508e-06, 4.443354e-06, 4.454344e-06, 4.464554e-06, 
    4.484754e-06, 4.510756e-06, 4.556577e-06, 4.596659e-06, 4.633421e-06, 
    4.630721e-06, 4.631672e-06, 4.639907e-06, 4.619525e-06, 4.643258e-06, 
    4.647249e-06, 4.63682e-06, 4.697522e-06, 4.680133e-06, 4.697927e-06, 
    4.6866e-06, 4.40698e-06, 4.420615e-06, 4.413244e-06, 4.427111e-06, 
    4.417341e-06, 4.460885e-06, 4.473988e-06, 4.535586e-06, 4.510244e-06, 
    4.550609e-06, 4.514334e-06, 4.52075e-06, 4.551936e-06, 4.516289e-06, 
    4.594446e-06, 4.54138e-06, 4.640227e-06, 4.586939e-06, 4.643579e-06, 
    4.633262e-06, 4.650349e-06, 4.665685e-06, 4.685017e-06, 4.720812e-06, 
    4.712509e-06, 4.742531e-06, 4.440986e-06, 4.458755e-06, 4.457186e-06, 
    4.475819e-06, 4.489628e-06, 4.519638e-06, 4.568013e-06, 4.549786e-06, 
    4.583275e-06, 4.590016e-06, 4.539149e-06, 4.570345e-06, 4.470667e-06, 
    4.48669e-06, 4.477144e-06, 4.442387e-06, 4.553986e-06, 4.496518e-06, 
    4.60296e-06, 4.571584e-06, 4.663497e-06, 4.617659e-06, 4.707942e-06, 
    4.746852e-06, 4.783626e-06, 4.826826e-06, 4.468467e-06, 4.456374e-06, 
    4.478037e-06, 4.508112e-06, 4.536113e-06, 4.573495e-06, 4.577328e-06, 
    4.584355e-06, 4.602582e-06, 4.61794e-06, 4.586581e-06, 4.621795e-06, 
    4.490416e-06, 4.558993e-06, 4.451809e-06, 4.483936e-06, 4.506335e-06, 
    4.496499e-06, 4.547705e-06, 4.559823e-06, 4.609257e-06, 4.583663e-06, 
    4.737234e-06, 4.668932e-06, 4.859859e-06, 4.806061e-06, 4.452154e-06, 
    4.468423e-06, 4.525315e-06, 4.498195e-06, 4.575995e-06, 4.595264e-06, 
    4.61096e-06, 4.631073e-06, 4.633245e-06, 4.645189e-06, 4.625627e-06, 
    4.644414e-06, 4.573575e-06, 4.605154e-06, 4.518789e-06, 4.539725e-06, 
    4.530086e-06, 4.519527e-06, 4.552158e-06, 4.587075e-06, 4.587818e-06, 
    4.599048e-06, 4.630786e-06, 4.576312e-06, 4.746099e-06, 4.640832e-06, 
    4.486204e-06, 4.517714e-06, 4.52222e-06, 4.509992e-06, 4.59333e-06, 
    4.563034e-06, 4.644897e-06, 4.622689e-06, 4.659107e-06, 4.64099e-06, 
    4.638328e-06, 4.615126e-06, 4.600715e-06, 4.564421e-06, 4.535011e-06, 
    4.511764e-06, 4.517163e-06, 4.54272e-06, 4.589214e-06, 4.633444e-06, 
    4.623735e-06, 4.656333e-06, 4.570329e-06, 4.606283e-06, 4.592369e-06, 
    4.628698e-06, 4.549303e-06, 4.616877e-06, 4.532124e-06, 4.539518e-06, 
    4.562434e-06, 4.60873e-06, 4.619002e-06, 4.629993e-06, 4.623208e-06, 
    4.590397e-06, 4.585032e-06, 4.561875e-06, 4.555495e-06, 4.537907e-06, 
    4.523378e-06, 4.536653e-06, 4.550619e-06, 4.590409e-06, 4.626439e-06, 
    4.665904e-06, 4.675589e-06, 4.722011e-06, 4.684208e-06, 4.746691e-06, 
    4.693548e-06, 4.785753e-06, 4.620803e-06, 4.691981e-06, 4.563477e-06, 
    4.577221e-06, 4.602147e-06, 4.659599e-06, 4.628527e-06, 4.664875e-06, 
    4.584822e-06, 4.543606e-06, 4.532971e-06, 4.513176e-06, 4.533424e-06, 
    4.531775e-06, 4.551195e-06, 4.544949e-06, 4.591734e-06, 4.566569e-06, 
    4.638262e-06, 4.664586e-06, 4.739381e-06, 4.785575e-06, 4.832855e-06, 
    4.853816e-06, 4.860206e-06, 4.862879e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SNOW_SOURCES =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SOIL1C =
  5.777963, 5.777943, 5.777946, 5.77793, 5.777939, 5.777928, 5.777958, 
    5.777942, 5.777952, 5.777961, 5.777898, 5.777929, 5.777866, 5.777886, 
    5.777837, 5.77787, 5.77783, 5.777838, 5.777815, 5.777822, 5.777792, 
    5.777812, 5.777777, 5.777797, 5.777794, 5.777812, 5.777923, 5.777902, 
    5.777925, 5.777921, 5.777923, 5.777939, 5.777947, 5.777964, 5.777961, 
    5.777948, 5.77792, 5.77793, 5.777905, 5.777906, 5.777879, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.777831, 5.777822, 5.777824, 5.777822, 
    5.777835, 5.777829, 5.777842, 5.777889, 5.777875, 5.777916, 5.777941, 
    5.777958, 5.777969, 5.777968, 5.777965, 5.777948, 5.777933, 5.777922, 
    5.777914, 5.777906, 5.777883, 5.777871, 5.777843, 5.777848, 5.77784, 
    5.777832, 5.777818, 5.77782, 5.777814, 5.77784, 5.777823, 5.777851, 
    5.777843, 5.777904, 5.777927, 5.777937, 5.777946, 5.777966, 5.777952, 
    5.777958, 5.777944, 5.777936, 5.77794, 5.777914, 5.777924, 5.77787, 
    5.777893, 5.777833, 5.777847, 5.777829, 5.777838, 5.777822, 5.777836, 
    5.777812, 5.777807, 5.77781, 5.777796, 5.777837, 5.777822, 5.77794, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777953, 5.777948, 
    5.777935, 5.777928, 5.777921, 5.777905, 5.777888, 5.777864, 5.777846, 
    5.777834, 5.777842, 5.777835, 5.777842, 5.777845, 5.777809, 5.777829, 
    5.777798, 5.7778, 5.777814, 5.7778, 5.777939, 5.777943, 5.777957, 
    5.777946, 5.777966, 5.777955, 5.777948, 5.777924, 5.777918, 5.777913, 
    5.777903, 5.77789, 5.777868, 5.777849, 5.777831, 5.777832, 5.777832, 
    5.777828, 5.777838, 5.777826, 5.777824, 5.777829, 5.7778, 5.777809, 
    5.7778, 5.777805, 5.777942, 5.777935, 5.777938, 5.777932, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.777891, 5.777871, 5.777889, 5.777885, 
    5.77787, 5.777888, 5.77785, 5.777875, 5.777828, 5.777853, 5.777826, 
    5.777831, 5.777823, 5.777815, 5.777806, 5.777789, 5.777793, 5.777779, 
    5.777925, 5.777916, 5.777917, 5.777907, 5.777901, 5.777886, 5.777863, 
    5.777872, 5.777855, 5.777852, 5.777876, 5.777862, 5.77791, 5.777902, 
    5.777907, 5.777924, 5.777869, 5.777897, 5.777846, 5.777861, 5.777816, 
    5.777839, 5.777795, 5.777777, 5.77776, 5.777739, 5.777911, 5.777917, 
    5.777906, 5.777892, 5.777878, 5.77786, 5.777858, 5.777854, 5.777846, 
    5.777838, 5.777853, 5.777837, 5.7779, 5.777867, 5.777919, 5.777904, 
    5.777893, 5.777897, 5.777873, 5.777866, 5.777843, 5.777855, 5.777781, 
    5.777814, 5.777724, 5.777749, 5.777919, 5.777911, 5.777884, 5.777896, 
    5.777859, 5.777849, 5.777842, 5.777832, 5.777831, 5.777825, 5.777835, 
    5.777826, 5.77786, 5.777844, 5.777886, 5.777876, 5.777881, 5.777886, 
    5.77787, 5.777853, 5.777853, 5.777848, 5.777832, 5.777859, 5.777777, 
    5.777827, 5.777903, 5.777887, 5.777885, 5.777891, 5.77785, 5.777865, 
    5.777825, 5.777836, 5.777819, 5.777827, 5.777829, 5.77784, 5.777847, 
    5.777864, 5.777879, 5.77789, 5.777887, 5.777875, 5.777852, 5.777831, 
    5.777836, 5.77782, 5.777862, 5.777844, 5.777851, 5.777833, 5.777872, 
    5.777839, 5.77788, 5.777876, 5.777865, 5.777843, 5.777838, 5.777833, 
    5.777836, 5.777852, 5.777854, 5.777865, 5.777869, 5.777877, 5.777884, 
    5.777878, 5.777871, 5.777852, 5.777834, 5.777815, 5.777811, 5.777789, 
    5.777807, 5.777777, 5.777802, 5.777759, 5.777837, 5.777803, 5.777865, 
    5.777858, 5.777846, 5.777818, 5.777833, 5.777816, 5.777854, 5.777874, 
    5.77788, 5.777889, 5.777879, 5.77788, 5.777871, 5.777874, 5.777851, 
    5.777864, 5.777829, 5.777816, 5.777781, 5.777759, 5.777736, 5.777726, 
    5.777723, 5.777722 ;

 SOIL1C_TO_SOIL2C =
  3.180121e-08, 3.194099e-08, 3.191381e-08, 3.202655e-08, 3.196401e-08, 
    3.203784e-08, 3.182955e-08, 3.194654e-08, 3.187186e-08, 3.181379e-08, 
    3.224534e-08, 3.203158e-08, 3.246734e-08, 3.233103e-08, 3.267344e-08, 
    3.244613e-08, 3.271928e-08, 3.266688e-08, 3.282457e-08, 3.277939e-08, 
    3.298108e-08, 3.284542e-08, 3.308563e-08, 3.294868e-08, 3.297011e-08, 
    3.284094e-08, 3.20746e-08, 3.221872e-08, 3.206605e-08, 3.208661e-08, 
    3.207738e-08, 3.196531e-08, 3.190883e-08, 3.179053e-08, 3.1812e-08, 
    3.189889e-08, 3.209585e-08, 3.202899e-08, 3.219749e-08, 3.219368e-08, 
    3.238127e-08, 3.229669e-08, 3.261196e-08, 3.252235e-08, 3.278128e-08, 
    3.271616e-08, 3.277822e-08, 3.27594e-08, 3.277847e-08, 3.268297e-08, 
    3.272389e-08, 3.263985e-08, 3.231253e-08, 3.240873e-08, 3.212181e-08, 
    3.194928e-08, 3.183468e-08, 3.175336e-08, 3.176486e-08, 3.178677e-08, 
    3.18994e-08, 3.200528e-08, 3.208597e-08, 3.213995e-08, 3.219314e-08, 
    3.235412e-08, 3.243932e-08, 3.263008e-08, 3.259565e-08, 3.265397e-08, 
    3.270969e-08, 3.280323e-08, 3.278783e-08, 3.282904e-08, 3.265243e-08, 
    3.276981e-08, 3.257604e-08, 3.262904e-08, 3.220761e-08, 3.204703e-08, 
    3.197878e-08, 3.191904e-08, 3.177369e-08, 3.187407e-08, 3.18345e-08, 
    3.192863e-08, 3.198844e-08, 3.195886e-08, 3.214143e-08, 3.207045e-08, 
    3.244437e-08, 3.228331e-08, 3.270319e-08, 3.260272e-08, 3.272727e-08, 
    3.266371e-08, 3.277261e-08, 3.26746e-08, 3.284438e-08, 3.288135e-08, 
    3.285609e-08, 3.295312e-08, 3.266917e-08, 3.277822e-08, 3.195803e-08, 
    3.196286e-08, 3.198533e-08, 3.188653e-08, 3.188049e-08, 3.178994e-08, 
    3.187051e-08, 3.190482e-08, 3.199191e-08, 3.204342e-08, 3.209239e-08, 
    3.220006e-08, 3.232031e-08, 3.248844e-08, 3.260923e-08, 3.26902e-08, 
    3.264055e-08, 3.268438e-08, 3.263538e-08, 3.261241e-08, 3.28675e-08, 
    3.272427e-08, 3.293917e-08, 3.292728e-08, 3.283002e-08, 3.292861e-08, 
    3.196624e-08, 3.193848e-08, 3.184208e-08, 3.191752e-08, 3.178008e-08, 
    3.185701e-08, 3.190125e-08, 3.207194e-08, 3.210943e-08, 3.214421e-08, 
    3.221288e-08, 3.230102e-08, 3.245562e-08, 3.259014e-08, 3.271293e-08, 
    3.270393e-08, 3.27071e-08, 3.273453e-08, 3.266658e-08, 3.274569e-08, 
    3.275896e-08, 3.272425e-08, 3.292568e-08, 3.286814e-08, 3.292702e-08, 
    3.288955e-08, 3.19475e-08, 3.199422e-08, 3.196898e-08, 3.201645e-08, 
    3.198301e-08, 3.213171e-08, 3.217629e-08, 3.23849e-08, 3.229928e-08, 
    3.243554e-08, 3.231312e-08, 3.233481e-08, 3.243998e-08, 3.231974e-08, 
    3.258272e-08, 3.240443e-08, 3.27356e-08, 3.255757e-08, 3.274675e-08, 
    3.27124e-08, 3.276928e-08, 3.282022e-08, 3.288431e-08, 3.300256e-08, 
    3.297518e-08, 3.307407e-08, 3.206386e-08, 3.212446e-08, 3.211912e-08, 
    3.218253e-08, 3.222942e-08, 3.233106e-08, 3.249407e-08, 3.243277e-08, 
    3.254531e-08, 3.25679e-08, 3.239693e-08, 3.250191e-08, 3.216501e-08, 
    3.221944e-08, 3.218703e-08, 3.206864e-08, 3.24469e-08, 3.225279e-08, 
    3.261123e-08, 3.250607e-08, 3.281296e-08, 3.266034e-08, 3.296011e-08, 
    3.308825e-08, 3.320885e-08, 3.334979e-08, 3.215752e-08, 3.211635e-08, 
    3.219007e-08, 3.229206e-08, 3.238669e-08, 3.251249e-08, 3.252536e-08, 
    3.254892e-08, 3.260996e-08, 3.266129e-08, 3.255638e-08, 3.267415e-08, 
    3.223207e-08, 3.246375e-08, 3.210079e-08, 3.221009e-08, 3.228605e-08, 
    3.225272e-08, 3.242577e-08, 3.246655e-08, 3.263228e-08, 3.254661e-08, 
    3.305663e-08, 3.283099e-08, 3.345709e-08, 3.328213e-08, 3.210197e-08, 
    3.215738e-08, 3.235024e-08, 3.225848e-08, 3.252088e-08, 3.258547e-08, 
    3.263797e-08, 3.27051e-08, 3.271234e-08, 3.275211e-08, 3.268694e-08, 
    3.274953e-08, 3.251276e-08, 3.261857e-08, 3.232819e-08, 3.239887e-08, 
    3.236635e-08, 3.233069e-08, 3.244076e-08, 3.255803e-08, 3.256053e-08, 
    3.259813e-08, 3.27041e-08, 3.252195e-08, 3.308576e-08, 3.273757e-08, 
    3.221781e-08, 3.232454e-08, 3.233978e-08, 3.229844e-08, 3.2579e-08, 
    3.247734e-08, 3.275114e-08, 3.267714e-08, 3.279838e-08, 3.273814e-08, 
    3.272927e-08, 3.265189e-08, 3.260372e-08, 3.2482e-08, 3.238297e-08, 
    3.230443e-08, 3.23227e-08, 3.240896e-08, 3.25652e-08, 3.2713e-08, 
    3.268062e-08, 3.278917e-08, 3.250186e-08, 3.262234e-08, 3.257577e-08, 
    3.269718e-08, 3.243115e-08, 3.265771e-08, 3.237323e-08, 3.239818e-08, 
    3.247532e-08, 3.263051e-08, 3.266484e-08, 3.270149e-08, 3.267887e-08, 
    3.256917e-08, 3.255119e-08, 3.247345e-08, 3.245199e-08, 3.239274e-08, 
    3.23437e-08, 3.238851e-08, 3.243557e-08, 3.256921e-08, 3.268964e-08, 
    3.282095e-08, 3.285308e-08, 3.30065e-08, 3.288161e-08, 3.30877e-08, 
    3.29125e-08, 3.321577e-08, 3.267083e-08, 3.290733e-08, 3.247883e-08, 
    3.2525e-08, 3.26085e-08, 3.28e-08, 3.269661e-08, 3.281752e-08, 
    3.255049e-08, 3.241194e-08, 3.237609e-08, 3.230921e-08, 3.237762e-08, 
    3.237206e-08, 3.243752e-08, 3.241648e-08, 3.257365e-08, 3.248923e-08, 
    3.272905e-08, 3.281657e-08, 3.306371e-08, 3.321521e-08, 3.336942e-08, 
    3.34375e-08, 3.345822e-08, 3.346688e-08 ;

 SOIL1C_TO_SOIL3C =
  3.771725e-10, 3.788308e-10, 3.785084e-10, 3.79846e-10, 3.79104e-10, 
    3.799799e-10, 3.775087e-10, 3.788967e-10, 3.780106e-10, 3.773217e-10, 
    3.824418e-10, 3.799057e-10, 3.85076e-10, 3.834586e-10, 3.875214e-10, 
    3.848243e-10, 3.880652e-10, 3.874436e-10, 3.893146e-10, 3.887785e-10, 
    3.911717e-10, 3.895619e-10, 3.924122e-10, 3.907873e-10, 3.910415e-10, 
    3.895088e-10, 3.80416e-10, 3.821261e-10, 3.803147e-10, 3.805586e-10, 
    3.804491e-10, 3.791193e-10, 3.784492e-10, 3.770457e-10, 3.773005e-10, 
    3.783313e-10, 3.806682e-10, 3.798749e-10, 3.818741e-10, 3.81829e-10, 
    3.840546e-10, 3.830511e-10, 3.867919e-10, 3.857287e-10, 3.888009e-10, 
    3.880283e-10, 3.887646e-10, 3.885414e-10, 3.887675e-10, 3.876344e-10, 
    3.881199e-10, 3.871228e-10, 3.832391e-10, 3.843805e-10, 3.809762e-10, 
    3.789293e-10, 3.775695e-10, 3.766047e-10, 3.767411e-10, 3.770011e-10, 
    3.783374e-10, 3.795937e-10, 3.805511e-10, 3.811915e-10, 3.818225e-10, 
    3.837326e-10, 3.847434e-10, 3.870069e-10, 3.865984e-10, 3.872904e-10, 
    3.879514e-10, 3.890613e-10, 3.888787e-10, 3.893676e-10, 3.872721e-10, 
    3.886648e-10, 3.863657e-10, 3.869945e-10, 3.819942e-10, 3.800889e-10, 
    3.792792e-10, 3.785704e-10, 3.76846e-10, 3.780369e-10, 3.775674e-10, 
    3.786842e-10, 3.793938e-10, 3.790429e-10, 3.81209e-10, 3.803669e-10, 
    3.848034e-10, 3.828924e-10, 3.878743e-10, 3.866822e-10, 3.881601e-10, 
    3.874059e-10, 3.886981e-10, 3.875352e-10, 3.895496e-10, 3.899883e-10, 
    3.896885e-10, 3.908399e-10, 3.874707e-10, 3.887647e-10, 3.79033e-10, 
    3.790903e-10, 3.79357e-10, 3.781847e-10, 3.78113e-10, 3.770387e-10, 
    3.779946e-10, 3.784017e-10, 3.79435e-10, 3.800462e-10, 3.806272e-10, 
    3.819047e-10, 3.833314e-10, 3.853263e-10, 3.867595e-10, 3.877202e-10, 
    3.871311e-10, 3.876512e-10, 3.870698e-10, 3.867973e-10, 3.898239e-10, 
    3.881244e-10, 3.906744e-10, 3.905332e-10, 3.893793e-10, 3.905491e-10, 
    3.791305e-10, 3.78801e-10, 3.776574e-10, 3.785524e-10, 3.769217e-10, 
    3.778345e-10, 3.783594e-10, 3.803845e-10, 3.808294e-10, 3.81242e-10, 
    3.820568e-10, 3.831025e-10, 3.849369e-10, 3.865329e-10, 3.879899e-10, 
    3.878831e-10, 3.879207e-10, 3.882462e-10, 3.8744e-10, 3.883786e-10, 
    3.885361e-10, 3.881242e-10, 3.905143e-10, 3.898315e-10, 3.905302e-10, 
    3.900856e-10, 3.789081e-10, 3.794624e-10, 3.791629e-10, 3.797261e-10, 
    3.793293e-10, 3.810937e-10, 3.816227e-10, 3.840978e-10, 3.830819e-10, 
    3.846986e-10, 3.832462e-10, 3.835035e-10, 3.847514e-10, 3.833246e-10, 
    3.86445e-10, 3.843295e-10, 3.882589e-10, 3.861465e-10, 3.883912e-10, 
    3.879836e-10, 3.886585e-10, 3.89263e-10, 3.900234e-10, 3.914266e-10, 
    3.911016e-10, 3.92275e-10, 3.802887e-10, 3.810076e-10, 3.809443e-10, 
    3.816966e-10, 3.822531e-10, 3.83459e-10, 3.853931e-10, 3.846658e-10, 
    3.86001e-10, 3.862691e-10, 3.842405e-10, 3.854861e-10, 3.814888e-10, 
    3.821346e-10, 3.8175e-10, 3.803454e-10, 3.848334e-10, 3.825302e-10, 
    3.867832e-10, 3.855355e-10, 3.891768e-10, 3.873659e-10, 3.909228e-10, 
    3.924434e-10, 3.938743e-10, 3.955467e-10, 3.814e-10, 3.809115e-10, 
    3.817861e-10, 3.829962e-10, 3.84119e-10, 3.856116e-10, 3.857643e-10, 
    3.860439e-10, 3.867682e-10, 3.873772e-10, 3.861324e-10, 3.875299e-10, 
    3.822845e-10, 3.850333e-10, 3.807268e-10, 3.820237e-10, 3.829249e-10, 
    3.825295e-10, 3.845826e-10, 3.850666e-10, 3.870329e-10, 3.860164e-10, 
    3.920681e-10, 3.893907e-10, 3.968199e-10, 3.947438e-10, 3.807408e-10, 
    3.813983e-10, 3.836865e-10, 3.825978e-10, 3.857112e-10, 3.864776e-10, 
    3.871006e-10, 3.87897e-10, 3.879829e-10, 3.884548e-10, 3.876816e-10, 
    3.884242e-10, 3.856148e-10, 3.868703e-10, 3.834249e-10, 3.842635e-10, 
    3.838777e-10, 3.834545e-10, 3.847606e-10, 3.86152e-10, 3.861817e-10, 
    3.866278e-10, 3.878852e-10, 3.857238e-10, 3.924137e-10, 3.882824e-10, 
    3.821152e-10, 3.833816e-10, 3.835625e-10, 3.830719e-10, 3.864008e-10, 
    3.851946e-10, 3.884433e-10, 3.875653e-10, 3.890039e-10, 3.88289e-10, 
    3.881838e-10, 3.872657e-10, 3.866941e-10, 3.852499e-10, 3.840749e-10, 
    3.83143e-10, 3.833597e-10, 3.843833e-10, 3.862371e-10, 3.879907e-10, 
    3.876066e-10, 3.888945e-10, 3.854855e-10, 3.86915e-10, 3.863625e-10, 
    3.878031e-10, 3.846465e-10, 3.873347e-10, 3.839594e-10, 3.842553e-10, 
    3.851707e-10, 3.87012e-10, 3.874193e-10, 3.878542e-10, 3.875858e-10, 
    3.862841e-10, 3.860709e-10, 3.851484e-10, 3.848938e-10, 3.841908e-10, 
    3.83609e-10, 3.841406e-10, 3.84699e-10, 3.862847e-10, 3.877136e-10, 
    3.892716e-10, 3.896528e-10, 3.914732e-10, 3.899914e-10, 3.924367e-10, 
    3.903579e-10, 3.939565e-10, 3.874903e-10, 3.902966e-10, 3.852123e-10, 
    3.857601e-10, 3.867508e-10, 3.890231e-10, 3.877963e-10, 3.89231e-10, 
    3.860625e-10, 3.844186e-10, 3.839933e-10, 3.831997e-10, 3.840114e-10, 
    3.839454e-10, 3.847221e-10, 3.844725e-10, 3.863373e-10, 3.853356e-10, 
    3.881812e-10, 3.892196e-10, 3.921521e-10, 3.939498e-10, 3.957796e-10, 
    3.965875e-10, 3.968333e-10, 3.969361e-10 ;

 SOIL1C_vr =
  19.97935, 19.9793, 19.97931, 19.97927, 19.97929, 19.97926, 19.97934, 
    19.9793, 19.97933, 19.97935, 19.97918, 19.97926, 19.9791, 19.97915, 
    19.97902, 19.9791, 19.979, 19.97902, 19.97896, 19.97898, 19.9789, 
    19.97895, 19.97886, 19.97891, 19.9789, 19.97895, 19.97925, 19.97919, 
    19.97925, 19.97924, 19.97925, 19.97929, 19.97931, 19.97936, 19.97935, 
    19.97931, 19.97924, 19.97927, 19.9792, 19.9792, 19.97913, 19.97916, 
    19.97904, 19.97907, 19.97898, 19.979, 19.97898, 19.97898, 19.97898, 
    19.97901, 19.979, 19.97903, 19.97916, 19.97912, 19.97923, 19.9793, 
    19.97934, 19.97937, 19.97937, 19.97936, 19.97931, 19.97927, 19.97924, 
    19.97922, 19.9792, 19.97914, 19.97911, 19.97903, 19.97905, 19.97902, 
    19.979, 19.97897, 19.97897, 19.97896, 19.97902, 19.97898, 19.97905, 
    19.97903, 19.9792, 19.97926, 19.97928, 19.97931, 19.97936, 19.97932, 
    19.97934, 19.9793, 19.97928, 19.97929, 19.97922, 19.97925, 19.9791, 
    19.97917, 19.97901, 19.97904, 19.979, 19.97902, 19.97898, 19.97902, 
    19.97895, 19.97894, 19.97895, 19.97891, 19.97902, 19.97898, 19.97929, 
    19.97929, 19.97928, 19.97932, 19.97932, 19.97936, 19.97933, 19.97931, 
    19.97928, 19.97926, 19.97924, 19.9792, 19.97915, 19.97909, 19.97904, 
    19.97901, 19.97903, 19.97901, 19.97903, 19.97904, 19.97894, 19.979, 
    19.97891, 19.97892, 19.97896, 19.97892, 19.97929, 19.9793, 19.97934, 
    19.97931, 19.97936, 19.97933, 19.97931, 19.97925, 19.97923, 19.97922, 
    19.97919, 19.97916, 19.9791, 19.97905, 19.979, 19.97901, 19.979, 
    19.97899, 19.97902, 19.97899, 19.97898, 19.979, 19.97892, 19.97894, 
    19.97892, 19.97893, 19.9793, 19.97928, 19.97929, 19.97927, 19.97928, 
    19.97923, 19.97921, 19.97913, 19.97916, 19.97911, 19.97916, 19.97915, 
    19.97911, 19.97915, 19.97905, 19.97912, 19.97899, 19.97906, 19.97899, 
    19.979, 19.97898, 19.97896, 19.97894, 19.97889, 19.9789, 19.97886, 
    19.97925, 19.97923, 19.97923, 19.97921, 19.97919, 19.97915, 19.97909, 
    19.97911, 19.97907, 19.97906, 19.97912, 19.97908, 19.97921, 19.97919, 
    19.9792, 19.97925, 19.9791, 19.97918, 19.97904, 19.97908, 19.97896, 
    19.97902, 19.97891, 19.97886, 19.97881, 19.97876, 19.97922, 19.97923, 
    19.9792, 19.97916, 19.97913, 19.97908, 19.97907, 19.97906, 19.97904, 
    19.97902, 19.97906, 19.97902, 19.97919, 19.9791, 19.97924, 19.97919, 
    19.97917, 19.97918, 19.97911, 19.9791, 19.97903, 19.97906, 19.97887, 
    19.97896, 19.97872, 19.97878, 19.97924, 19.97922, 19.97914, 19.97918, 
    19.97908, 19.97905, 19.97903, 19.979, 19.979, 19.97899, 19.97901, 
    19.97899, 19.97908, 19.97904, 19.97915, 19.97912, 19.97914, 19.97915, 
    19.97911, 19.97906, 19.97906, 19.97905, 19.97901, 19.97907, 19.97886, 
    19.97899, 19.97919, 19.97915, 19.97915, 19.97916, 19.97905, 19.97909, 
    19.97899, 19.97902, 19.97897, 19.97899, 19.979, 19.97902, 19.97904, 
    19.97909, 19.97913, 19.97916, 19.97915, 19.97912, 19.97906, 19.979, 
    19.97901, 19.97897, 19.97908, 19.97904, 19.97906, 19.97901, 19.97911, 
    19.97902, 19.97913, 19.97912, 19.97909, 19.97903, 19.97902, 19.97901, 
    19.97902, 19.97906, 19.97906, 19.97909, 19.9791, 19.97912, 19.97914, 
    19.97913, 19.97911, 19.97906, 19.97901, 19.97896, 19.97895, 19.97889, 
    19.97894, 19.97886, 19.97893, 19.97881, 19.97902, 19.97893, 19.97909, 
    19.97907, 19.97904, 19.97897, 19.97901, 19.97896, 19.97906, 19.97912, 
    19.97913, 19.97916, 19.97913, 19.97913, 19.97911, 19.97912, 19.97906, 
    19.97909, 19.979, 19.97896, 19.97887, 19.97881, 19.97875, 19.97873, 
    19.97872, 19.97871,
  19.98101, 19.98094, 19.98095, 19.98089, 19.98092, 19.98089, 19.98099, 
    19.98093, 19.98097, 19.981, 19.98078, 19.98089, 19.98067, 19.98074, 
    19.98057, 19.98068, 19.98054, 19.98057, 19.98049, 19.98051, 19.98041, 
    19.98048, 19.98036, 19.98043, 19.98042, 19.98048, 19.98087, 19.98079, 
    19.98087, 19.98086, 19.98087, 19.98092, 19.98095, 19.98101, 19.981, 
    19.98096, 19.98086, 19.98089, 19.98081, 19.98081, 19.98071, 19.98076, 
    19.9806, 19.98064, 19.98051, 19.98054, 19.98051, 19.98052, 19.98051, 
    19.98056, 19.98054, 19.98058, 19.98075, 19.9807, 19.98084, 19.98093, 
    19.98099, 19.98103, 19.98103, 19.98101, 19.98096, 19.9809, 19.98086, 
    19.98083, 19.98081, 19.98073, 19.98068, 19.98059, 19.9806, 19.98058, 
    19.98055, 19.9805, 19.98051, 19.98049, 19.98058, 19.98052, 19.98061, 
    19.98059, 19.9808, 19.98088, 19.98092, 19.98095, 19.98102, 19.98097, 
    19.98099, 19.98094, 19.98091, 19.98093, 19.98083, 19.98087, 19.98068, 
    19.98076, 19.98055, 19.9806, 19.98054, 19.98057, 19.98051, 19.98056, 
    19.98048, 19.98046, 19.98047, 19.98042, 19.98057, 19.98051, 19.98093, 
    19.98092, 19.98091, 19.98096, 19.98097, 19.98101, 19.98097, 19.98096, 
    19.98091, 19.98088, 19.98086, 19.9808, 19.98074, 19.98066, 19.9806, 
    19.98056, 19.98058, 19.98056, 19.98059, 19.9806, 19.98047, 19.98054, 
    19.98043, 19.98044, 19.98049, 19.98044, 19.98092, 19.98094, 19.98099, 
    19.98095, 19.98102, 19.98098, 19.98096, 19.98087, 19.98085, 19.98083, 
    19.9808, 19.98075, 19.98067, 19.98061, 19.98055, 19.98055, 19.98055, 
    19.98053, 19.98057, 19.98053, 19.98052, 19.98054, 19.98044, 19.98047, 
    19.98044, 19.98046, 19.98093, 19.98091, 19.98092, 19.9809, 19.98092, 
    19.98084, 19.98082, 19.98071, 19.98075, 19.98069, 19.98075, 19.98074, 
    19.98068, 19.98074, 19.98061, 19.9807, 19.98053, 19.98062, 19.98053, 
    19.98055, 19.98052, 19.98049, 19.98046, 19.9804, 19.98041, 19.98036, 
    19.98087, 19.98084, 19.98085, 19.98081, 19.98079, 19.98074, 19.98066, 
    19.98069, 19.98063, 19.98062, 19.98071, 19.98065, 19.98082, 19.98079, 
    19.98081, 19.98087, 19.98068, 19.98078, 19.9806, 19.98065, 19.9805, 
    19.98057, 19.98042, 19.98036, 19.9803, 19.98022, 19.98083, 19.98085, 
    19.98081, 19.98076, 19.98071, 19.98065, 19.98064, 19.98063, 19.9806, 
    19.98057, 19.98063, 19.98056, 19.98079, 19.98067, 19.98086, 19.9808, 
    19.98076, 19.98078, 19.98069, 19.98067, 19.98059, 19.98063, 19.98037, 
    19.98049, 19.98017, 19.98026, 19.98085, 19.98083, 19.98073, 19.98078, 
    19.98064, 19.98061, 19.98058, 19.98055, 19.98055, 19.98053, 19.98056, 
    19.98053, 19.98065, 19.98059, 19.98074, 19.9807, 19.98072, 19.98074, 
    19.98068, 19.98062, 19.98062, 19.9806, 19.98055, 19.98064, 19.98036, 
    19.98053, 19.9808, 19.98074, 19.98073, 19.98075, 19.98061, 19.98067, 
    19.98053, 19.98056, 19.9805, 19.98053, 19.98054, 19.98058, 19.9806, 
    19.98066, 19.98071, 19.98075, 19.98074, 19.9807, 19.98062, 19.98055, 
    19.98056, 19.98051, 19.98065, 19.98059, 19.98062, 19.98055, 19.98069, 
    19.98057, 19.98072, 19.98071, 19.98067, 19.98059, 19.98057, 19.98055, 
    19.98056, 19.98062, 19.98063, 19.98067, 19.98068, 19.98071, 19.98073, 
    19.98071, 19.98069, 19.98062, 19.98056, 19.98049, 19.98047, 19.9804, 
    19.98046, 19.98036, 19.98044, 19.98029, 19.98057, 19.98045, 19.98066, 
    19.98064, 19.9806, 19.9805, 19.98055, 19.98049, 19.98063, 19.9807, 
    19.98071, 19.98075, 19.98071, 19.98072, 19.98068, 19.9807, 19.98062, 
    19.98066, 19.98054, 19.98049, 19.98037, 19.98029, 19.98022, 19.98018, 
    19.98017, 19.98017,
  19.98273, 19.98265, 19.98267, 19.98261, 19.98264, 19.9826, 19.98271, 
    19.98265, 19.98269, 19.98272, 19.98249, 19.9826, 19.98237, 19.98244, 
    19.98226, 19.98238, 19.98223, 19.98226, 19.98217, 19.9822, 19.98209, 
    19.98216, 19.98203, 19.98211, 19.9821, 19.98217, 19.98258, 19.9825, 
    19.98258, 19.98257, 19.98258, 19.98264, 19.98267, 19.98273, 19.98272, 
    19.98268, 19.98257, 19.9826, 19.98251, 19.98252, 19.98241, 19.98246, 
    19.98229, 19.98234, 19.9822, 19.98223, 19.9822, 19.98221, 19.9822, 
    19.98225, 19.98223, 19.98228, 19.98245, 19.9824, 19.98255, 19.98265, 
    19.98271, 19.98275, 19.98275, 19.98274, 19.98268, 19.98262, 19.98257, 
    19.98254, 19.98252, 19.98243, 19.98238, 19.98228, 19.9823, 19.98227, 
    19.98224, 19.98219, 19.98219, 19.98217, 19.98227, 19.9822, 19.98231, 
    19.98228, 19.98251, 19.9826, 19.98263, 19.98266, 19.98274, 19.98269, 
    19.98271, 19.98266, 19.98263, 19.98264, 19.98254, 19.98258, 19.98238, 
    19.98247, 19.98224, 19.98229, 19.98223, 19.98226, 19.9822, 19.98226, 
    19.98216, 19.98214, 19.98216, 19.98211, 19.98226, 19.9822, 19.98264, 
    19.98264, 19.98263, 19.98268, 19.98269, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.9826, 19.98257, 19.98251, 19.98245, 19.98236, 19.98229, 
    19.98225, 19.98227, 19.98225, 19.98228, 19.98229, 19.98215, 19.98223, 
    19.98211, 19.98212, 19.98217, 19.98212, 19.98264, 19.98265, 19.98271, 
    19.98266, 19.98274, 19.9827, 19.98267, 19.98258, 19.98256, 19.98254, 
    19.98251, 19.98246, 19.98237, 19.9823, 19.98223, 19.98224, 19.98224, 
    19.98222, 19.98226, 19.98222, 19.98221, 19.98223, 19.98212, 19.98215, 
    19.98212, 19.98214, 19.98265, 19.98262, 19.98264, 19.98261, 19.98263, 
    19.98255, 19.98252, 19.98241, 19.98246, 19.98238, 19.98245, 19.98244, 
    19.98238, 19.98245, 19.98231, 19.9824, 19.98222, 19.98232, 19.98222, 
    19.98223, 19.9822, 19.98218, 19.98214, 19.98208, 19.98209, 19.98204, 
    19.98259, 19.98255, 19.98256, 19.98252, 19.9825, 19.98244, 19.98235, 
    19.98239, 19.98232, 19.98231, 19.9824, 19.98235, 19.98253, 19.9825, 
    19.98252, 19.98258, 19.98238, 19.98248, 19.98229, 19.98235, 19.98218, 
    19.98226, 19.9821, 19.98203, 19.98197, 19.98189, 19.98253, 19.98256, 
    19.98252, 19.98246, 19.98241, 19.98234, 19.98234, 19.98232, 19.98229, 
    19.98226, 19.98232, 19.98226, 19.98249, 19.98237, 19.98256, 19.98251, 
    19.98247, 19.98248, 19.98239, 19.98237, 19.98228, 19.98232, 19.98205, 
    19.98217, 19.98183, 19.98193, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98234, 19.9823, 19.98228, 19.98224, 19.98223, 19.98221, 19.98225, 
    19.98222, 19.98234, 19.98229, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98232, 19.98232, 19.9823, 19.98224, 19.98234, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98244, 19.98246, 19.98231, 19.98236, 
    19.98221, 19.98225, 19.98219, 19.98222, 19.98223, 19.98227, 19.98229, 
    19.98236, 19.98241, 19.98246, 19.98244, 19.9824, 19.98232, 19.98223, 
    19.98225, 19.98219, 19.98235, 19.98228, 19.98231, 19.98224, 19.98239, 
    19.98227, 19.98242, 19.9824, 19.98236, 19.98228, 19.98226, 19.98224, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98238, 19.98241, 19.98243, 
    19.98241, 19.98238, 19.98231, 19.98225, 19.98218, 19.98216, 19.98208, 
    19.98214, 19.98203, 19.98213, 19.98196, 19.98226, 19.98213, 19.98236, 
    19.98234, 19.98229, 19.98219, 19.98224, 19.98218, 19.98232, 19.9824, 
    19.98242, 19.98245, 19.98242, 19.98242, 19.98238, 19.9824, 19.98231, 
    19.98236, 19.98223, 19.98218, 19.98205, 19.98196, 19.98188, 19.98184, 
    19.98183, 19.98183,
  19.9841, 19.98403, 19.98404, 19.98398, 19.98401, 19.98397, 19.98409, 
    19.98402, 19.98406, 19.9841, 19.98386, 19.98398, 19.98375, 19.98382, 
    19.98363, 19.98376, 19.98361, 19.98364, 19.98355, 19.98358, 19.98347, 
    19.98354, 19.98341, 19.98349, 19.98347, 19.98355, 19.98396, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98405, 19.98411, 19.9841, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98384, 
    19.98367, 19.98372, 19.98358, 19.98361, 19.98358, 19.98359, 19.98358, 
    19.98363, 19.98361, 19.98365, 19.98383, 19.98378, 19.98393, 19.98402, 
    19.98409, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98366, 19.98368, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98365, 19.98358, 19.98369, 
    19.98366, 19.98388, 19.98397, 19.98401, 19.98404, 19.98412, 19.98406, 
    19.98409, 19.98403, 19.984, 19.98402, 19.98392, 19.98396, 19.98376, 
    19.98384, 19.98362, 19.98367, 19.98361, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98354, 19.98348, 19.98364, 19.98358, 19.98402, 
    19.98402, 19.984, 19.98406, 19.98406, 19.98411, 19.98407, 19.98405, 
    19.984, 19.98397, 19.98395, 19.98389, 19.98382, 19.98373, 19.98367, 
    19.98363, 19.98365, 19.98363, 19.98365, 19.98367, 19.98353, 19.98361, 
    19.98349, 19.9835, 19.98355, 19.9835, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98396, 19.98394, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98362, 19.98362, 
    19.9836, 19.98364, 19.98359, 19.98359, 19.98361, 19.9835, 19.98353, 
    19.9835, 19.98352, 19.98402, 19.984, 19.98401, 19.98399, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98384, 19.98376, 19.98383, 19.98382, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.9837, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98346, 19.98347, 19.98342, 
    19.98396, 19.98393, 19.98393, 19.9839, 19.98387, 19.98382, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98373, 19.98391, 19.98388, 
    19.98389, 19.98396, 19.98376, 19.98386, 19.98367, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98335, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.9837, 19.98363, 19.98387, 19.98375, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98377, 19.98375, 19.98366, 19.9837, 19.98343, 
    19.98355, 19.98322, 19.98331, 19.98394, 19.98391, 19.98381, 19.98386, 
    19.98372, 19.98368, 19.98365, 19.98362, 19.98361, 19.98359, 19.98363, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98382, 
    19.98376, 19.9837, 19.98369, 19.98368, 19.98362, 19.98372, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98384, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98357, 19.9836, 19.9836, 19.98365, 19.98367, 
    19.98374, 19.98379, 19.98383, 19.98382, 19.98378, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98373, 19.98366, 19.98369, 19.98362, 19.98376, 
    19.98364, 19.9838, 19.98378, 19.98374, 19.98366, 19.98364, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98379, 19.98381, 
    19.98379, 19.98376, 19.98369, 19.98363, 19.98355, 19.98354, 19.98346, 
    19.98352, 19.98341, 19.98351, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98357, 19.98362, 19.98356, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.9838, 19.98376, 19.98377, 19.98369, 
    19.98373, 19.9836, 19.98356, 19.98343, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.98571, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98558, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98529, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98564, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98522, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98565, 19.98562, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98527, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98567, 19.98567, 19.98571, 19.98567, 19.98566, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98522, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98572, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98528, 
    19.98526, 19.98529, 19.98526, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98563, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98535, 19.98526, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98556, 19.98553, 19.9855, 19.98545, 19.98538, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98554, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.9853, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98548, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98522, 19.98492, 19.985, 19.98556, 19.98554, 19.98545, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98528, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98535, 19.98534, 19.98533, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98534, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98542, 19.98534, 19.98527, 
    19.98529, 19.98524, 19.98537, 19.98532, 19.98534, 19.98528, 19.98541, 
    19.9853, 19.98543, 19.98542, 19.98539, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98539, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98518, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98493, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222428, 0.7222433, 0.7222413, 0.7222424, 0.722241, 0.7222448, 
    0.7222427, 0.722244, 0.7222451, 0.7222373, 0.7222412, 0.7222333, 
    0.7222357, 0.7222296, 0.7222337, 0.7222288, 0.7222297, 0.7222269, 
    0.7222277, 0.7222241, 0.7222265, 0.7222221, 0.7222246, 0.7222242, 
    0.7222266, 0.7222404, 0.7222378, 0.7222406, 0.7222401, 0.7222403, 
    0.7222424, 0.7222434, 0.7222455, 0.7222452, 0.7222435, 0.72224, 
    0.7222412, 0.7222382, 0.7222382, 0.7222348, 0.7222364, 0.7222307, 
    0.7222323, 0.7222276, 0.7222288, 0.7222277, 0.7222281, 0.7222277, 
    0.7222294, 0.7222286, 0.7222302, 0.7222361, 0.7222344, 0.7222396, 
    0.7222427, 0.7222447, 0.7222462, 0.722246, 0.7222456, 0.7222435, 
    0.7222416, 0.7222402, 0.7222392, 0.7222382, 0.7222353, 0.7222338, 
    0.7222304, 0.722231, 0.72223, 0.7222289, 0.7222272, 0.7222275, 0.7222268, 
    0.72223, 0.7222279, 0.7222313, 0.7222304, 0.722238, 0.7222409, 0.7222421, 
    0.7222432, 0.7222458, 0.722244, 0.7222447, 0.722243, 0.7222419, 
    0.7222425, 0.7222392, 0.7222404, 0.7222337, 0.7222366, 0.7222291, 
    0.7222309, 0.7222286, 0.7222298, 0.7222278, 0.7222295, 0.7222265, 
    0.7222258, 0.7222263, 0.7222245, 0.7222297, 0.7222277, 0.7222425, 
    0.7222424, 0.722242, 0.7222438, 0.7222439, 0.7222455, 0.7222441, 
    0.7222435, 0.7222419, 0.722241, 0.7222401, 0.7222381, 0.722236, 
    0.7222329, 0.7222307, 0.7222293, 0.7222302, 0.7222294, 0.7222303, 
    0.7222307, 0.7222261, 0.7222286, 0.7222248, 0.722225, 0.7222267, 
    0.722225, 0.7222424, 0.7222428, 0.7222446, 0.7222432, 0.7222457, 
    0.7222443, 0.7222435, 0.7222404, 0.7222398, 0.7222391, 0.7222379, 
    0.7222363, 0.7222335, 0.7222311, 0.7222289, 0.722229, 0.722229, 
    0.7222285, 0.7222297, 0.7222283, 0.7222281, 0.7222286, 0.722225, 
    0.7222261, 0.722225, 0.7222257, 0.7222427, 0.7222418, 0.7222423, 
    0.7222415, 0.7222421, 0.7222394, 0.7222385, 0.7222348, 0.7222363, 
    0.7222339, 0.7222361, 0.7222357, 0.7222338, 0.722236, 0.7222312, 
    0.7222344, 0.7222285, 0.7222317, 0.7222283, 0.7222289, 0.7222279, 
    0.7222269, 0.7222258, 0.7222236, 0.7222241, 0.7222223, 0.7222406, 
    0.7222395, 0.7222396, 0.7222384, 0.7222376, 0.7222357, 0.7222328, 
    0.722234, 0.7222319, 0.7222315, 0.7222345, 0.7222327, 0.7222388, 
    0.7222378, 0.7222384, 0.7222405, 0.7222337, 0.7222372, 0.7222307, 
    0.7222326, 0.722227, 0.7222298, 0.7222244, 0.7222221, 0.7222199, 
    0.7222174, 0.7222389, 0.7222396, 0.7222383, 0.7222365, 0.7222348, 
    0.7222325, 0.7222323, 0.7222318, 0.7222307, 0.7222298, 0.7222317, 
    0.7222296, 0.7222375, 0.7222334, 0.7222399, 0.7222379, 0.7222366, 
    0.7222372, 0.7222341, 0.7222333, 0.7222303, 0.7222319, 0.7222227, 
    0.7222267, 0.7222155, 0.7222186, 0.7222399, 0.7222389, 0.7222354, 
    0.7222371, 0.7222323, 0.7222311, 0.7222302, 0.722229, 0.7222289, 
    0.7222282, 0.7222294, 0.7222282, 0.7222325, 0.7222306, 0.7222358, 
    0.7222345, 0.7222351, 0.7222358, 0.7222338, 0.7222317, 0.7222316, 
    0.722231, 0.722229, 0.7222323, 0.7222221, 0.7222284, 0.7222378, 
    0.7222359, 0.7222356, 0.7222363, 0.7222313, 0.7222331, 0.7222282, 
    0.7222295, 0.7222273, 0.7222284, 0.7222286, 0.72223, 0.7222309, 
    0.7222331, 0.7222348, 0.7222362, 0.7222359, 0.7222344, 0.7222315, 
    0.7222289, 0.7222295, 0.7222275, 0.7222327, 0.7222305, 0.7222313, 
    0.7222292, 0.722234, 0.7222298, 0.722235, 0.7222345, 0.7222332, 
    0.7222304, 0.7222297, 0.7222291, 0.7222295, 0.7222314, 0.7222318, 
    0.7222332, 0.7222336, 0.7222347, 0.7222356, 0.7222347, 0.7222339, 
    0.7222314, 0.7222293, 0.7222269, 0.7222263, 0.7222236, 0.7222258, 
    0.7222221, 0.7222252, 0.7222198, 0.7222297, 0.7222254, 0.7222331, 
    0.7222323, 0.7222307, 0.7222273, 0.7222292, 0.722227, 0.7222318, 
    0.7222343, 0.722235, 0.7222362, 0.7222349, 0.722235, 0.7222338, 
    0.7222342, 0.7222314, 0.7222329, 0.7222286, 0.722227, 0.7222226, 
    0.7222198, 0.722217, 0.7222158, 0.7222154, 0.7222153 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  2.055969e-20, 0, 5.139921e-21, -2.569961e-20, 3.083953e-20, -2.569961e-20, 
    3.083953e-20, -5.139921e-21, 2.055969e-20, -5.139921e-21, -1.027984e-20, 
    2.569961e-20, -2.569961e-20, 2.006177e-36, -2.006177e-36, -2.569961e-20, 
    -1.027984e-20, -2.055969e-20, -3.083953e-20, -1.541976e-20, 
    -1.541976e-20, 1.027984e-20, 3.083953e-20, 2.055969e-20, -1.541976e-20, 
    3.083953e-20, 2.055969e-20, -2.055969e-20, 1.027984e-20, -1.027984e-20, 
    2.006177e-36, -2.055969e-20, 2.006177e-36, 2.569961e-20, 5.139921e-21, 
    -5.139921e-21, -2.569961e-20, 2.055969e-20, 0, -2.569961e-20, 
    2.055969e-20, -1.027984e-20, -5.139921e-21, -4.111937e-20, 1.541976e-20, 
    -1.027984e-20, 3.083953e-20, -1.027984e-20, -5.139921e-21, 0, 
    -2.006177e-36, -2.569961e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    2.055969e-20, 1.541976e-20, 3.597945e-20, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, -2.006177e-36, -4.625929e-20, -1.027984e-20, 1.027984e-20, 
    -2.055969e-20, 2.006177e-36, -2.569961e-20, 2.569961e-20, 3.083953e-20, 
    -2.569961e-20, -2.569961e-20, -1.541976e-20, 0, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.541976e-20, 1.027984e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, -5.139921e-21, 
    2.055969e-20, 0, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    5.653913e-20, -1.541976e-20, -1.027984e-20, -2.006177e-36, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, -1.541976e-20, -1.027984e-20, 
    1.027984e-20, 2.569961e-20, 2.055969e-20, -3.597945e-20, -5.139921e-20, 
    1.027984e-20, 2.055969e-20, -2.569961e-20, 2.055969e-20, 2.006177e-36, 
    -2.055969e-20, 2.569961e-20, 3.083953e-20, -5.139921e-21, 2.006177e-36, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 0, 
    -1.027984e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, -2.055969e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, 1.027984e-20, -3.083953e-20, 
    -5.653913e-20, 0, 5.139921e-21, 2.569961e-20, 3.083953e-20, 0, 
    -2.569961e-20, 3.083953e-20, 2.569961e-20, -5.139921e-21, 2.006177e-36, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 2.006177e-36, 
    -5.139921e-21, -1.027984e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    0, 2.569961e-20, 2.006177e-36, 3.597945e-20, 0, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    1.541976e-20, 2.006177e-36, -5.139921e-21, -3.597945e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-20, -2.569961e-20, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, -4.111937e-20, -3.083953e-20, -1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 3.083953e-20, 3.083953e-20, -5.139921e-21, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, -1.541976e-20, 2.569961e-20, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, -2.569961e-20, -5.139921e-21, 1.541976e-20, 
    -1.027984e-20, -5.139921e-21, 0, -1.027984e-20, 2.006177e-36, 0, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -3.083953e-20, -1.541976e-20, 0, 3.083953e-20, 5.139921e-21, 
    2.055969e-20, 1.027984e-20, 2.569961e-20, 2.055969e-20, 5.139921e-21, 
    2.055969e-20, 1.027984e-20, 3.597945e-20, -1.541976e-20, 2.055969e-20, 
    -5.653913e-20, 1.541976e-20, -5.139921e-21, -2.569961e-20, 1.027984e-20, 
    2.006177e-36, -5.139921e-21, 3.083953e-20, -3.597945e-20, -1.541976e-20, 
    -1.027984e-20, -2.569961e-20, 3.083953e-20, -2.569961e-20, -2.055969e-20, 
    -4.111937e-20, 2.055969e-20, -3.083953e-20, 2.006177e-36, 2.055969e-20, 
    2.569961e-20, -1.541976e-20, 2.569961e-20, 1.027984e-20, 2.055969e-20, 
    -3.083953e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, -2.055969e-20, 0, -2.569961e-20, 6.681898e-20, 
    -5.139921e-21, 4.111937e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, -2.569961e-20, 2.055969e-20, 
    1.541976e-20, -4.111937e-20, -2.055969e-20, 1.541976e-20, 0, 
    1.027984e-20, 4.111937e-20, 1.541976e-20, 2.006177e-36, -1.027984e-20, 
    -2.569961e-20, 1.027984e-20, -2.055969e-20, -2.055969e-20, -2.055969e-20, 
    -2.569961e-20, 4.625929e-20, -2.569961e-20, 1.541976e-20, -2.569961e-20, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, -2.006177e-36, 5.139921e-20, -5.139921e-21, 
    0, 1.541976e-20, 2.006177e-36, 4.111937e-20, -2.006177e-36, 
    -5.139921e-21, 5.139921e-21, -2.055969e-20, -5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-20, 
    -1.027984e-20, -2.006177e-36, 1.027984e-20, 2.006177e-36, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 1.541976e-20, 1.541976e-20, 0, 
    -5.139921e-21, -2.006177e-36, 2.055969e-20, -3.597945e-20,
  1.027984e-20, -5.139921e-21, -3.083953e-20, -1.027984e-20, 0, 
    -1.027984e-20, -2.569961e-20, -1.027984e-20, 2.569961e-20, -5.139921e-21, 
    -3.083953e-20, -5.139921e-21, 1.541976e-20, 2.055969e-20, 5.139921e-21, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 0, 5.139921e-21, 
    1.027984e-20, 0, -5.139921e-21, 2.569961e-20, 2.055969e-20, 
    -5.139921e-21, 2.006177e-36, -2.006177e-36, -2.055969e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -2.569961e-20, 1.027984e-20, -3.597945e-20, 
    4.625929e-20, 2.055969e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    2.569961e-20, 2.055969e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, 
    -5.139921e-21, -2.006177e-36, -5.139921e-21, 2.569961e-20, -1.027984e-20, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 0, 
    1.541976e-20, 5.139921e-21, 3.083953e-20, 1.541976e-20, 0, -2.006177e-36, 
    2.055969e-20, 2.055969e-20, -1.027984e-20, -2.006177e-36, 0, 
    1.027984e-20, 0, -1.027984e-20, -1.541976e-20, 5.139921e-21, 
    -2.569961e-20, -2.569961e-20, -3.083953e-20, 0, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 0, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 2.055969e-20, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, -2.569961e-20, -2.569961e-20, -3.597945e-20, 
    1.027984e-20, 0, -1.027984e-20, 5.139921e-21, 0, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -2.055969e-20, 1.541976e-20, 1.541976e-20, 
    -1.027984e-20, -5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 0, 5.139921e-21, -1.027984e-20, 
    -2.006177e-36, 1.541976e-20, -2.569961e-20, 5.139921e-21, 3.083953e-20, 
    5.139921e-21, 0, 2.569961e-20, 1.027984e-20, 2.055969e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -1.541976e-20, 5.139921e-21, 1.027984e-20, 0, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 0, 1.027984e-20, -2.006177e-36, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -3.083953e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, 5.139921e-21, 5.139921e-21, 2.569961e-20, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -3.083953e-20, 2.055969e-20, 2.055969e-20, 5.139921e-21, 
    -5.139921e-21, 0, 0, -3.597945e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 3.083953e-20, 5.139921e-21, 0, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, -5.139921e-21, 0, 
    -1.027984e-20, 2.055969e-20, -3.597945e-20, 1.541976e-20, -1.541976e-20, 
    -1.027984e-20, 2.569961e-20, 0, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, -2.055969e-20, -3.597945e-20, -2.006177e-36, 
    -2.569961e-20, 1.027984e-20, 3.083953e-20, -2.055969e-20, -5.139921e-21, 
    0, -1.027984e-20, -1.541976e-20, -2.055969e-20, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, 2.569961e-20, -3.597945e-20, 
    3.597945e-20, 1.027984e-20, 2.569961e-20, -2.055969e-20, -3.083953e-20, 
    1.027984e-20, 5.139921e-21, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -2.055969e-20, 2.006177e-36, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, -5.139921e-21, 
    2.569961e-20, -3.597945e-20, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    2.055969e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, -2.006177e-36, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 2.055969e-20, 
    2.055969e-20, -1.027984e-20, 3.083953e-20, -3.083953e-20, 0, 
    3.083953e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -3.597945e-20, -3.597945e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, 0, 5.139921e-21, 1.027984e-20, -5.139921e-21, 2.569961e-20, 
    -1.541976e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, 3.083953e-20, 
    -1.027984e-20, 1.541976e-20, 0, 1.027984e-20, -2.569961e-20, 
    1.027984e-20, -5.139921e-21, 2.006177e-36, 2.055969e-20, 5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 1.541976e-20, 4.111937e-20, 5.139921e-21, 
    -2.569961e-20, 2.569961e-20, 0, 1.027984e-20, -2.569961e-20, 
    2.055969e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, 1.027984e-20, 
    -3.083953e-20, 1.541976e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    2.569961e-20, -2.055969e-20,
  5.139921e-21, -2.055969e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 
    -1.541976e-20, 0, 2.006177e-36, 3.083953e-20, -3.083953e-20, 0, 
    3.597945e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, -2.569961e-20, 2.569961e-20, -1.027984e-20, -2.055969e-20, 
    0, -5.139921e-21, 1.541976e-20, 5.139921e-21, -2.006177e-36, 
    1.027984e-20, 2.055969e-20, 5.139921e-21, -2.006177e-36, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, 2.055969e-20, 2.055969e-20, 2.569961e-20, 
    5.139921e-21, 2.006177e-36, -2.006177e-36, 2.055969e-20, -1.541976e-20, 
    2.569961e-20, -1.027984e-20, 2.055969e-20, 0, 2.055969e-20, 
    -5.139921e-21, -2.569961e-20, 1.541976e-20, 5.139921e-21, 0, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -2.569961e-20, 
    -1.027984e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    0, 2.006177e-36, -2.569961e-20, 1.541976e-20, -2.006177e-36, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, -3.083953e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.569961e-20, -3.597945e-20, 5.139921e-21, 0, -2.006177e-36, 
    5.139921e-21, 2.055969e-20, -3.083953e-20, -2.055969e-20, -2.006177e-36, 
    0, 0, 1.541976e-20, 1.027984e-20, 0, 2.006177e-36, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -5.139921e-21, -1.027984e-20, 0, -1.541976e-20, 2.569961e-20, 
    1.027984e-20, -1.027984e-20, 2.055969e-20, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, 0, 
    3.083953e-20, -2.055969e-20, 0, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -3.597945e-20, 0, 2.055969e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-20, 
    2.055969e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 0, 
    -2.055969e-20, 1.027984e-20, 2.055969e-20, -1.027984e-20, -2.569961e-20, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, 2.569961e-20, 5.139921e-21, 
    -2.006177e-36, 0, -2.055969e-20, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 1.027984e-20, 1.027984e-20, 
    2.006177e-36, 0, -5.139921e-21, 0, -1.541976e-20, -2.055969e-20, 
    1.541976e-20, -1.027984e-20, 0, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, 
    5.139921e-21, 0, 2.055969e-20, 1.541976e-20, 1.027984e-20, -2.055969e-20, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, -3.083953e-20, 2.055969e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    0, 1.027984e-20, -2.055969e-20, -2.006177e-36, -1.027984e-20, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, -2.006177e-36, -2.006177e-36, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, -2.055969e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -4.625929e-20, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-20, -1.541976e-20, 
    0, -2.006177e-36, 3.083953e-20, 1.541976e-20, -1.541976e-20, 
    -3.083953e-20, -2.055969e-20, 2.006177e-36, 2.055969e-20, -1.027984e-20, 
    2.055969e-20, 2.006177e-36, 1.027984e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    2.569961e-20, -2.006177e-36, -1.027984e-20, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, -2.569961e-20, 5.139921e-21, 1.541976e-20, 2.569961e-20, 
    -2.006177e-36, 1.541976e-20, -2.569961e-20, -2.055969e-20, 5.139921e-21, 
    1.541976e-20, 2.055969e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, -5.139921e-20, -5.139921e-21, -1.027984e-20, 2.055969e-20, 
    -1.027984e-20, -2.055969e-20, 1.541976e-20, 2.006177e-36, -2.055969e-20, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    0, 1.541976e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, -1.541976e-20, 0, -2.569961e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, 2.569961e-20, -2.055969e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -2.569961e-20, 1.541976e-20, 
    -5.139921e-21, 0, -1.027984e-20, 1.541976e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, -3.083953e-20, 1.027984e-20, 
    3.597945e-20, 5.139921e-21, -1.541976e-20, 2.055969e-20, -3.597945e-20, 
    -2.055969e-20, -1.027984e-20, 2.055969e-20, 2.006177e-36, 2.055969e-20, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, -3.597945e-20, 
    0, -2.055969e-20, -4.111937e-20, -2.569961e-20, -2.006177e-36, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, 3.083953e-20, 2.055969e-20, 
    -2.569961e-20, -5.139921e-21,
  2.569961e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 0, -2.569961e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 1.541976e-20, -1.027984e-20, 
    1.541976e-20, 2.055969e-20, 0, 2.055969e-20, -5.139921e-21, 
    -1.027984e-20, 0, -4.111937e-20, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 0, -2.006177e-36, 1.027984e-20, -1.541976e-20, 
    -2.006177e-36, -1.541976e-20, -2.055969e-20, -1.027984e-20, 0, 
    -1.541976e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, -3.083953e-20, 
    3.083953e-20, -2.055969e-20, -1.541976e-20, -4.111937e-20, -5.139921e-21, 
    1.541976e-20, 0, 2.055969e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    -2.569961e-20, -2.006177e-36, 1.541976e-20, 4.111937e-20, -3.597945e-20, 
    -5.139921e-21, -3.083953e-20, 5.139921e-21, -3.597945e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, 4.111937e-20, 
    2.569961e-20, -2.569961e-20, -5.139921e-21, 1.027984e-20, -3.083953e-20, 
    2.055969e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    1.541976e-20, -3.083953e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, 
    0, 1.027984e-20, 1.541976e-20, 5.139921e-21, 2.569961e-20, -1.541976e-20, 
    -2.055969e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, 
    2.006177e-36, 0, 2.569961e-20, 1.027984e-20, 5.139921e-20, -2.006177e-36, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, 5.139921e-21, 0, 1.027984e-20, 
    3.597945e-20, 1.541976e-20, 3.597945e-20, 5.139921e-21, -1.541976e-20, 
    1.541976e-20, -3.083953e-20, 1.027984e-20, 0, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 5.139921e-21, -3.083953e-20, -1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -3.597945e-20, 0, 1.027984e-20, 
    -3.597945e-20, -1.027984e-20, -5.139921e-21, 4.111937e-20, 3.597945e-20, 
    2.055969e-20, -5.139921e-21, 2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 1.027984e-20, -1.027984e-20, 0, 
    -5.139921e-21, -2.055969e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    3.083953e-20, -5.139921e-21, -2.055969e-20, -1.541976e-20, -3.597945e-20, 
    -2.006177e-36, -5.139921e-21, 4.625929e-20, 0, -3.597945e-20, 0, 
    -5.139921e-21, 1.541976e-20, -3.597945e-20, 0, -3.083953e-20, 
    4.625929e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -2.569961e-20, 3.597945e-20, -3.083953e-20, 5.139921e-21, 5.139921e-21, 
    3.597945e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, -4.111937e-20, 
    0, -1.541976e-20, 2.006177e-36, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, 0, 5.139921e-21, 0, 
    -2.569961e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 0, 
    3.083953e-20, 2.006177e-36, -2.006177e-36, 1.541976e-20, -2.569961e-20, 
    2.006177e-36, -5.139921e-21, -2.055969e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -3.083953e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.541976e-20, -1.541976e-20, -5.139921e-21, 0, 5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    2.569961e-20, -2.055969e-20, 2.569961e-20, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -2.569961e-20, 2.055969e-20, 5.139921e-21, 2.569961e-20, 
    -2.569961e-20, -2.006177e-36, 1.541976e-20, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, -5.139921e-21, 3.597945e-20, 3.083953e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.055969e-20, 2.055969e-20, 
    5.139921e-21, -2.569961e-20, 5.139921e-21, 0, 3.083953e-20, 1.027984e-20, 
    -3.083953e-20, 3.083953e-20, 2.055969e-20, -2.569961e-20, 3.597945e-20, 
    -1.027984e-20, -2.055969e-20, 1.027984e-20, -4.111937e-20, 1.027984e-20, 
    2.006177e-36, -5.139921e-21, 5.139921e-21, 0, 5.139921e-21, 
    -3.597945e-20, -5.139921e-21, 4.625929e-20, -2.055969e-20, 5.653913e-20, 
    -3.597945e-20, -3.083953e-20, 2.055969e-20, 0, 1.027984e-20, 
    3.083953e-20, 1.541976e-20, -5.139921e-21, 0, 1.027984e-20, 
    -2.569961e-20, -4.111937e-20, 4.625929e-20, 0, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 3.597945e-20, 5.139921e-21, 5.139921e-21, 
    3.083953e-20, 5.139921e-21, -1.027984e-20, 4.111937e-20, 1.027984e-20, 0, 
    1.027984e-20, -5.139921e-21, 2.006177e-36, 2.569961e-20, -2.055969e-20, 
    2.569961e-20, 5.139921e-21, 5.139921e-20, -1.027984e-20, 5.139921e-21, 
    2.006177e-36, -5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -3.597945e-20, -2.055969e-20, 
    -3.083953e-20, -1.027984e-20, -2.055969e-20, -1.027984e-20, 2.055969e-20, 
    2.006177e-36, 1.541976e-20, -1.541976e-20, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, -4.111937e-20, 0, -2.006177e-36, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, 3.083953e-20, -1.541976e-20,
  5.139921e-21, 5.139921e-21, 0, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -4.625929e-20, -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -2.055969e-20, 5.139921e-21, 0, 
    1.541976e-20, -2.006177e-36, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 1.027984e-20, 5.139921e-21, 2.055969e-20, 1.027984e-20, 
    2.055969e-20, 5.139921e-21, 3.083953e-20, -2.055969e-20, 5.139921e-21, 
    1.027984e-20, 3.597945e-20, 5.139921e-21, -2.006177e-36, -1.027984e-20, 
    1.541976e-20, -2.006177e-36, -1.027984e-20, 0, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, 2.055969e-20, 5.139921e-21, -1.027984e-20, 
    2.006177e-36, -2.006177e-36, 0, 5.139921e-21, 1.027984e-20, 3.083953e-20, 
    5.139921e-21, 0, -1.027984e-20, 3.083953e-20, 2.569961e-20, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 3.083953e-20, 4.625929e-20, 2.006177e-36, -5.139921e-21, 
    -2.055969e-20, 1.541976e-20, -3.083953e-20, 0, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, -2.569961e-20, -2.569961e-20, 1.027984e-20, 
    1.541976e-20, 1.027984e-20, 2.006177e-36, -1.541976e-20, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, -1.027984e-20, 0, -1.027984e-20, 
    -5.139921e-21, 0, 1.541976e-20, -3.083953e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, -1.541976e-20, 4.625929e-20, 3.083953e-20, 4.111937e-20, 
    -5.139921e-21, -2.055969e-20, -5.139921e-21, 5.139921e-21, 3.083953e-20, 
    2.006177e-36, 5.139921e-21, 2.006177e-36, 0, -3.083953e-20, 5.139921e-21, 
    2.055969e-20, -2.006177e-36, -2.569961e-20, 1.541976e-20, 4.111937e-20, 
    -1.027984e-20, 2.569961e-20, 2.006177e-36, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 1.027984e-20, -2.055969e-20, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -2.569961e-20, -1.541976e-20, 0, 
    1.541976e-20, -5.139921e-21, -2.006177e-36, -5.139921e-21, -1.541976e-20, 
    4.111937e-20, 0, 1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -2.055969e-20, -2.569961e-20, 1.027984e-20, 1.027984e-20, -4.625929e-20, 
    3.083953e-20, -2.569961e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 0, -2.055969e-20, -2.055969e-20, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, -4.625929e-20, 1.027984e-20, 
    -1.027984e-20, 3.083953e-20, 1.027984e-20, -3.083953e-20, -2.055969e-20, 
    -5.139921e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 0, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -1.541976e-20, 3.083953e-20, -2.055969e-20, 
    -5.139921e-21, 0, -1.541976e-20, 1.541976e-20, 1.541976e-20, 
    -1.027984e-20, -2.006177e-36, 2.569961e-20, -5.139921e-21, 1.541976e-20, 
    2.569961e-20, -3.083953e-20, -4.625929e-20, -1.027984e-20, -2.006177e-36, 
    -2.055969e-20, 1.027984e-20, 1.541976e-20, 0, -5.139921e-21, 
    -2.006177e-36, -2.055969e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, -2.569961e-20, 
    5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    2.055969e-20, 1.541976e-20, -2.006177e-36, 3.597945e-20, -2.055969e-20, 
    1.027984e-20, 5.139921e-21, -2.055969e-20, 0, -2.055969e-20, 
    2.569961e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 1.541976e-20, 
    3.083953e-20, 1.027984e-20, 0, 3.597945e-20, -2.055969e-20, 1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, 5.139921e-21, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 3.597945e-20, 1.027984e-20, 
    2.006177e-36, -1.541976e-20, 0, -1.027984e-20, -2.006177e-36, 
    -2.006177e-36, 0, 4.111937e-20, -1.027984e-20, -1.027984e-20, 0, 
    -2.006177e-36, -5.139921e-21, 2.569961e-20, 5.139921e-21, 1.541976e-20, 
    3.083953e-20, -5.139921e-21, 2.055969e-20, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 0, 3.597945e-20, -5.139921e-21, 2.006177e-36, 
    1.541976e-20, 1.541976e-20, -2.055969e-20, 1.027984e-20, -1.027984e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 3.083953e-20, -1.541976e-20, 
    -5.139921e-21, -2.006177e-36, -1.027984e-20, -1.027984e-20, 
    -2.569961e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.006177e-36, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 2.055969e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 2.055969e-20, -5.139921e-21, 2.055969e-20, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, -2.006177e-36, 5.139921e-21, 
    3.083953e-20, 0, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, 
    1.541976e-20, -2.569961e-20, 0, -2.055969e-20,
  8.598664e-29, 8.598635e-29, 8.598641e-29, 8.598618e-29, 8.59863e-29, 
    8.598615e-29, 8.598658e-29, 8.598634e-29, 8.598649e-29, 8.598662e-29, 
    8.598573e-29, 8.598617e-29, 8.598527e-29, 8.598556e-29, 8.598485e-29, 
    8.598532e-29, 8.598476e-29, 8.598486e-29, 8.598454e-29, 8.598463e-29, 
    8.598422e-29, 8.59845e-29, 8.5984e-29, 8.598429e-29, 8.598424e-29, 
    8.598451e-29, 8.598608e-29, 8.598578e-29, 8.59861e-29, 8.598606e-29, 
    8.598607e-29, 8.59863e-29, 8.598642e-29, 8.598666e-29, 8.598662e-29, 
    8.598644e-29, 8.598604e-29, 8.598617e-29, 8.598583e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598498e-29, 8.598516e-29, 8.598463e-29, 
    8.598476e-29, 8.598463e-29, 8.598468e-29, 8.598463e-29, 8.598483e-29, 
    8.598475e-29, 8.598492e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598674e-29, 8.598671e-29, 8.598667e-29, 
    8.598643e-29, 8.598622e-29, 8.598606e-29, 8.598595e-29, 8.598584e-29, 
    8.598551e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598478e-29, 8.598459e-29, 8.598462e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598505e-29, 8.598494e-29, 8.598581e-29, 8.598613e-29, 
    8.598627e-29, 8.59864e-29, 8.598669e-29, 8.598649e-29, 8.598657e-29, 
    8.598638e-29, 8.598625e-29, 8.598631e-29, 8.598594e-29, 8.598609e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.5985e-29, 8.598474e-29, 
    8.598487e-29, 8.598465e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598448e-29, 8.598427e-29, 8.598486e-29, 8.598463e-29, 8.598632e-29, 
    8.598631e-29, 8.598626e-29, 8.598646e-29, 8.598648e-29, 8.598666e-29, 
    8.598649e-29, 8.598643e-29, 8.598625e-29, 8.598614e-29, 8.598604e-29, 
    8.598582e-29, 8.598557e-29, 8.598523e-29, 8.598498e-29, 8.598482e-29, 
    8.598492e-29, 8.598483e-29, 8.598493e-29, 8.598498e-29, 8.598445e-29, 
    8.598475e-29, 8.59843e-29, 8.598433e-29, 8.598453e-29, 8.598433e-29, 
    8.59863e-29, 8.598636e-29, 8.598655e-29, 8.59864e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598609e-29, 8.598601e-29, 8.598593e-29, 
    8.59858e-29, 8.598562e-29, 8.59853e-29, 8.598502e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598473e-29, 8.598486e-29, 8.59847e-29, 
    8.598468e-29, 8.598475e-29, 8.598433e-29, 8.598445e-29, 8.598433e-29, 
    8.598441e-29, 8.598634e-29, 8.598624e-29, 8.59863e-29, 8.59862e-29, 
    8.598627e-29, 8.598596e-29, 8.598587e-29, 8.598544e-29, 8.598562e-29, 
    8.598534e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598504e-29, 8.598541e-29, 8.598473e-29, 8.598509e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598455e-29, 8.598442e-29, 8.598418e-29, 
    8.598423e-29, 8.598403e-29, 8.59861e-29, 8.598598e-29, 8.598599e-29, 
    8.598586e-29, 8.598576e-29, 8.598556e-29, 8.598522e-29, 8.598535e-29, 
    8.598512e-29, 8.598507e-29, 8.598542e-29, 8.59852e-29, 8.598589e-29, 
    8.598578e-29, 8.598585e-29, 8.598609e-29, 8.598532e-29, 8.598571e-29, 
    8.598498e-29, 8.598519e-29, 8.598456e-29, 8.598488e-29, 8.598426e-29, 
    8.5984e-29, 8.598375e-29, 8.598346e-29, 8.598591e-29, 8.5986e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598488e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598528e-29, 8.598603e-29, 8.59858e-29, 8.598565e-29, 
    8.598571e-29, 8.598536e-29, 8.598527e-29, 8.598494e-29, 8.598511e-29, 
    8.598406e-29, 8.598453e-29, 8.598324e-29, 8.59836e-29, 8.598603e-29, 
    8.598591e-29, 8.598551e-29, 8.59857e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598479e-29, 8.598477e-29, 8.598469e-29, 8.598482e-29, 
    8.59847e-29, 8.598518e-29, 8.598497e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598556e-29, 8.598533e-29, 8.598509e-29, 8.598508e-29, 
    8.598501e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598472e-29, 
    8.598578e-29, 8.598557e-29, 8.598554e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598469e-29, 8.598485e-29, 8.598459e-29, 8.598472e-29, 
    8.598474e-29, 8.598489e-29, 8.5985e-29, 8.598524e-29, 8.598545e-29, 
    8.598561e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598477e-29, 
    8.598483e-29, 8.598461e-29, 8.59852e-29, 8.598495e-29, 8.598505e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598547e-29, 8.598542e-29, 
    8.598525e-29, 8.598494e-29, 8.598487e-29, 8.598479e-29, 8.598484e-29, 
    8.598506e-29, 8.59851e-29, 8.598526e-29, 8.59853e-29, 8.598543e-29, 
    8.598553e-29, 8.598544e-29, 8.598534e-29, 8.598506e-29, 8.598482e-29, 
    8.598455e-29, 8.598448e-29, 8.598417e-29, 8.598442e-29, 8.5984e-29, 
    8.598436e-29, 8.598374e-29, 8.598486e-29, 8.598437e-29, 8.598525e-29, 
    8.598516e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598456e-29, 
    8.59851e-29, 8.598539e-29, 8.598546e-29, 8.59856e-29, 8.598546e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598506e-29, 8.598523e-29, 
    8.598474e-29, 8.598456e-29, 8.598405e-29, 8.598374e-29, 8.598342e-29, 
    8.598328e-29, 8.598324e-29, 8.598322e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.164843e-08, 1.169965e-08, 1.168969e-08, 1.1731e-08, 1.170809e-08, 
    1.173514e-08, 1.165882e-08, 1.170168e-08, 1.167432e-08, 1.165304e-08, 
    1.181117e-08, 1.173285e-08, 1.189252e-08, 1.184257e-08, 1.196805e-08, 
    1.188475e-08, 1.198484e-08, 1.196564e-08, 1.202342e-08, 1.200687e-08, 
    1.208078e-08, 1.203106e-08, 1.211909e-08, 1.206891e-08, 1.207676e-08, 
    1.202942e-08, 1.174861e-08, 1.180142e-08, 1.174548e-08, 1.175301e-08, 
    1.174963e-08, 1.170856e-08, 1.168787e-08, 1.164452e-08, 1.165239e-08, 
    1.168423e-08, 1.17564e-08, 1.17319e-08, 1.179364e-08, 1.179224e-08, 
    1.186098e-08, 1.182999e-08, 1.194551e-08, 1.191268e-08, 1.200756e-08, 
    1.19837e-08, 1.200644e-08, 1.199954e-08, 1.200653e-08, 1.197153e-08, 
    1.198653e-08, 1.195573e-08, 1.183579e-08, 1.187104e-08, 1.176591e-08, 
    1.170269e-08, 1.16607e-08, 1.16309e-08, 1.163511e-08, 1.164314e-08, 
    1.168441e-08, 1.172321e-08, 1.175278e-08, 1.177256e-08, 1.179204e-08, 
    1.185103e-08, 1.188225e-08, 1.195215e-08, 1.193954e-08, 1.196091e-08, 
    1.198133e-08, 1.20156e-08, 1.200996e-08, 1.202506e-08, 1.196035e-08, 
    1.200336e-08, 1.193235e-08, 1.195177e-08, 1.179735e-08, 1.173851e-08, 
    1.17135e-08, 1.169161e-08, 1.163835e-08, 1.167513e-08, 1.166063e-08, 
    1.169512e-08, 1.171704e-08, 1.17062e-08, 1.17731e-08, 1.174709e-08, 
    1.18841e-08, 1.182509e-08, 1.197894e-08, 1.194213e-08, 1.198777e-08, 
    1.196448e-08, 1.200439e-08, 1.196847e-08, 1.203068e-08, 1.204423e-08, 
    1.203497e-08, 1.207053e-08, 1.196648e-08, 1.200644e-08, 1.17059e-08, 
    1.170766e-08, 1.17159e-08, 1.16797e-08, 1.167748e-08, 1.16443e-08, 
    1.167382e-08, 1.16864e-08, 1.171831e-08, 1.173719e-08, 1.175513e-08, 
    1.179458e-08, 1.183864e-08, 1.190025e-08, 1.194451e-08, 1.197418e-08, 
    1.195599e-08, 1.197205e-08, 1.19541e-08, 1.194568e-08, 1.203916e-08, 
    1.198667e-08, 1.206542e-08, 1.206106e-08, 1.202542e-08, 1.206155e-08, 
    1.17089e-08, 1.169873e-08, 1.166341e-08, 1.169105e-08, 1.164069e-08, 
    1.166888e-08, 1.168509e-08, 1.174763e-08, 1.176137e-08, 1.177412e-08, 
    1.179928e-08, 1.183157e-08, 1.188823e-08, 1.193752e-08, 1.198251e-08, 
    1.197922e-08, 1.198038e-08, 1.199043e-08, 1.196553e-08, 1.199452e-08, 
    1.199938e-08, 1.198666e-08, 1.206048e-08, 1.203939e-08, 1.206097e-08, 
    1.204724e-08, 1.170204e-08, 1.171916e-08, 1.170991e-08, 1.17273e-08, 
    1.171505e-08, 1.176954e-08, 1.178587e-08, 1.186231e-08, 1.183094e-08, 
    1.188087e-08, 1.183601e-08, 1.184396e-08, 1.18825e-08, 1.183843e-08, 
    1.19348e-08, 1.186947e-08, 1.199082e-08, 1.192558e-08, 1.199491e-08, 
    1.198232e-08, 1.200316e-08, 1.202183e-08, 1.204532e-08, 1.208865e-08, 
    1.207862e-08, 1.211485e-08, 1.174467e-08, 1.176688e-08, 1.176492e-08, 
    1.178816e-08, 1.180534e-08, 1.184258e-08, 1.190232e-08, 1.187985e-08, 
    1.192109e-08, 1.192937e-08, 1.186672e-08, 1.190519e-08, 1.178174e-08, 
    1.180168e-08, 1.178981e-08, 1.174643e-08, 1.188503e-08, 1.18139e-08, 
    1.194525e-08, 1.190671e-08, 1.201917e-08, 1.196324e-08, 1.207309e-08, 
    1.212005e-08, 1.216424e-08, 1.221589e-08, 1.177899e-08, 1.176391e-08, 
    1.179092e-08, 1.182829e-08, 1.186297e-08, 1.190906e-08, 1.191378e-08, 
    1.192242e-08, 1.194478e-08, 1.196359e-08, 1.192515e-08, 1.196831e-08, 
    1.180631e-08, 1.189121e-08, 1.175821e-08, 1.179826e-08, 1.182609e-08, 
    1.181388e-08, 1.187729e-08, 1.189223e-08, 1.195296e-08, 1.192157e-08, 
    1.210846e-08, 1.202578e-08, 1.225522e-08, 1.21911e-08, 1.175864e-08, 
    1.177894e-08, 1.184961e-08, 1.181599e-08, 1.191214e-08, 1.193581e-08, 
    1.195505e-08, 1.197964e-08, 1.19823e-08, 1.199687e-08, 1.197299e-08, 
    1.199593e-08, 1.190916e-08, 1.194794e-08, 1.184153e-08, 1.186743e-08, 
    1.185552e-08, 1.184245e-08, 1.188278e-08, 1.192575e-08, 1.192667e-08, 
    1.194045e-08, 1.197928e-08, 1.191253e-08, 1.211914e-08, 1.199155e-08, 
    1.180108e-08, 1.18402e-08, 1.184578e-08, 1.183063e-08, 1.193344e-08, 
    1.189619e-08, 1.199652e-08, 1.19694e-08, 1.201383e-08, 1.199175e-08, 
    1.19885e-08, 1.196015e-08, 1.194249e-08, 1.189789e-08, 1.18616e-08, 
    1.183283e-08, 1.183952e-08, 1.187113e-08, 1.192838e-08, 1.198254e-08, 
    1.197068e-08, 1.201045e-08, 1.190517e-08, 1.194932e-08, 1.193225e-08, 
    1.197674e-08, 1.187926e-08, 1.196228e-08, 1.185804e-08, 1.186718e-08, 
    1.189545e-08, 1.195231e-08, 1.196489e-08, 1.197832e-08, 1.197003e-08, 
    1.192983e-08, 1.192325e-08, 1.189476e-08, 1.188689e-08, 1.186519e-08, 
    1.184721e-08, 1.186364e-08, 1.188088e-08, 1.192985e-08, 1.197398e-08, 
    1.20221e-08, 1.203387e-08, 1.209009e-08, 1.204433e-08, 1.211985e-08, 
    1.205565e-08, 1.216678e-08, 1.196709e-08, 1.205375e-08, 1.189673e-08, 
    1.191365e-08, 1.194425e-08, 1.201442e-08, 1.197654e-08, 1.202084e-08, 
    1.192299e-08, 1.187222e-08, 1.185908e-08, 1.183458e-08, 1.185964e-08, 
    1.185761e-08, 1.188159e-08, 1.187388e-08, 1.193148e-08, 1.190054e-08, 
    1.198842e-08, 1.202049e-08, 1.211106e-08, 1.216658e-08, 1.222309e-08, 
    1.224804e-08, 1.225563e-08, 1.22588e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382049e-10, 1.388128e-10, 1.386946e-10, 1.39185e-10, 1.38913e-10, 
    1.39234e-10, 1.383282e-10, 1.38837e-10, 1.385122e-10, 1.382596e-10, 
    1.401365e-10, 1.392068e-10, 1.411021e-10, 1.405092e-10, 1.419986e-10, 
    1.410098e-10, 1.421979e-10, 1.4197e-10, 1.426559e-10, 1.424594e-10, 
    1.433367e-10, 1.427466e-10, 1.437915e-10, 1.431958e-10, 1.43289e-10, 
    1.427271e-10, 1.393939e-10, 1.400208e-10, 1.393568e-10, 1.394461e-10, 
    1.39406e-10, 1.389186e-10, 1.386729e-10, 1.381585e-10, 1.382519e-10, 
    1.386297e-10, 1.394864e-10, 1.391956e-10, 1.399284e-10, 1.399118e-10, 
    1.407277e-10, 1.403598e-10, 1.417311e-10, 1.413414e-10, 1.424676e-10, 
    1.421844e-10, 1.424543e-10, 1.423724e-10, 1.424554e-10, 1.4204e-10, 
    1.422179e-10, 1.418524e-10, 1.404288e-10, 1.408472e-10, 1.395992e-10, 
    1.388489e-10, 1.383505e-10, 1.379968e-10, 1.380468e-10, 1.381421e-10, 
    1.386319e-10, 1.390925e-10, 1.394434e-10, 1.396782e-10, 1.399095e-10, 
    1.406096e-10, 1.409802e-10, 1.418099e-10, 1.416602e-10, 1.419139e-10, 
    1.421562e-10, 1.425631e-10, 1.424961e-10, 1.426753e-10, 1.419072e-10, 
    1.424177e-10, 1.415749e-10, 1.418054e-10, 1.399724e-10, 1.39274e-10, 
    1.389772e-10, 1.387174e-10, 1.380853e-10, 1.385218e-10, 1.383497e-10, 
    1.387591e-10, 1.390192e-10, 1.388906e-10, 1.396846e-10, 1.393759e-10, 
    1.410022e-10, 1.403017e-10, 1.421279e-10, 1.416909e-10, 1.422327e-10, 
    1.419562e-10, 1.424299e-10, 1.420036e-10, 1.427421e-10, 1.429029e-10, 
    1.42793e-10, 1.432151e-10, 1.4198e-10, 1.424543e-10, 1.388869e-10, 
    1.389079e-10, 1.390057e-10, 1.38576e-10, 1.385497e-10, 1.381559e-10, 
    1.385063e-10, 1.386555e-10, 1.390343e-10, 1.392583e-10, 1.394713e-10, 
    1.399396e-10, 1.404626e-10, 1.411939e-10, 1.417192e-10, 1.420714e-10, 
    1.418555e-10, 1.420461e-10, 1.41833e-10, 1.417331e-10, 1.428426e-10, 
    1.422196e-10, 1.431544e-10, 1.431026e-10, 1.426796e-10, 1.431085e-10, 
    1.389227e-10, 1.388019e-10, 1.383827e-10, 1.387108e-10, 1.38113e-10, 
    1.384476e-10, 1.3864e-10, 1.393823e-10, 1.395454e-10, 1.396967e-10, 
    1.399953e-10, 1.403787e-10, 1.410511e-10, 1.416362e-10, 1.421703e-10, 
    1.421311e-10, 1.421449e-10, 1.422642e-10, 1.419687e-10, 1.423128e-10, 
    1.423705e-10, 1.422195e-10, 1.430957e-10, 1.428454e-10, 1.431015e-10, 
    1.429385e-10, 1.388412e-10, 1.390443e-10, 1.389345e-10, 1.39141e-10, 
    1.389956e-10, 1.396423e-10, 1.398362e-10, 1.407435e-10, 1.403711e-10, 
    1.409638e-10, 1.404313e-10, 1.405257e-10, 1.409831e-10, 1.404601e-10, 
    1.41604e-10, 1.408285e-10, 1.422689e-10, 1.414945e-10, 1.423174e-10, 
    1.42168e-10, 1.424154e-10, 1.42637e-10, 1.429157e-10, 1.434301e-10, 
    1.43311e-10, 1.437412e-10, 1.393472e-10, 1.396108e-10, 1.395875e-10, 
    1.398633e-10, 1.400673e-10, 1.405094e-10, 1.412184e-10, 1.409517e-10, 
    1.414412e-10, 1.415395e-10, 1.407958e-10, 1.412524e-10, 1.397871e-10, 
    1.400239e-10, 1.398829e-10, 1.39368e-10, 1.410132e-10, 1.401689e-10, 
    1.417279e-10, 1.412706e-10, 1.426054e-10, 1.419416e-10, 1.432454e-10, 
    1.438029e-10, 1.443274e-10, 1.449405e-10, 1.397546e-10, 1.395755e-10, 
    1.398961e-10, 1.403397e-10, 1.407513e-10, 1.412984e-10, 1.413544e-10, 
    1.414569e-10, 1.417224e-10, 1.419457e-10, 1.414893e-10, 1.420016e-10, 
    1.400788e-10, 1.410865e-10, 1.395078e-10, 1.399832e-10, 1.403136e-10, 
    1.401686e-10, 1.409213e-10, 1.410986e-10, 1.418195e-10, 1.414468e-10, 
    1.436653e-10, 1.426838e-10, 1.454073e-10, 1.446462e-10, 1.39513e-10, 
    1.39754e-10, 1.405927e-10, 1.401936e-10, 1.41335e-10, 1.416159e-10, 
    1.418443e-10, 1.421362e-10, 1.421677e-10, 1.423407e-10, 1.420573e-10, 
    1.423295e-10, 1.412996e-10, 1.417598e-10, 1.404969e-10, 1.408043e-10, 
    1.406628e-10, 1.405077e-10, 1.409865e-10, 1.414965e-10, 1.415074e-10, 
    1.41671e-10, 1.421319e-10, 1.413396e-10, 1.43792e-10, 1.422775e-10, 
    1.400168e-10, 1.40481e-10, 1.405473e-10, 1.403675e-10, 1.415877e-10, 
    1.411456e-10, 1.423365e-10, 1.420146e-10, 1.42542e-10, 1.422799e-10, 
    1.422414e-10, 1.419048e-10, 1.416953e-10, 1.411659e-10, 1.407351e-10, 
    1.403935e-10, 1.40473e-10, 1.408482e-10, 1.415277e-10, 1.421706e-10, 
    1.420298e-10, 1.425019e-10, 1.412522e-10, 1.417762e-10, 1.415737e-10, 
    1.421018e-10, 1.409447e-10, 1.419301e-10, 1.406928e-10, 1.408013e-10, 
    1.411368e-10, 1.418118e-10, 1.419611e-10, 1.421206e-10, 1.420222e-10, 
    1.41545e-10, 1.414668e-10, 1.411287e-10, 1.410353e-10, 1.407776e-10, 
    1.405643e-10, 1.407592e-10, 1.409639e-10, 1.415452e-10, 1.42069e-10, 
    1.426401e-10, 1.427799e-10, 1.434472e-10, 1.42904e-10, 1.438005e-10, 
    1.430383e-10, 1.443576e-10, 1.419872e-10, 1.430159e-10, 1.411521e-10, 
    1.413529e-10, 1.417161e-10, 1.42549e-10, 1.420993e-10, 1.426252e-10, 
    1.414637e-10, 1.408611e-10, 1.407052e-10, 1.404143e-10, 1.407118e-10, 
    1.406876e-10, 1.409724e-10, 1.408809e-10, 1.415645e-10, 1.411973e-10, 
    1.422404e-10, 1.426211e-10, 1.436961e-10, 1.443551e-10, 1.450259e-10, 
    1.453221e-10, 1.454122e-10, 1.454499e-10 ;

 SOIL1N_vr =
  2.497419, 2.497412, 2.497414, 2.497408, 2.497411, 2.497408, 2.497418, 
    2.497412, 2.497416, 2.497419, 2.497398, 2.497408, 2.497387, 2.497394, 
    2.497377, 2.497388, 2.497375, 2.497377, 2.49737, 2.497372, 2.497362, 
    2.497369, 2.497357, 2.497364, 2.497363, 2.497369, 2.497406, 2.497399, 
    2.497406, 2.497405, 2.497406, 2.497411, 2.497414, 2.49742, 2.497419, 
    2.497414, 2.497405, 2.497408, 2.4974, 2.4974, 2.497391, 2.497395, 
    2.49738, 2.497384, 2.497372, 2.497375, 2.497372, 2.497373, 2.497372, 
    2.497377, 2.497375, 2.497379, 2.497395, 2.49739, 2.497404, 2.497412, 
    2.497417, 2.497422, 2.497421, 2.49742, 2.497414, 2.497409, 2.497405, 
    2.497403, 2.4974, 2.497392, 2.497388, 2.497379, 2.497381, 2.497378, 
    2.497375, 2.497371, 2.497372, 2.49737, 2.497378, 2.497372, 2.497382, 
    2.497379, 2.4974, 2.497407, 2.497411, 2.497413, 2.497421, 2.497416, 
    2.497417, 2.497413, 2.49741, 2.497411, 2.497403, 2.497406, 2.497388, 
    2.497396, 2.497376, 2.49738, 2.497375, 2.497378, 2.497372, 2.497377, 
    2.497369, 2.497367, 2.497368, 2.497364, 2.497377, 2.497372, 2.497411, 
    2.497411, 2.49741, 2.497415, 2.497415, 2.49742, 2.497416, 2.497414, 
    2.49741, 2.497407, 2.497405, 2.4974, 2.497394, 2.497386, 2.49738, 
    2.497376, 2.497379, 2.497377, 2.497379, 2.49738, 2.497368, 2.497375, 
    2.497364, 2.497365, 2.49737, 2.497365, 2.497411, 2.497412, 2.497417, 
    2.497414, 2.49742, 2.497416, 2.497414, 2.497406, 2.497404, 2.497403, 
    2.497399, 2.497395, 2.497388, 2.497381, 2.497375, 2.497376, 2.497375, 
    2.497374, 2.497377, 2.497374, 2.497373, 2.497375, 2.497365, 2.497368, 
    2.497365, 2.497367, 2.497412, 2.49741, 2.497411, 2.497409, 2.49741, 
    2.497403, 2.497401, 2.497391, 2.497395, 2.497389, 2.497395, 2.497393, 
    2.497388, 2.497394, 2.497381, 2.49739, 2.497374, 2.497383, 2.497374, 
    2.497375, 2.497373, 2.49737, 2.497367, 2.497361, 2.497363, 2.497358, 
    2.497406, 2.497404, 2.497404, 2.497401, 2.497398, 2.497394, 2.497386, 
    2.497389, 2.497383, 2.497382, 2.497391, 2.497385, 2.497401, 2.497399, 
    2.497401, 2.497406, 2.497388, 2.497397, 2.49738, 2.497385, 2.49737, 
    2.497378, 2.497363, 2.497357, 2.497351, 2.497345, 2.497402, 2.497404, 
    2.4974, 2.497396, 2.497391, 2.497385, 2.497384, 2.497383, 2.49738, 
    2.497378, 2.497383, 2.497377, 2.497398, 2.497387, 2.497405, 2.497399, 
    2.497396, 2.497397, 2.497389, 2.497387, 2.497379, 2.497383, 2.497359, 
    2.49737, 2.49734, 2.497348, 2.497405, 2.497402, 2.497393, 2.497397, 
    2.497385, 2.497381, 2.497379, 2.497375, 2.497375, 2.497373, 2.497376, 
    2.497374, 2.497385, 2.49738, 2.497394, 2.49739, 2.497392, 2.497394, 
    2.497388, 2.497383, 2.497383, 2.497381, 2.497376, 2.497384, 2.497357, 
    2.497374, 2.497399, 2.497394, 2.497393, 2.497395, 2.497382, 2.497386, 
    2.497373, 2.497377, 2.497371, 2.497374, 2.497375, 2.497378, 2.49738, 
    2.497386, 2.497391, 2.497395, 2.497394, 2.49739, 2.497382, 2.497375, 
    2.497377, 2.497372, 2.497385, 2.49738, 2.497382, 2.497376, 2.497389, 
    2.497378, 2.497391, 2.49739, 2.497387, 2.497379, 2.497378, 2.497376, 
    2.497377, 2.497382, 2.497383, 2.497387, 2.497388, 2.497391, 2.497393, 
    2.497391, 2.497389, 2.497382, 2.497376, 2.49737, 2.497369, 2.497361, 
    2.497367, 2.497357, 2.497366, 2.497351, 2.497377, 2.497366, 2.497386, 
    2.497384, 2.49738, 2.497371, 2.497376, 2.49737, 2.497383, 2.49739, 
    2.497391, 2.497395, 2.497391, 2.497392, 2.497388, 2.49739, 2.497382, 
    2.497386, 2.497375, 2.49737, 2.497358, 2.497351, 2.497344, 2.497341, 
    2.49734, 2.497339,
  2.497626, 2.497617, 2.497619, 2.497612, 2.497616, 2.497611, 2.497624, 
    2.497617, 2.497622, 2.497625, 2.497598, 2.497611, 2.497584, 2.497592, 
    2.497571, 2.497585, 2.497568, 2.497571, 2.497561, 2.497564, 2.497551, 
    2.49756, 2.497545, 2.497553, 2.497552, 2.49756, 2.497609, 2.497599, 
    2.497609, 2.497608, 2.497608, 2.497616, 2.497619, 2.497627, 2.497625, 
    2.49762, 2.497607, 2.497612, 2.497601, 2.497601, 2.497589, 2.497595, 
    2.497575, 2.49758, 2.497564, 2.497568, 2.497564, 2.497565, 2.497564, 
    2.49757, 2.497567, 2.497573, 2.497593, 2.497587, 2.497606, 2.497617, 
    2.497624, 2.497629, 2.497628, 2.497627, 2.49762, 2.497613, 2.497608, 
    2.497604, 2.497601, 2.497591, 2.497586, 2.497573, 2.497576, 2.497572, 
    2.497568, 2.497562, 2.497563, 2.497561, 2.497572, 2.497565, 2.497577, 
    2.497573, 2.4976, 2.49761, 2.497615, 2.497618, 2.497628, 2.497621, 
    2.497624, 2.497618, 2.497614, 2.497616, 2.497604, 2.497609, 2.497585, 
    2.497595, 2.497569, 2.497575, 2.497567, 2.497571, 2.497564, 2.497571, 
    2.49756, 2.497558, 2.497559, 2.497553, 2.497571, 2.497564, 2.497616, 
    2.497616, 2.497614, 2.497621, 2.497621, 2.497627, 2.497622, 2.497619, 
    2.497614, 2.497611, 2.497607, 2.497601, 2.497593, 2.497582, 2.497575, 
    2.49757, 2.497573, 2.49757, 2.497573, 2.497575, 2.497558, 2.497567, 
    2.497554, 2.497555, 2.497561, 2.497555, 2.497615, 2.497617, 2.497623, 
    2.497618, 2.497627, 2.497622, 2.49762, 2.497609, 2.497606, 2.497604, 
    2.4976, 2.497594, 2.497584, 2.497576, 2.497568, 2.497569, 2.497569, 
    2.497567, 2.497571, 2.497566, 2.497565, 2.497567, 2.497555, 2.497558, 
    2.497555, 2.497557, 2.497617, 2.497614, 2.497615, 2.497612, 2.497614, 
    2.497605, 2.497602, 2.497589, 2.497594, 2.497586, 2.497593, 2.497592, 
    2.497586, 2.497593, 2.497576, 2.497588, 2.497567, 2.497578, 2.497566, 
    2.497568, 2.497565, 2.497561, 2.497557, 2.49755, 2.497552, 2.497545, 
    2.497609, 2.497605, 2.497606, 2.497602, 2.497599, 2.497592, 2.497582, 
    2.497586, 2.497579, 2.497577, 2.497588, 2.497581, 2.497603, 2.497599, 
    2.497602, 2.497609, 2.497585, 2.497597, 2.497575, 2.497581, 2.497562, 
    2.497571, 2.497553, 2.497545, 2.497537, 2.497528, 2.497603, 2.497606, 
    2.497601, 2.497595, 2.497589, 2.497581, 2.49758, 2.497579, 2.497575, 
    2.497571, 2.497578, 2.497571, 2.497599, 2.497584, 2.497607, 2.4976, 
    2.497595, 2.497597, 2.497586, 2.497584, 2.497573, 2.497579, 2.497546, 
    2.497561, 2.497521, 2.497532, 2.497607, 2.497603, 2.497591, 2.497597, 
    2.49758, 2.497576, 2.497573, 2.497569, 2.497568, 2.497566, 2.49757, 
    2.497566, 2.497581, 2.497574, 2.497592, 2.497588, 2.49759, 2.497592, 
    2.497585, 2.497578, 2.497578, 2.497576, 2.497569, 2.49758, 2.497545, 
    2.497567, 2.4976, 2.497593, 2.497592, 2.497594, 2.497577, 2.497583, 
    2.497566, 2.497571, 2.497563, 2.497567, 2.497567, 2.497572, 2.497575, 
    2.497583, 2.497589, 2.497594, 2.497593, 2.497587, 2.497577, 2.497568, 
    2.49757, 2.497563, 2.497581, 2.497574, 2.497577, 2.497569, 2.497586, 
    2.497572, 2.49759, 2.497588, 2.497583, 2.497573, 2.497571, 2.497569, 
    2.49757, 2.497577, 2.497578, 2.497583, 2.497585, 2.497588, 2.497591, 
    2.497589, 2.497586, 2.497577, 2.49757, 2.497561, 2.497559, 2.49755, 
    2.497558, 2.497545, 2.497555, 2.497536, 2.497571, 2.497556, 2.497583, 
    2.49758, 2.497575, 2.497563, 2.497569, 2.497562, 2.497578, 2.497587, 
    2.497589, 2.497594, 2.497589, 2.49759, 2.497586, 2.497587, 2.497577, 
    2.497582, 2.497567, 2.497562, 2.497546, 2.497536, 2.497527, 2.497523, 
    2.497521, 2.497521,
  2.497841, 2.497832, 2.497833, 2.497826, 2.49783, 2.497825, 2.497839, 
    2.497831, 2.497836, 2.49784, 2.497811, 2.497825, 2.497796, 2.497805, 
    2.497782, 2.497797, 2.497779, 2.497782, 2.497772, 2.497775, 2.497761, 
    2.49777, 2.497754, 2.497763, 2.497762, 2.497771, 2.497823, 2.497813, 
    2.497823, 2.497822, 2.497822, 2.49783, 2.497834, 2.497842, 2.49784, 
    2.497834, 2.497821, 2.497826, 2.497814, 2.497814, 2.497802, 2.497808, 
    2.497786, 2.497792, 2.497775, 2.497779, 2.497775, 2.497776, 2.497775, 
    2.497781, 2.497779, 2.497784, 2.497806, 2.4978, 2.497819, 2.497831, 
    2.497839, 2.497844, 2.497844, 2.497842, 2.497834, 2.497827, 2.497822, 
    2.497818, 2.497814, 2.497804, 2.497798, 2.497785, 2.497787, 2.497783, 
    2.49778, 2.497773, 2.497774, 2.497772, 2.497783, 2.497776, 2.497789, 
    2.497785, 2.497813, 2.497824, 2.497829, 2.497833, 2.497843, 2.497836, 
    2.497839, 2.497832, 2.497828, 2.49783, 2.497818, 2.497823, 2.497797, 
    2.497808, 2.49778, 2.497787, 2.497778, 2.497783, 2.497775, 2.497782, 
    2.497771, 2.497768, 2.49777, 2.497763, 2.497782, 2.497775, 2.49783, 
    2.49783, 2.497828, 2.497835, 2.497836, 2.497842, 2.497836, 2.497834, 
    2.497828, 2.497825, 2.497821, 2.497814, 2.497806, 2.497794, 2.497786, 
    2.497781, 2.497784, 2.497781, 2.497785, 2.497786, 2.497769, 2.497779, 
    2.497764, 2.497765, 2.497772, 2.497765, 2.49783, 2.497832, 2.497838, 
    2.497833, 2.497843, 2.497837, 2.497834, 2.497823, 2.49782, 2.497818, 
    2.497813, 2.497807, 2.497797, 2.497788, 2.497779, 2.49778, 2.49778, 
    2.497778, 2.497782, 2.497777, 2.497776, 2.497779, 2.497765, 2.497769, 
    2.497765, 2.497767, 2.497831, 2.497828, 2.49783, 2.497826, 2.497829, 
    2.497819, 2.497816, 2.497802, 2.497807, 2.497798, 2.497806, 2.497805, 
    2.497798, 2.497806, 2.497788, 2.4978, 2.497778, 2.49779, 2.497777, 
    2.497779, 2.497776, 2.497772, 2.497768, 2.49776, 2.497762, 2.497755, 
    2.497823, 2.497819, 2.497819, 2.497815, 2.497812, 2.497805, 2.497794, 
    2.497798, 2.497791, 2.497789, 2.497801, 2.497794, 2.497816, 2.497813, 
    2.497815, 2.497823, 2.497797, 2.49781, 2.497786, 2.497793, 2.497773, 
    2.497783, 2.497763, 2.497754, 2.497746, 2.497736, 2.497817, 2.49782, 
    2.497815, 2.497808, 2.497801, 2.497793, 2.497792, 2.49779, 2.497786, 
    2.497783, 2.49779, 2.497782, 2.497812, 2.497796, 2.497821, 2.497813, 
    2.497808, 2.49781, 2.497799, 2.497796, 2.497785, 2.497791, 2.497756, 
    2.497771, 2.497729, 2.497741, 2.497821, 2.497817, 2.497804, 2.49781, 
    2.497792, 2.497788, 2.497784, 2.49778, 2.497779, 2.497777, 2.497781, 
    2.497777, 2.497793, 2.497786, 2.497805, 2.497801, 2.497803, 2.497805, 
    2.497798, 2.49779, 2.49779, 2.497787, 2.49778, 2.497792, 2.497754, 
    2.497778, 2.497813, 2.497806, 2.497805, 2.497807, 2.497788, 2.497795, 
    2.497777, 2.497782, 2.497774, 2.497778, 2.497778, 2.497783, 2.497787, 
    2.497795, 2.497802, 2.497807, 2.497806, 2.4978, 2.497789, 2.497779, 
    2.497782, 2.497774, 2.497794, 2.497786, 2.497789, 2.49778, 2.497798, 
    2.497783, 2.497802, 2.497801, 2.497795, 2.497785, 2.497783, 2.49778, 
    2.497782, 2.497789, 2.49779, 2.497796, 2.497797, 2.497801, 2.497804, 
    2.497801, 2.497798, 2.497789, 2.497781, 2.497772, 2.49777, 2.49776, 
    2.497768, 2.497754, 2.497766, 2.497746, 2.497782, 2.497766, 2.497795, 
    2.497792, 2.497786, 2.497773, 2.497781, 2.497772, 2.49779, 2.4978, 
    2.497802, 2.497807, 2.497802, 2.497802, 2.497798, 2.497799, 2.497789, 
    2.497794, 2.497778, 2.497772, 2.497756, 2.497746, 2.497735, 2.49773, 
    2.497729, 2.497729,
  2.498013, 2.498003, 2.498005, 2.497998, 2.498002, 2.497997, 2.498011, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.49797, 2.497951, 2.497955, 2.497944, 2.497947, 2.497934, 
    2.497943, 2.497927, 2.497936, 2.497934, 2.497943, 2.497994, 2.497985, 
    2.497995, 2.497994, 2.497994, 2.498002, 2.498006, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497998, 2.497986, 2.497987, 2.497974, 2.49798, 
    2.497958, 2.497964, 2.497947, 2.497952, 2.497947, 2.497948, 2.497947, 
    2.497954, 2.497951, 2.497957, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.498011, 2.498016, 2.498015, 2.498014, 2.498006, 2.497999, 2.497994, 
    2.49799, 2.497987, 2.497976, 2.49797, 2.497957, 2.49796, 2.497956, 
    2.497952, 2.497946, 2.497947, 2.497944, 2.497956, 2.497948, 2.497961, 
    2.497957, 2.497986, 2.497996, 2.498001, 2.498005, 2.498015, 2.498008, 
    2.498011, 2.498004, 2.498, 2.498002, 2.49799, 2.497995, 2.49797, 2.49798, 
    2.497952, 2.497959, 2.497951, 2.497955, 2.497948, 2.497954, 2.497943, 
    2.49794, 2.497942, 2.497936, 2.497955, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498008, 2.498013, 2.498008, 2.498006, 2.498, 2.497997, 
    2.497993, 2.497986, 2.497978, 2.497967, 2.497959, 2.497953, 2.497957, 
    2.497954, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497944, 2.497937, 2.498002, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497995, 2.497992, 2.49799, 2.497985, 2.497979, 
    2.497969, 2.49796, 2.497952, 2.497952, 2.497952, 2.49795, 2.497955, 
    2.497949, 2.497949, 2.497951, 2.497937, 2.497941, 2.497937, 2.49794, 
    2.498003, 2.498, 2.498002, 2.497998, 2.498001, 2.497991, 2.497988, 
    2.497974, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497978, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497952, 2.497948, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497992, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497963, 
    2.497961, 2.497973, 2.497966, 2.497988, 2.497985, 2.497987, 2.497995, 
    2.497969, 2.497983, 2.497958, 2.497966, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497989, 2.497992, 2.497987, 2.49798, 
    2.497973, 2.497965, 2.497964, 2.497963, 2.497959, 2.497955, 2.497962, 
    2.497954, 2.497984, 2.497968, 2.497993, 2.497985, 2.49798, 2.497983, 
    2.497971, 2.497968, 2.497957, 2.497963, 2.497929, 2.497944, 2.497902, 
    2.497914, 2.497993, 2.497989, 2.497976, 2.497982, 2.497965, 2.49796, 
    2.497957, 2.497952, 2.497952, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497958, 2.497977, 2.497973, 2.497975, 2.497977, 2.49797, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497927, 2.49795, 2.497985, 
    2.497978, 2.497977, 2.497979, 2.497961, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.497951, 2.497956, 2.497959, 2.497967, 2.497974, 
    2.497979, 2.497978, 2.497972, 2.497962, 2.497952, 2.497954, 2.497947, 
    2.497966, 2.497958, 2.497961, 2.497953, 2.497971, 2.497955, 2.497974, 
    2.497973, 2.497967, 2.497957, 2.497955, 2.497952, 2.497954, 2.497961, 
    2.497962, 2.497968, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497932, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497939, 2.497967, 2.497964, 2.497959, 
    2.497946, 2.497953, 2.497945, 2.497962, 2.497972, 2.497974, 2.497979, 
    2.497974, 2.497974, 2.49797, 2.497972, 2.497961, 2.497967, 2.497951, 
    2.497945, 2.497928, 2.497918, 2.497908, 2.497903, 2.497902, 2.497901,
  2.498213, 2.498205, 2.498207, 2.4982, 2.498204, 2.498199, 2.498212, 
    2.498205, 2.498209, 2.498213, 2.498187, 2.498199, 2.498174, 2.498182, 
    2.498161, 2.498175, 2.498159, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498144, 2.498151, 2.498197, 2.498188, 
    2.498198, 2.498196, 2.498197, 2.498204, 2.498207, 2.498214, 2.498213, 
    2.498207, 2.498196, 2.4982, 2.49819, 2.49819, 2.498179, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498163, 
    2.498159, 2.498154, 2.498154, 2.498152, 2.498163, 2.498156, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498206, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498185, 2.49816, 2.498166, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498145, 2.498162, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498209, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498164, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498204, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498189, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498184, 2.498175, 2.498183, 2.498182, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498156, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.498191, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498172, 2.498192, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498137, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498169, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498174, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498115, 2.498125, 2.498195, 2.498192, 2.498181, 2.498186, 
    2.49817, 2.498167, 2.498163, 2.498159, 2.498159, 2.498157, 2.498161, 
    2.498157, 2.498171, 2.498165, 2.498182, 2.498178, 2.49818, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498158, 2.498188, 2.498182, 2.498181, 2.498184, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498158, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498179, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498172, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.49816, 
    2.498161, 2.498168, 2.498169, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498168, 2.49816, 2.498152, 2.498151, 2.498142, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498162, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498153, 2.498169, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.138626e-08, 6.165622e-08, 6.160374e-08, 6.182147e-08, 6.170069e-08, 
    6.184327e-08, 6.144099e-08, 6.166694e-08, 6.15227e-08, 6.141056e-08, 
    6.224403e-08, 6.183119e-08, 6.267283e-08, 6.240955e-08, 6.307092e-08, 
    6.263187e-08, 6.315945e-08, 6.305824e-08, 6.336283e-08, 6.327556e-08, 
    6.366515e-08, 6.340309e-08, 6.386709e-08, 6.360256e-08, 6.364395e-08, 
    6.339445e-08, 6.191426e-08, 6.219263e-08, 6.189777e-08, 6.193746e-08, 
    6.191966e-08, 6.170318e-08, 6.15941e-08, 6.136563e-08, 6.14071e-08, 
    6.157491e-08, 6.195532e-08, 6.182618e-08, 6.215162e-08, 6.214427e-08, 
    6.250657e-08, 6.234322e-08, 6.295216e-08, 6.277909e-08, 6.327921e-08, 
    6.315344e-08, 6.32733e-08, 6.323695e-08, 6.327377e-08, 6.308932e-08, 
    6.316835e-08, 6.300603e-08, 6.237381e-08, 6.255962e-08, 6.200545e-08, 
    6.167224e-08, 6.14509e-08, 6.129384e-08, 6.131604e-08, 6.135837e-08, 
    6.157589e-08, 6.17804e-08, 6.193624e-08, 6.204049e-08, 6.214322e-08, 
    6.245415e-08, 6.26187e-08, 6.298716e-08, 6.292066e-08, 6.303331e-08, 
    6.314092e-08, 6.33216e-08, 6.329186e-08, 6.337147e-08, 6.303033e-08, 
    6.325705e-08, 6.288278e-08, 6.298515e-08, 6.217116e-08, 6.186102e-08, 
    6.172921e-08, 6.161383e-08, 6.133311e-08, 6.152697e-08, 6.145055e-08, 
    6.163235e-08, 6.174787e-08, 6.169073e-08, 6.204335e-08, 6.190626e-08, 
    6.262845e-08, 6.231738e-08, 6.312837e-08, 6.29343e-08, 6.317489e-08, 
    6.305212e-08, 6.326247e-08, 6.307316e-08, 6.340109e-08, 6.34725e-08, 
    6.34237e-08, 6.361115e-08, 6.306266e-08, 6.32733e-08, 6.168914e-08, 
    6.169845e-08, 6.174186e-08, 6.155104e-08, 6.153937e-08, 6.136449e-08, 
    6.152009e-08, 6.158636e-08, 6.175456e-08, 6.185406e-08, 6.194864e-08, 
    6.215659e-08, 6.238884e-08, 6.271359e-08, 6.294689e-08, 6.310327e-08, 
    6.300738e-08, 6.309205e-08, 6.29974e-08, 6.295304e-08, 6.344575e-08, 
    6.316909e-08, 6.358418e-08, 6.356122e-08, 6.337336e-08, 6.35638e-08, 
    6.170499e-08, 6.165137e-08, 6.14652e-08, 6.16109e-08, 6.134544e-08, 
    6.149403e-08, 6.157947e-08, 6.190913e-08, 6.198155e-08, 6.204871e-08, 
    6.218136e-08, 6.235158e-08, 6.265019e-08, 6.291001e-08, 6.314718e-08, 
    6.31298e-08, 6.313592e-08, 6.318891e-08, 6.305766e-08, 6.321046e-08, 
    6.32361e-08, 6.316905e-08, 6.355814e-08, 6.344698e-08, 6.356073e-08, 
    6.348835e-08, 6.16688e-08, 6.175902e-08, 6.171027e-08, 6.180196e-08, 
    6.173737e-08, 6.202458e-08, 6.211068e-08, 6.251359e-08, 6.234824e-08, 
    6.26114e-08, 6.237497e-08, 6.241686e-08, 6.262e-08, 6.238774e-08, 
    6.289569e-08, 6.255132e-08, 6.319097e-08, 6.28471e-08, 6.321252e-08, 
    6.314615e-08, 6.325602e-08, 6.335443e-08, 6.347822e-08, 6.370664e-08, 
    6.365374e-08, 6.384476e-08, 6.189354e-08, 6.201056e-08, 6.200026e-08, 
    6.212273e-08, 6.22133e-08, 6.240961e-08, 6.272446e-08, 6.260606e-08, 
    6.282342e-08, 6.286705e-08, 6.253683e-08, 6.273959e-08, 6.208889e-08, 
    6.219403e-08, 6.213142e-08, 6.190277e-08, 6.263335e-08, 6.225842e-08, 
    6.295075e-08, 6.274764e-08, 6.33404e-08, 6.304561e-08, 6.362463e-08, 
    6.387216e-08, 6.41051e-08, 6.437735e-08, 6.207443e-08, 6.199491e-08, 
    6.213729e-08, 6.233429e-08, 6.251705e-08, 6.276003e-08, 6.278488e-08, 
    6.283041e-08, 6.294831e-08, 6.304744e-08, 6.28448e-08, 6.30723e-08, 
    6.221842e-08, 6.266589e-08, 6.196485e-08, 6.217596e-08, 6.232267e-08, 
    6.225831e-08, 6.259253e-08, 6.26713e-08, 6.29914e-08, 6.282593e-08, 
    6.381107e-08, 6.337522e-08, 6.458463e-08, 6.424666e-08, 6.196713e-08, 
    6.207416e-08, 6.244665e-08, 6.226941e-08, 6.277624e-08, 6.2901e-08, 
    6.300241e-08, 6.313206e-08, 6.314605e-08, 6.322286e-08, 6.309699e-08, 
    6.321789e-08, 6.276054e-08, 6.296492e-08, 6.240406e-08, 6.254058e-08, 
    6.247777e-08, 6.240889e-08, 6.262149e-08, 6.2848e-08, 6.285283e-08, 
    6.292546e-08, 6.313014e-08, 6.27783e-08, 6.386734e-08, 6.319479e-08, 
    6.219086e-08, 6.239702e-08, 6.242645e-08, 6.23466e-08, 6.28885e-08, 
    6.269214e-08, 6.322099e-08, 6.307806e-08, 6.331224e-08, 6.319588e-08, 
    6.317875e-08, 6.302929e-08, 6.293624e-08, 6.270115e-08, 6.250987e-08, 
    6.235818e-08, 6.239345e-08, 6.256008e-08, 6.286185e-08, 6.314732e-08, 
    6.308479e-08, 6.329444e-08, 6.27395e-08, 6.29722e-08, 6.288226e-08, 
    6.311677e-08, 6.260291e-08, 6.304052e-08, 6.249106e-08, 6.253924e-08, 
    6.268825e-08, 6.298799e-08, 6.305429e-08, 6.31251e-08, 6.308141e-08, 
    6.286951e-08, 6.283479e-08, 6.268463e-08, 6.264317e-08, 6.252875e-08, 
    6.243402e-08, 6.252057e-08, 6.261147e-08, 6.28696e-08, 6.310221e-08, 
    6.335583e-08, 6.341789e-08, 6.371423e-08, 6.347301e-08, 6.387109e-08, 
    6.353267e-08, 6.411849e-08, 6.306586e-08, 6.35227e-08, 6.269503e-08, 
    6.27842e-08, 6.294547e-08, 6.331538e-08, 6.311567e-08, 6.334922e-08, 
    6.283343e-08, 6.256583e-08, 6.249658e-08, 6.236741e-08, 6.249954e-08, 
    6.248879e-08, 6.261523e-08, 6.257459e-08, 6.287816e-08, 6.27151e-08, 
    6.317833e-08, 6.334737e-08, 6.382474e-08, 6.411739e-08, 6.441527e-08, 
    6.454679e-08, 6.458681e-08, 6.460355e-08 ;

 SOIL1_HR_S3 =
  7.28467e-10, 7.316718e-10, 7.310487e-10, 7.336336e-10, 7.321997e-10, 
    7.338923e-10, 7.291167e-10, 7.31799e-10, 7.300867e-10, 7.287554e-10, 
    7.386501e-10, 7.33749e-10, 7.437408e-10, 7.406151e-10, 7.48467e-10, 
    7.432545e-10, 7.495179e-10, 7.483165e-10, 7.519325e-10, 7.508966e-10, 
    7.555219e-10, 7.524106e-10, 7.579194e-10, 7.547788e-10, 7.552701e-10, 
    7.52308e-10, 7.347352e-10, 7.3804e-10, 7.345394e-10, 7.350107e-10, 
    7.347992e-10, 7.322293e-10, 7.309344e-10, 7.28222e-10, 7.287144e-10, 
    7.307065e-10, 7.352225e-10, 7.336895e-10, 7.37553e-10, 7.374658e-10, 
    7.41767e-10, 7.398276e-10, 7.47057e-10, 7.450023e-10, 7.509398e-10, 
    7.494466e-10, 7.508696e-10, 7.504382e-10, 7.508753e-10, 7.486853e-10, 
    7.496236e-10, 7.476965e-10, 7.401909e-10, 7.423968e-10, 7.358177e-10, 
    7.31862e-10, 7.292343e-10, 7.273698e-10, 7.276334e-10, 7.281359e-10, 
    7.307182e-10, 7.331459e-10, 7.349961e-10, 7.362337e-10, 7.374532e-10, 
    7.411446e-10, 7.430981e-10, 7.474725e-10, 7.46683e-10, 7.480204e-10, 
    7.49298e-10, 7.514431e-10, 7.5109e-10, 7.520351e-10, 7.479851e-10, 
    7.506767e-10, 7.462333e-10, 7.474486e-10, 7.377851e-10, 7.341031e-10, 
    7.325384e-10, 7.311685e-10, 7.278361e-10, 7.301374e-10, 7.292302e-10, 
    7.313884e-10, 7.327598e-10, 7.320815e-10, 7.362676e-10, 7.346402e-10, 
    7.432139e-10, 7.395209e-10, 7.49149e-10, 7.46845e-10, 7.497012e-10, 
    7.482437e-10, 7.507411e-10, 7.484935e-10, 7.523868e-10, 7.532346e-10, 
    7.526553e-10, 7.548807e-10, 7.483689e-10, 7.508697e-10, 7.320625e-10, 
    7.321732e-10, 7.326885e-10, 7.304232e-10, 7.302846e-10, 7.282085e-10, 
    7.300557e-10, 7.308424e-10, 7.328393e-10, 7.340205e-10, 7.351433e-10, 
    7.37612e-10, 7.403692e-10, 7.442246e-10, 7.469944e-10, 7.48851e-10, 
    7.477126e-10, 7.487177e-10, 7.47594e-10, 7.470674e-10, 7.52917e-10, 
    7.496324e-10, 7.545606e-10, 7.542879e-10, 7.520576e-10, 7.543186e-10, 
    7.322508e-10, 7.316142e-10, 7.294041e-10, 7.311337e-10, 7.279824e-10, 
    7.297464e-10, 7.307607e-10, 7.346743e-10, 7.35534e-10, 7.363313e-10, 
    7.37906e-10, 7.399269e-10, 7.434721e-10, 7.465565e-10, 7.493723e-10, 
    7.49166e-10, 7.492387e-10, 7.498677e-10, 7.483095e-10, 7.501235e-10, 
    7.50428e-10, 7.49632e-10, 7.542513e-10, 7.529316e-10, 7.54282e-10, 
    7.534228e-10, 7.318212e-10, 7.328923e-10, 7.323135e-10, 7.334019e-10, 
    7.326351e-10, 7.360447e-10, 7.37067e-10, 7.418503e-10, 7.398872e-10, 
    7.430114e-10, 7.402045e-10, 7.407019e-10, 7.431135e-10, 7.403562e-10, 
    7.463866e-10, 7.422983e-10, 7.498921e-10, 7.458097e-10, 7.50148e-10, 
    7.493601e-10, 7.506645e-10, 7.518328e-10, 7.533025e-10, 7.560144e-10, 
    7.553864e-10, 7.576543e-10, 7.344891e-10, 7.358785e-10, 7.357561e-10, 
    7.3721e-10, 7.382853e-10, 7.406158e-10, 7.443537e-10, 7.429481e-10, 
    7.455285e-10, 7.460466e-10, 7.421262e-10, 7.445333e-10, 7.368082e-10, 
    7.380564e-10, 7.373132e-10, 7.345987e-10, 7.432721e-10, 7.388209e-10, 
    7.470402e-10, 7.446289e-10, 7.516662e-10, 7.481665e-10, 7.550407e-10, 
    7.579796e-10, 7.607452e-10, 7.639777e-10, 7.366366e-10, 7.356926e-10, 
    7.373829e-10, 7.397216e-10, 7.418913e-10, 7.44776e-10, 7.450711e-10, 
    7.456115e-10, 7.470113e-10, 7.481882e-10, 7.457824e-10, 7.484833e-10, 
    7.38346e-10, 7.436584e-10, 7.353358e-10, 7.37842e-10, 7.395837e-10, 
    7.388196e-10, 7.427874e-10, 7.437226e-10, 7.475229e-10, 7.455583e-10, 
    7.572543e-10, 7.520797e-10, 7.664386e-10, 7.624259e-10, 7.353628e-10, 
    7.366334e-10, 7.410555e-10, 7.389515e-10, 7.449685e-10, 7.464496e-10, 
    7.476536e-10, 7.491928e-10, 7.493589e-10, 7.502708e-10, 7.487764e-10, 
    7.502118e-10, 7.447821e-10, 7.472085e-10, 7.4055e-10, 7.421707e-10, 
    7.41425e-10, 7.406072e-10, 7.431312e-10, 7.458203e-10, 7.458777e-10, 
    7.467399e-10, 7.4917e-10, 7.449928e-10, 7.579224e-10, 7.499376e-10, 
    7.380189e-10, 7.404664e-10, 7.408158e-10, 7.398677e-10, 7.463011e-10, 
    7.439701e-10, 7.502486e-10, 7.485517e-10, 7.51332e-10, 7.499504e-10, 
    7.497472e-10, 7.479727e-10, 7.46868e-10, 7.44077e-10, 7.418061e-10, 
    7.400052e-10, 7.404239e-10, 7.424021e-10, 7.459848e-10, 7.49374e-10, 
    7.486315e-10, 7.511207e-10, 7.445322e-10, 7.472949e-10, 7.462272e-10, 
    7.490113e-10, 7.429107e-10, 7.48106e-10, 7.415829e-10, 7.421547e-10, 
    7.439238e-10, 7.474824e-10, 7.482695e-10, 7.491102e-10, 7.485914e-10, 
    7.460758e-10, 7.456635e-10, 7.438808e-10, 7.433886e-10, 7.420302e-10, 
    7.409056e-10, 7.419331e-10, 7.430123e-10, 7.460768e-10, 7.488384e-10, 
    7.518495e-10, 7.525863e-10, 7.561046e-10, 7.532407e-10, 7.579669e-10, 
    7.539489e-10, 7.609041e-10, 7.484069e-10, 7.538306e-10, 7.440043e-10, 
    7.450628e-10, 7.469776e-10, 7.513691e-10, 7.489982e-10, 7.517709e-10, 
    7.456474e-10, 7.424704e-10, 7.416484e-10, 7.401147e-10, 7.416834e-10, 
    7.415558e-10, 7.430569e-10, 7.425745e-10, 7.461785e-10, 7.442426e-10, 
    7.49742e-10, 7.51749e-10, 7.574166e-10, 7.608911e-10, 7.644279e-10, 
    7.659893e-10, 7.664646e-10, 7.666632e-10 ;

 SOIL2C =
  5.784044, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784102, 5.784096, 5.784097, 5.784091, 5.784057, 5.784063, 
    5.784057, 5.784057, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.78407, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784084, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784057, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784088, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784052, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784051, 5.78406, 5.784057, 5.784073, 
    5.784066, 5.784085, 5.784081, 5.784086, 5.784083, 5.784089, 5.784084, 
    5.784091, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784051, 
    5.784052, 5.784053, 5.784048, 5.784048, 5.784044, 5.784048, 5.784049, 
    5.784053, 5.784055, 5.784058, 5.784062, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784084, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784095, 5.784091, 5.784095, 5.784052, 5.78405, 5.784046, 
    5.78405, 5.784043, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.78408, 5.784086, 5.784085, 5.784085, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784095, 5.784093, 
    5.784095, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784087, 
    5.784086, 5.784088, 5.784091, 5.784093, 5.784099, 5.784098, 5.784102, 
    5.784056, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.784079, 5.784071, 5.784076, 5.784061, 5.784063, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784076, 5.78409, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784114, 5.78406, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784077, 5.784078, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784074, 5.784058, 5.784063, 
    5.784066, 5.784065, 5.784073, 5.784075, 5.784082, 5.784078, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.78406, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784085, 5.784086, 5.784088, 5.784084, 
    5.784087, 5.784077, 5.784081, 5.784068, 5.784071, 5.78407, 5.784069, 
    5.784073, 5.784079, 5.784079, 5.784081, 5.784085, 5.784077, 5.784102, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784067, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.784089, 5.784076, 5.784081, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784083, 5.784085, 
    5.784084, 5.784079, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.784079, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784094, 5.784075, 
    5.784077, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.78407, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784086, 5.784091, 5.784101, 5.784109, 5.784115, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086043e-09, 1.090822e-09, 1.089893e-09, 1.093748e-09, 1.09161e-09, 
    1.094134e-09, 1.087011e-09, 1.091012e-09, 1.088458e-09, 1.086473e-09, 
    1.10123e-09, 1.09392e-09, 1.108822e-09, 1.10416e-09, 1.11587e-09, 
    1.108096e-09, 1.117437e-09, 1.115646e-09, 1.121038e-09, 1.119493e-09, 
    1.126391e-09, 1.121751e-09, 1.129967e-09, 1.125283e-09, 1.126016e-09, 
    1.121598e-09, 1.095391e-09, 1.10032e-09, 1.095099e-09, 1.095802e-09, 
    1.095486e-09, 1.091654e-09, 1.089722e-09, 1.085677e-09, 1.086412e-09, 
    1.089383e-09, 1.096118e-09, 1.093831e-09, 1.099593e-09, 1.099463e-09, 
    1.105878e-09, 1.102986e-09, 1.113767e-09, 1.110703e-09, 1.119558e-09, 
    1.117331e-09, 1.119453e-09, 1.11881e-09, 1.119462e-09, 1.116196e-09, 
    1.117595e-09, 1.114721e-09, 1.103527e-09, 1.106817e-09, 1.097005e-09, 
    1.091106e-09, 1.087187e-09, 1.084406e-09, 1.084799e-09, 1.085549e-09, 
    1.0894e-09, 1.093021e-09, 1.09578e-09, 1.097626e-09, 1.099445e-09, 
    1.10495e-09, 1.107863e-09, 1.114387e-09, 1.11321e-09, 1.115204e-09, 
    1.11711e-09, 1.120309e-09, 1.119782e-09, 1.121191e-09, 1.115151e-09, 
    1.119166e-09, 1.112539e-09, 1.114351e-09, 1.099939e-09, 1.094448e-09, 
    1.092115e-09, 1.090072e-09, 1.085102e-09, 1.088534e-09, 1.087181e-09, 
    1.0904e-09, 1.092445e-09, 1.091433e-09, 1.097676e-09, 1.095249e-09, 
    1.108036e-09, 1.102528e-09, 1.116887e-09, 1.113451e-09, 1.117711e-09, 
    1.115537e-09, 1.119262e-09, 1.11591e-09, 1.121716e-09, 1.12298e-09, 
    1.122116e-09, 1.125435e-09, 1.115724e-09, 1.119453e-09, 1.091405e-09, 
    1.09157e-09, 1.092339e-09, 1.08896e-09, 1.088753e-09, 1.085657e-09, 
    1.088412e-09, 1.089585e-09, 1.092563e-09, 1.094325e-09, 1.096e-09, 
    1.099681e-09, 1.103794e-09, 1.109543e-09, 1.113674e-09, 1.116443e-09, 
    1.114745e-09, 1.116244e-09, 1.114568e-09, 1.113783e-09, 1.122507e-09, 
    1.117608e-09, 1.124958e-09, 1.124551e-09, 1.121225e-09, 1.124597e-09, 
    1.091686e-09, 1.090736e-09, 1.08744e-09, 1.09002e-09, 1.08532e-09, 
    1.087951e-09, 1.089463e-09, 1.0953e-09, 1.096582e-09, 1.097771e-09, 
    1.10012e-09, 1.103134e-09, 1.108421e-09, 1.113021e-09, 1.11722e-09, 
    1.116913e-09, 1.117021e-09, 1.117959e-09, 1.115635e-09, 1.118341e-09, 
    1.118795e-09, 1.117607e-09, 1.124496e-09, 1.122528e-09, 1.124542e-09, 
    1.123261e-09, 1.091045e-09, 1.092643e-09, 1.091779e-09, 1.093402e-09, 
    1.092259e-09, 1.097344e-09, 1.098869e-09, 1.106002e-09, 1.103075e-09, 
    1.107734e-09, 1.103548e-09, 1.10429e-09, 1.107886e-09, 1.103774e-09, 
    1.112768e-09, 1.10667e-09, 1.117996e-09, 1.111907e-09, 1.118377e-09, 
    1.117202e-09, 1.119147e-09, 1.12089e-09, 1.123082e-09, 1.127126e-09, 
    1.126189e-09, 1.129571e-09, 1.095024e-09, 1.097096e-09, 1.096914e-09, 
    1.099082e-09, 1.100686e-09, 1.104161e-09, 1.109736e-09, 1.10764e-09, 
    1.111488e-09, 1.112261e-09, 1.106414e-09, 1.110004e-09, 1.098483e-09, 
    1.100344e-09, 1.099236e-09, 1.095187e-09, 1.108123e-09, 1.101484e-09, 
    1.113742e-09, 1.110146e-09, 1.120641e-09, 1.115422e-09, 1.125674e-09, 
    1.130056e-09, 1.134181e-09, 1.139001e-09, 1.098227e-09, 1.096819e-09, 
    1.09934e-09, 1.102828e-09, 1.106063e-09, 1.110366e-09, 1.110806e-09, 
    1.111612e-09, 1.113699e-09, 1.115454e-09, 1.111867e-09, 1.115894e-09, 
    1.100776e-09, 1.108699e-09, 1.096287e-09, 1.100024e-09, 1.102622e-09, 
    1.101482e-09, 1.1074e-09, 1.108795e-09, 1.114462e-09, 1.111532e-09, 
    1.128975e-09, 1.121258e-09, 1.142671e-09, 1.136687e-09, 1.096327e-09, 
    1.098222e-09, 1.104817e-09, 1.101679e-09, 1.110653e-09, 1.112862e-09, 
    1.114657e-09, 1.116953e-09, 1.1172e-09, 1.11856e-09, 1.116332e-09, 
    1.118472e-09, 1.110375e-09, 1.113993e-09, 1.104063e-09, 1.10648e-09, 
    1.105368e-09, 1.104148e-09, 1.107913e-09, 1.111923e-09, 1.112009e-09, 
    1.113295e-09, 1.116919e-09, 1.110689e-09, 1.129971e-09, 1.118063e-09, 
    1.100288e-09, 1.103938e-09, 1.10446e-09, 1.103046e-09, 1.11264e-09, 
    1.109164e-09, 1.118527e-09, 1.115997e-09, 1.120143e-09, 1.118082e-09, 
    1.117779e-09, 1.115133e-09, 1.113486e-09, 1.109323e-09, 1.105936e-09, 
    1.103251e-09, 1.103875e-09, 1.106825e-09, 1.112168e-09, 1.117223e-09, 
    1.116116e-09, 1.119828e-09, 1.110002e-09, 1.114122e-09, 1.11253e-09, 
    1.116682e-09, 1.107584e-09, 1.115332e-09, 1.105603e-09, 1.106456e-09, 
    1.109095e-09, 1.114402e-09, 1.115576e-09, 1.116829e-09, 1.116056e-09, 
    1.112304e-09, 1.111689e-09, 1.109031e-09, 1.108297e-09, 1.106271e-09, 
    1.104593e-09, 1.106126e-09, 1.107735e-09, 1.112305e-09, 1.116424e-09, 
    1.120915e-09, 1.122013e-09, 1.12726e-09, 1.122989e-09, 1.130038e-09, 
    1.124046e-09, 1.134418e-09, 1.115781e-09, 1.123869e-09, 1.109215e-09, 
    1.110793e-09, 1.113649e-09, 1.120198e-09, 1.116662e-09, 1.120797e-09, 
    1.111665e-09, 1.106927e-09, 1.105701e-09, 1.103414e-09, 1.105753e-09, 
    1.105563e-09, 1.107802e-09, 1.107082e-09, 1.112457e-09, 1.10957e-09, 
    1.117772e-09, 1.120765e-09, 1.129217e-09, 1.134398e-09, 1.139673e-09, 
    1.142001e-09, 1.14271e-09, 1.143006e-09 ;

 SOIL2C_TO_SOIL3C =
  7.757447e-11, 7.791587e-11, 7.78495e-11, 7.812487e-11, 7.797211e-11, 
    7.815242e-11, 7.764368e-11, 7.792943e-11, 7.774701e-11, 7.76052e-11, 
    7.865926e-11, 7.813715e-11, 7.920156e-11, 7.886858e-11, 7.970501e-11, 
    7.914974e-11, 7.981697e-11, 7.968898e-11, 8.007417e-11, 7.996382e-11, 
    8.045652e-11, 8.01251e-11, 8.071191e-11, 8.037736e-11, 8.04297e-11, 
    8.011417e-11, 7.824221e-11, 7.859426e-11, 7.822135e-11, 7.827156e-11, 
    7.824903e-11, 7.797527e-11, 7.783731e-11, 7.754837e-11, 7.760082e-11, 
    7.781304e-11, 7.829413e-11, 7.813081e-11, 7.854239e-11, 7.853309e-11, 
    7.899129e-11, 7.87847e-11, 7.955481e-11, 7.933593e-11, 7.996842e-11, 
    7.980936e-11, 7.996095e-11, 7.991498e-11, 7.996155e-11, 7.972827e-11, 
    7.982822e-11, 7.962294e-11, 7.882339e-11, 7.905838e-11, 7.835754e-11, 
    7.793614e-11, 7.765621e-11, 7.745758e-11, 7.748566e-11, 7.75392e-11, 
    7.781428e-11, 7.807292e-11, 7.827001e-11, 7.840185e-11, 7.853176e-11, 
    7.892498e-11, 7.91331e-11, 7.959908e-11, 7.951497e-11, 7.965744e-11, 
    7.979353e-11, 8.002204e-11, 7.998443e-11, 8.00851e-11, 7.965367e-11, 
    7.99404e-11, 7.946707e-11, 7.959653e-11, 7.85671e-11, 7.817488e-11, 
    7.800818e-11, 7.786226e-11, 7.750726e-11, 7.775242e-11, 7.765577e-11, 
    7.788568e-11, 7.803178e-11, 7.795952e-11, 7.840546e-11, 7.823209e-11, 
    7.914543e-11, 7.875203e-11, 7.977766e-11, 7.953223e-11, 7.983648e-11, 
    7.968123e-11, 7.994726e-11, 7.970784e-11, 8.012256e-11, 8.021287e-11, 
    8.015116e-11, 8.038822e-11, 7.969456e-11, 7.996095e-11, 7.795749e-11, 
    7.796928e-11, 7.802418e-11, 7.778286e-11, 7.776809e-11, 7.754693e-11, 
    7.774372e-11, 7.782752e-11, 7.804024e-11, 7.816608e-11, 7.828569e-11, 
    7.854867e-11, 7.884239e-11, 7.92531e-11, 7.954814e-11, 7.974593e-11, 
    7.962465e-11, 7.973171e-11, 7.961203e-11, 7.955592e-11, 8.017904e-11, 
    7.982915e-11, 8.035412e-11, 8.032507e-11, 8.008749e-11, 8.032834e-11, 
    7.797755e-11, 7.790974e-11, 7.76743e-11, 7.785855e-11, 7.752285e-11, 
    7.771076e-11, 7.781881e-11, 7.823572e-11, 7.832731e-11, 7.841225e-11, 
    7.858e-11, 7.879528e-11, 7.917293e-11, 7.95015e-11, 7.980145e-11, 
    7.977947e-11, 7.978721e-11, 7.985422e-11, 7.968824e-11, 7.988147e-11, 
    7.99139e-11, 7.982911e-11, 8.032118e-11, 8.01806e-11, 8.032445e-11, 
    8.023292e-11, 7.793179e-11, 7.804589e-11, 7.798423e-11, 7.810018e-11, 
    7.801849e-11, 7.838172e-11, 7.849062e-11, 7.900017e-11, 7.879104e-11, 
    7.912386e-11, 7.882484e-11, 7.887783e-11, 7.913473e-11, 7.8841e-11, 
    7.94834e-11, 7.904789e-11, 7.985683e-11, 7.942194e-11, 7.988408e-11, 
    7.980015e-11, 7.99391e-11, 8.006355e-11, 8.022011e-11, 8.050898e-11, 
    8.044209e-11, 8.068367e-11, 7.8216e-11, 7.8364e-11, 7.835096e-11, 
    7.850585e-11, 7.862039e-11, 7.886866e-11, 7.926684e-11, 7.911711e-11, 
    7.939199e-11, 7.944718e-11, 7.902956e-11, 7.928598e-11, 7.846305e-11, 
    7.859602e-11, 7.851685e-11, 7.822767e-11, 7.915162e-11, 7.867746e-11, 
    7.955302e-11, 7.929615e-11, 8.004581e-11, 7.9673e-11, 8.040527e-11, 
    8.071832e-11, 8.101292e-11, 8.135723e-11, 7.844477e-11, 7.834421e-11, 
    7.852427e-11, 7.87734e-11, 7.900453e-11, 7.931183e-11, 7.934326e-11, 
    7.940083e-11, 7.954994e-11, 7.967531e-11, 7.941904e-11, 7.970674e-11, 
    7.862686e-11, 7.919278e-11, 7.830619e-11, 7.857318e-11, 7.875871e-11, 
    7.867731e-11, 7.909999e-11, 7.919961e-11, 7.960444e-11, 7.939516e-11, 
    8.064106e-11, 8.008984e-11, 8.161938e-11, 8.119194e-11, 7.830907e-11, 
    7.844442e-11, 7.89155e-11, 7.869136e-11, 7.933233e-11, 7.949011e-11, 
    7.961836e-11, 7.978232e-11, 7.980002e-11, 7.989717e-11, 7.973797e-11, 
    7.989087e-11, 7.931248e-11, 7.957095e-11, 7.886165e-11, 7.903429e-11, 
    7.895486e-11, 7.886775e-11, 7.913662e-11, 7.942308e-11, 7.942919e-11, 
    7.952104e-11, 7.97799e-11, 7.933493e-11, 8.071223e-11, 7.986166e-11, 
    7.859201e-11, 7.885274e-11, 7.888996e-11, 7.878897e-11, 7.94743e-11, 
    7.922598e-11, 7.989479e-11, 7.971403e-11, 8.00102e-11, 7.986303e-11, 
    7.984138e-11, 7.965235e-11, 7.953468e-11, 7.923737e-11, 7.899546e-11, 
    7.880362e-11, 7.884823e-11, 7.905895e-11, 7.944059e-11, 7.980162e-11, 
    7.972254e-11, 7.998769e-11, 7.928586e-11, 7.958015e-11, 7.946641e-11, 
    7.976299e-11, 7.911313e-11, 7.966656e-11, 7.897168e-11, 7.90326e-11, 
    7.922105e-11, 7.960013e-11, 7.968397e-11, 7.977353e-11, 7.971827e-11, 
    7.945028e-11, 7.940637e-11, 7.921647e-11, 7.916404e-11, 7.901933e-11, 
    7.889953e-11, 7.900899e-11, 7.912394e-11, 7.945039e-11, 7.974458e-11, 
    8.006532e-11, 8.014382e-11, 8.051859e-11, 8.021352e-11, 8.071696e-11, 
    8.028896e-11, 8.102984e-11, 7.969861e-11, 8.027636e-11, 7.922962e-11, 
    7.934239e-11, 7.954636e-11, 8.001416e-11, 7.97616e-11, 8.005696e-11, 
    7.940465e-11, 7.906623e-11, 7.897865e-11, 7.881528e-11, 7.898239e-11, 
    7.89688e-11, 7.91287e-11, 7.907731e-11, 7.946123e-11, 7.925501e-11, 
    7.984084e-11, 8.005462e-11, 8.065835e-11, 8.102846e-11, 8.14052e-11, 
    8.157151e-11, 8.162214e-11, 8.16433e-11 ;

 SOIL2C_vr =
  20.00646, 20.00647, 20.00647, 20.00648, 20.00648, 20.00648, 20.00646, 
    20.00647, 20.00646, 20.00646, 20.00651, 20.00648, 20.00654, 20.00652, 
    20.00656, 20.00653, 20.00657, 20.00656, 20.00658, 20.00657, 20.0066, 
    20.00658, 20.00661, 20.00659, 20.0066, 20.00658, 20.00649, 20.00651, 
    20.00649, 20.00649, 20.00649, 20.00648, 20.00647, 20.00645, 20.00646, 
    20.00647, 20.00649, 20.00648, 20.0065, 20.0065, 20.00653, 20.00652, 
    20.00655, 20.00654, 20.00657, 20.00657, 20.00657, 20.00657, 20.00657, 
    20.00656, 20.00657, 20.00656, 20.00652, 20.00653, 20.00649, 20.00647, 
    20.00646, 20.00645, 20.00645, 20.00645, 20.00647, 20.00648, 20.00649, 
    20.0065, 20.0065, 20.00652, 20.00653, 20.00656, 20.00655, 20.00656, 
    20.00657, 20.00658, 20.00657, 20.00658, 20.00656, 20.00657, 20.00655, 
    20.00656, 20.00651, 20.00648, 20.00648, 20.00647, 20.00645, 20.00646, 
    20.00646, 20.00647, 20.00648, 20.00648, 20.0065, 20.00649, 20.00653, 
    20.00651, 20.00657, 20.00655, 20.00657, 20.00656, 20.00657, 20.00656, 
    20.00658, 20.00659, 20.00658, 20.0066, 20.00656, 20.00657, 20.00648, 
    20.00648, 20.00648, 20.00647, 20.00647, 20.00645, 20.00646, 20.00647, 
    20.00648, 20.00648, 20.00649, 20.0065, 20.00652, 20.00654, 20.00655, 
    20.00656, 20.00656, 20.00656, 20.00656, 20.00655, 20.00658, 20.00657, 
    20.00659, 20.00659, 20.00658, 20.00659, 20.00648, 20.00647, 20.00646, 
    20.00647, 20.00645, 20.00646, 20.00647, 20.00649, 20.00649, 20.0065, 
    20.00651, 20.00652, 20.00653, 20.00655, 20.00657, 20.00657, 20.00657, 
    20.00657, 20.00656, 20.00657, 20.00657, 20.00657, 20.00659, 20.00658, 
    20.00659, 20.00659, 20.00647, 20.00648, 20.00648, 20.00648, 20.00648, 
    20.0065, 20.0065, 20.00653, 20.00652, 20.00653, 20.00652, 20.00652, 
    20.00653, 20.00652, 20.00655, 20.00653, 20.00657, 20.00655, 20.00657, 
    20.00657, 20.00657, 20.00658, 20.00659, 20.0066, 20.0066, 20.00661, 
    20.00649, 20.00649, 20.00649, 20.0065, 20.00651, 20.00652, 20.00654, 
    20.00653, 20.00655, 20.00655, 20.00653, 20.00654, 20.0065, 20.00651, 
    20.0065, 20.00649, 20.00653, 20.00651, 20.00655, 20.00654, 20.00658, 
    20.00656, 20.0066, 20.00661, 20.00663, 20.00664, 20.0065, 20.00649, 
    20.0065, 20.00652, 20.00653, 20.00654, 20.00654, 20.00655, 20.00655, 
    20.00656, 20.00655, 20.00656, 20.00651, 20.00654, 20.00649, 20.00651, 
    20.00652, 20.00651, 20.00653, 20.00654, 20.00656, 20.00655, 20.00661, 
    20.00658, 20.00665, 20.00663, 20.00649, 20.0065, 20.00652, 20.00651, 
    20.00654, 20.00655, 20.00656, 20.00657, 20.00657, 20.00657, 20.00656, 
    20.00657, 20.00654, 20.00656, 20.00652, 20.00653, 20.00653, 20.00652, 
    20.00653, 20.00655, 20.00655, 20.00655, 20.00657, 20.00654, 20.00661, 
    20.00657, 20.00651, 20.00652, 20.00652, 20.00652, 20.00655, 20.00654, 
    20.00657, 20.00656, 20.00658, 20.00657, 20.00657, 20.00656, 20.00655, 
    20.00654, 20.00653, 20.00652, 20.00652, 20.00653, 20.00655, 20.00657, 
    20.00656, 20.00657, 20.00654, 20.00656, 20.00655, 20.00656, 20.00653, 
    20.00656, 20.00653, 20.00653, 20.00654, 20.00656, 20.00656, 20.00657, 
    20.00656, 20.00655, 20.00655, 20.00654, 20.00653, 20.00653, 20.00652, 
    20.00653, 20.00653, 20.00655, 20.00656, 20.00658, 20.00658, 20.0066, 
    20.00659, 20.00661, 20.00659, 20.00663, 20.00656, 20.00659, 20.00654, 
    20.00654, 20.00655, 20.00658, 20.00656, 20.00658, 20.00655, 20.00653, 
    20.00653, 20.00652, 20.00653, 20.00653, 20.00653, 20.00653, 20.00655, 
    20.00654, 20.00657, 20.00658, 20.00661, 20.00663, 20.00665, 20.00665, 
    20.00665, 20.00666,
  20.00607, 20.00609, 20.00609, 20.00611, 20.0061, 20.00611, 20.00607, 
    20.00609, 20.00608, 20.00607, 20.00614, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00617, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00625, 20.00626, 20.00624, 20.00611, 20.00614, 
    20.00611, 20.00611, 20.00611, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00608, 20.00612, 20.00611, 20.00613, 20.00613, 20.00616, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00622, 20.00623, 
    20.00621, 20.00622, 20.0062, 20.00615, 20.00617, 20.00612, 20.00609, 
    20.00607, 20.00606, 20.00606, 20.00607, 20.00608, 20.0061, 20.00611, 
    20.00612, 20.00613, 20.00616, 20.00617, 20.0062, 20.0062, 20.00621, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.0062, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00607, 20.00609, 20.0061, 20.00609, 20.00612, 20.00611, 20.00617, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00624, 20.00624, 20.00626, 20.00621, 20.00623, 20.00609, 
    20.0061, 20.0061, 20.00608, 20.00608, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00613, 20.00615, 20.00618, 20.0062, 
    20.00621, 20.0062, 20.00621, 20.0062, 20.0062, 20.00624, 20.00622, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00607, 
    20.00609, 20.00607, 20.00608, 20.00608, 20.00611, 20.00612, 20.00612, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00622, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00624, 20.00609, 20.0061, 20.0061, 20.0061, 20.0061, 
    20.00612, 20.00613, 20.00616, 20.00615, 20.00617, 20.00615, 20.00616, 
    20.00617, 20.00615, 20.0062, 20.00617, 20.00622, 20.00619, 20.00622, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00626, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00618, 
    20.00617, 20.00619, 20.00619, 20.00617, 20.00618, 20.00613, 20.00614, 
    20.00613, 20.00611, 20.00617, 20.00614, 20.0062, 20.00618, 20.00623, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00613, 20.00615, 20.00616, 20.00618, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.00619, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00614, 20.00617, 20.00618, 20.0062, 20.00619, 20.00627, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00614, 
    20.00619, 20.0062, 20.0062, 20.00622, 20.00622, 20.00622, 20.00621, 
    20.00622, 20.00618, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00617, 20.00619, 20.00619, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00615, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00622, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00616, 20.00615, 20.00615, 20.00617, 20.00619, 20.00622, 
    20.00621, 20.00623, 20.00618, 20.0062, 20.0062, 20.00621, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.0062, 20.00621, 20.00621, 
    20.00621, 20.00619, 20.00619, 20.00618, 20.00617, 20.00616, 20.00616, 
    20.00616, 20.00617, 20.00619, 20.00621, 20.00623, 20.00624, 20.00626, 
    20.00624, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00623, 20.00621, 20.00623, 20.00619, 20.00617, 
    20.00616, 20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00623, 20.00627, 20.0063, 20.00632, 20.00633, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00552, 
    20.00554, 20.00553, 20.00552, 20.0056, 20.00556, 20.00563, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00572, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00564, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00566, 20.00561, 20.00562, 20.00558, 20.00554, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00555, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.00569, 20.00569, 20.0057, 20.00567, 20.00569, 20.00565, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00551, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00567, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00553, 20.00553, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00566, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00571, 20.0057, 20.00571, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00557, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00571, 20.0057, 
    20.00571, 20.00571, 20.00554, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00558, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00558, 20.00559, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.00569, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00557, 
    20.00559, 20.0056, 20.00562, 20.00564, 20.00564, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.00559, 20.00563, 20.00557, 20.00559, 
    20.0056, 20.0056, 20.00563, 20.00563, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.0058, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00564, 20.00566, 20.00566, 20.00568, 20.00568, 20.00568, 20.00567, 
    20.00568, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00564, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00561, 20.00561, 20.00565, 20.00564, 
    20.00568, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00562, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00565, 20.00567, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00567, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00561, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00576, 20.00567, 20.00571, 20.00564, 
    20.00564, 20.00566, 20.00569, 20.00567, 20.0057, 20.00565, 20.00562, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00565, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00576, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.0051, 20.0051, 20.00512, 20.00511, 20.00512, 20.00508, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.00519, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00525, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.0052, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00518, 20.00513, 20.00511, 
    20.00508, 20.00507, 20.00507, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00517, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00508, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.00509, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00521, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00514, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00525, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00513, 20.00515, 20.00515, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00515, 20.00519, 20.00513, 20.00515, 
    20.00516, 20.00516, 20.00519, 20.00519, 20.00522, 20.00521, 20.00529, 
    20.00526, 20.00536, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.0052, 20.00521, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.0052, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00518, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00523, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00523, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00525, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00523, 20.00525, 20.00521, 20.00518, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00536, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00446, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00438, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.00439, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00445, 20.00448, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00442, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00445, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00444, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258258, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.5258269, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258233, 0.5258234, 
    0.5258234, 0.5258229, 0.5258226, 0.5258222, 0.5258223, 0.5258226, 
    0.5258234, 0.5258232, 0.5258238, 0.5258238, 0.5258246, 0.5258242, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258262, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258243, 0.5258247, 
    0.5258235, 0.5258228, 0.5258223, 0.525822, 0.525822, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258236, 0.5258238, 0.5258245, 
    0.5258248, 0.5258256, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.5258229, 0.5258227, 0.5258221, 0.5258225, 
    0.5258223, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258248, 0.5258242, 0.5258259, 0.5258255, 0.525826, 0.5258258, 
    0.5258262, 0.5258258, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258262, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258225, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.525825, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.5258239, 0.5258243, 0.5258249, 0.5258254, 
    0.525826, 0.5258259, 0.525826, 0.525826, 0.5258258, 0.5258261, 0.5258262, 
    0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 0.5258228, 
    0.525823, 0.5258229, 0.5258231, 0.525823, 0.5258236, 0.5258238, 
    0.5258246, 0.5258242, 0.5258248, 0.5258243, 0.5258244, 0.5258248, 
    0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258253, 0.5258261, 
    0.525826, 0.5258262, 0.5258264, 0.5258267, 0.5258272, 0.5258271, 
    0.5258275, 0.5258233, 0.5258235, 0.5258235, 0.5258238, 0.525824, 
    0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 0.5258247, 
    0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258233, 0.5258249, 
    0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258257, 0.525827, 
    0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 0.5258238, 
    0.5258242, 0.5258246, 0.5258251, 0.5258252, 0.5258253, 0.5258256, 
    0.5258257, 0.5258253, 0.5258258, 0.525824, 0.525825, 0.5258235, 
    0.5258239, 0.5258242, 0.5258241, 0.5258248, 0.525825, 0.5258256, 
    0.5258253, 0.5258274, 0.5258265, 0.525829, 0.5258283, 0.5258235, 
    0.5258237, 0.5258245, 0.5258241, 0.5258252, 0.5258254, 0.5258257, 
    0.5258259, 0.525826, 0.5258262, 0.5258259, 0.5258262, 0.5258251, 
    0.5258256, 0.5258244, 0.5258247, 0.5258245, 0.5258244, 0.5258248, 
    0.5258253, 0.5258253, 0.5258255, 0.5258259, 0.5258252, 0.5258275, 
    0.5258261, 0.525824, 0.5258244, 0.5258244, 0.5258242, 0.5258254, 
    0.525825, 0.5258262, 0.5258259, 0.5258263, 0.5258261, 0.525826, 
    0.5258257, 0.5258255, 0.525825, 0.5258246, 0.5258243, 0.5258244, 
    0.5258247, 0.5258254, 0.525826, 0.5258259, 0.5258263, 0.5258251, 
    0.5258256, 0.5258254, 0.5258259, 0.5258248, 0.5258257, 0.5258246, 
    0.5258247, 0.525825, 0.5258256, 0.5258258, 0.5258259, 0.5258259, 
    0.5258254, 0.5258253, 0.525825, 0.5258249, 0.5258247, 0.5258244, 
    0.5258247, 0.5258248, 0.5258254, 0.5258259, 0.5258264, 0.5258266, 
    0.5258272, 0.5258267, 0.5258275, 0.5258268, 0.5258281, 0.5258258, 
    0.5258268, 0.525825, 0.5258252, 0.5258256, 0.5258263, 0.5258259, 
    0.5258264, 0.5258253, 0.5258247, 0.5258246, 0.5258243, 0.5258246, 
    0.5258245, 0.5258248, 0.5258248, 0.5258254, 0.5258251, 0.525826, 
    0.5258264, 0.5258274, 0.5258281, 0.5258287, 0.525829, 0.525829, 0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -1.28498e-20, -2.569961e-21, -1.027984e-20, -2.569961e-21, 1.28498e-20, 
    1.027984e-20, -1.027984e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    0, -1.28498e-20, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    2.055969e-20, 1.027984e-20, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -1.003089e-36, 7.709882e-21, 1.541976e-20, -1.28498e-20, 
    1.28498e-20, -1.28498e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, -1.003089e-36, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 1.798972e-20, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 1.798972e-20, -1.003089e-36, -1.027984e-20, -5.139921e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 1.798972e-20, 
    -5.139921e-21, 1.003089e-36, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 0, -5.139921e-21, 0, -1.027984e-20, -2.569961e-21, 
    -1.798972e-20, 2.312965e-20, 1.28498e-20, 2.569961e-21, -1.027984e-20, 
    1.28498e-20, 2.569961e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -7.709882e-21, -5.139921e-21, -1.28498e-20, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, -1.28498e-20, -7.709882e-21, 1.28498e-20, 1.28498e-20, 
    -1.027984e-20, 0, 5.139921e-21, -7.709882e-21, 1.027984e-20, 
    1.027984e-20, 1.541976e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 0, 2.569961e-21, -1.28498e-20, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, -1.28498e-20, 1.541976e-20, 1.798972e-20, 
    1.28498e-20, -1.003089e-36, 1.28498e-20, 1.798972e-20, -2.312965e-20, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, -2.055969e-20, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.798972e-20, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 0, 5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    0, 5.139921e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 0, -2.569961e-21, 1.798972e-20, -5.139921e-21, 
    1.798972e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, -1.798972e-20, 5.139921e-21, 
    1.28498e-20, -3.083953e-20, 1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -5.139921e-21, 1.003089e-36, 1.28498e-20, -5.139921e-21, 1.798972e-20, 
    2.569961e-21, 2.312965e-20, -1.798972e-20, -2.569961e-21, 1.027984e-20, 
    1.28498e-20, 1.027984e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -1.003089e-36, 2.312965e-20, 5.139921e-21, 7.709882e-21, -2.569961e-20, 
    -7.709882e-21, -5.139921e-21, 0, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, 0, 
    1.027984e-20, -7.709882e-21, 1.541976e-20, 5.139921e-21, -2.569961e-21, 
    -1.541976e-20, -5.139921e-21, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 1.541976e-20, 
    1.28498e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, 1.003089e-36, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, -1.003089e-36, 5.139921e-21, -1.28498e-20, 
    -1.541976e-20, 7.709882e-21, -1.027984e-20, 2.569961e-21, -1.027984e-20, 
    -1.003089e-36, 5.139921e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 1.798972e-20, -1.003089e-36, 5.139921e-21, -1.28498e-20, 
    1.027984e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    1.027984e-20, 1.28498e-20, -2.569961e-21, -5.139921e-21, 0, 
    -7.709882e-21, 0, 5.139921e-21, -1.541976e-20, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 1.28498e-20, 1.541976e-20, 1.28498e-20, 1.541976e-20, 
    -7.709882e-21, 2.055969e-20, 2.569961e-20, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    1.798972e-20, -1.541976e-20, 2.569961e-21, 1.027984e-20, 1.28498e-20, 
    -1.28498e-20, -1.798972e-20, -7.709882e-21, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -1.28498e-20, -2.569961e-21, 1.28498e-20, 
    1.798972e-20, 1.28498e-20, 5.139921e-21, 0, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 0, 1.541976e-20, 5.139921e-21, -1.798972e-20, 
    -1.28498e-20, 1.28498e-20, 0, -7.709882e-21, -1.027984e-20, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, 0, 2.569961e-21, -2.312965e-20, 
    -2.569961e-21, 1.798972e-20,
  1.027984e-20, 2.569961e-21, -1.003089e-36, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 0, -2.569961e-21, 2.569961e-21, 0, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, 1.798972e-20, 5.139921e-21, 
    -1.003089e-36, 5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 
    1.003089e-36, 5.139921e-21, 1.027984e-20, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, 1.027984e-20, 0, 0, -2.569961e-21, 0, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -1.003089e-36, 
    -2.569961e-21, -1.027984e-20, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 0, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    1.027984e-20, 0, 7.709882e-21, -1.027984e-20, 1.28498e-20, 7.709882e-21, 
    1.541976e-20, 0, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -2.569961e-20, 5.139921e-21, -2.569961e-21, -1.541976e-20, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.541976e-20, -7.709882e-21, 1.003089e-36, 
    -5.139921e-21, 2.569961e-21, 1.28498e-20, 7.709882e-21, -1.28498e-20, 0, 
    -5.139921e-21, -1.003089e-36, -7.709882e-21, -5.139921e-21, 1.003089e-36, 
    7.709882e-21, -7.709882e-21, -5.139921e-21, -1.28498e-20, 1.541976e-20, 
    -2.569961e-21, 0, -5.139921e-21, -5.139921e-21, -1.28498e-20, 
    1.798972e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, -1.027984e-20, -1.003089e-36, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, -1.541976e-20, 2.569961e-21, -2.569961e-21, 
    0, -5.139921e-21, 1.798972e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, 1.28498e-20, 0, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    0, -5.139921e-21, 5.139921e-21, 1.003089e-36, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, 0, 0, -7.709882e-21, 
    -5.139921e-21, 0, -2.569961e-21, -2.569961e-21, -5.139921e-21, 0, 
    -2.569961e-21, 2.569961e-21, 0, -2.569961e-21, 1.027984e-20, 
    1.541976e-20, -2.569961e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 0, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 0, 0, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 1.003089e-36, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 1.28498e-20, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, 1.28498e-20, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, -7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 0, 
    -7.709882e-21, -1.027984e-20, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    -7.709882e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 0, 1.027984e-20, 0, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, 0, -1.28498e-20, 
    2.569961e-21, 2.569961e-21, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    0, 2.569961e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, -2.569961e-21, -1.541976e-20, -5.139921e-21, 0, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 
    7.709882e-21, -5.139921e-21, -1.027984e-20, 0, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 0, 1.28498e-20, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -2.055969e-20, 7.709882e-21, -1.003089e-36, -7.709882e-21,
  1.027984e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 0, 1.027984e-20, 
    2.569961e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, 2.569961e-21, -2.569961e-21, -1.027984e-20, 0, 
    1.027984e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -1.798972e-20, -1.798972e-20, 7.709882e-21, -1.027984e-20, 
    -1.027984e-20, -1.798972e-20, 7.709882e-21, -2.569961e-21, 0, 
    1.541976e-20, 1.28498e-20, -1.003089e-36, 1.28498e-20, 7.709882e-21, 
    1.003089e-36, 1.003089e-36, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -2.569961e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -1.027984e-20, 1.28498e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 1.28498e-20, -2.569961e-21, 0, 
    -1.027984e-20, 1.541976e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    0, -1.003089e-36, -2.569961e-21, -1.28498e-20, 1.541976e-20, 
    7.709882e-21, -1.003089e-36, -1.28498e-20, -1.541976e-20, 0, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 0, 5.139921e-21, 1.28498e-20, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, 0, -1.541976e-20, -1.28498e-20, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, 1.28498e-20, -2.569961e-21, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 0, 
    -1.28498e-20, 2.569961e-21, 1.027984e-20, 1.003089e-36, -1.027984e-20, 
    -5.139921e-21, 0, -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.28498e-20, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, 
    0, -2.569961e-21, -1.28498e-20, 1.798972e-20, -2.569961e-21, 
    -1.798972e-20, -2.569961e-21, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    1.541976e-20, 2.569961e-21, 7.709882e-21, 1.28498e-20, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 1.28498e-20, 0, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, -1.003089e-36, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, 7.709882e-21, 
    1.28498e-20, 1.28498e-20, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -1.28498e-20, 0, 2.569961e-21, -1.28498e-20, -7.709882e-21, 
    -7.709882e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 0, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.003089e-36, 7.709882e-21, -5.139921e-21, -5.139921e-21, 1.798972e-20, 
    -1.28498e-20, 2.569961e-21, -7.709882e-21, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, -1.798972e-20, 
    -2.569961e-21, 2.569961e-21, -1.003089e-36, 7.709882e-21, 1.541976e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -2.569961e-21, -1.541976e-20, 
    -5.139921e-21, -1.003089e-36, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    0, -7.709882e-21, -5.139921e-21, -5.139921e-21, 0, -5.139921e-21, 
    1.28498e-20, 7.709882e-21, 2.569961e-21, 2.055969e-20, 1.027984e-20, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 0, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 
    2.569961e-21, 5.139921e-21, -1.027984e-20, 2.569961e-21, 1.003089e-36, 
    2.569961e-21, 0, 1.003089e-36, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    1.28498e-20, -1.28498e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, 0, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, -1.003089e-36, 
    0, 0, -2.569961e-21, -1.003089e-36, -5.139921e-21, 1.003089e-36, 0, 
    1.003089e-36, -1.027984e-20, 1.28498e-20, -5.139921e-21, -1.28498e-20, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, -1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -1.798972e-20, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, -1.003089e-36, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    0, 7.709882e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 1.003089e-36, 7.709882e-21, 0, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 0, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21,
  5.139921e-21, 1.541976e-20, 2.569961e-21, 0, 1.027984e-20, 1.541976e-20, 
    1.28498e-20, -7.709882e-21, -5.139921e-21, 1.003089e-36, 0, 
    -2.569961e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -1.027984e-20, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 1.027984e-20, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, 0, 0, 2.569961e-21, 5.139921e-21, 1.28498e-20, 0, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 2.055969e-20, 
    0, -2.055969e-20, -1.28498e-20, -2.569961e-21, -1.541976e-20, 0, 0, 
    -1.541976e-20, -1.28498e-20, 1.027984e-20, -1.798972e-20, -1.541976e-20, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 1.027984e-20, 
    1.28498e-20, 7.709882e-21, -7.709882e-21, -1.003089e-36, 1.003089e-36, 0, 
    1.541976e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, 1.28498e-20, 
    1.28498e-20, -5.139921e-21, 2.569961e-21, -1.798972e-20, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, -1.003089e-36, 2.569961e-21, 0, 
    0, 1.798972e-20, 0, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 0, 1.027984e-20, 0, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, -1.027984e-20, 0, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -1.28498e-20, 0, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -1.003089e-36, -1.027984e-20, -2.055969e-20, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, -2.055969e-20, 
    -5.139921e-21, -1.798972e-20, -1.027984e-20, 2.055969e-20, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, -2.055969e-20, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 1.003089e-36, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 0, 
    1.003089e-36, 5.139921e-21, -1.28498e-20, 1.003089e-36, -1.28498e-20, 
    2.569961e-21, 1.28498e-20, 1.28498e-20, -1.027984e-20, -7.709882e-21, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -1.003089e-36, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    2.055969e-20, 7.709882e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    0, -7.709882e-21, 3.083953e-20, -2.569961e-21, -1.027984e-20, 
    -7.709882e-21, -7.709882e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 0, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    1.28498e-20, 5.139921e-21, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 1.541976e-20, 
    7.709882e-21, 2.569961e-21, -1.541976e-20, 7.709882e-21, -1.28498e-20, 
    -2.569961e-21, 1.798972e-20, -7.709882e-21, 0, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 1.003089e-36, 
    -1.28498e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 0, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -2.055969e-20, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, 
    1.541976e-20, 1.28498e-20, 0, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    0, -2.569961e-21, 7.709882e-21, 0, 1.003089e-36, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 2.055969e-20, 2.569961e-21, 2.312965e-20, 5.139921e-21, 
    -2.569961e-21, -1.003089e-36, 1.027984e-20, -5.139921e-21, 1.798972e-20, 
    2.569961e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 1.027984e-20, 0, -1.027984e-20, -2.569961e-21, 
    1.541976e-20, -2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.28498e-20, 5.139921e-21, -1.027984e-20, 
    2.055969e-20, -2.569961e-21, 5.139921e-21, 1.541976e-20, -1.003089e-36, 
    2.055969e-20, -7.709882e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, -1.28498e-20, 7.709882e-21, 
    -1.027984e-20, -1.28498e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, 1.541976e-20, 1.003089e-36, 
    1.798972e-20, -2.569961e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, 
    1.28498e-20,
  2.569961e-21, 1.28498e-20, 2.569961e-21, -1.28498e-20, -2.569961e-21, 
    1.003089e-36, -1.003089e-36, 1.798972e-20, -5.139921e-21, -1.28498e-20, 
    -2.312965e-20, 2.569961e-21, 7.709882e-21, 1.541976e-20, -7.709882e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, -1.28498e-20, -1.027984e-20, 
    1.28498e-20, -1.027984e-20, 2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-20, 0, 
    -7.709882e-21, -7.709882e-21, 1.28498e-20, -1.541976e-20, 1.28498e-20, 
    2.569961e-21, 5.139921e-21, -1.541976e-20, 2.569961e-21, 1.798972e-20, 
    -5.139921e-21, -1.28498e-20, 1.798972e-20, -7.709882e-21, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, -2.569961e-21, 1.541976e-20, 1.003089e-36, 
    1.541976e-20, -2.569961e-21, -1.541976e-20, -7.709882e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 7.709882e-21, 1.541976e-20, 1.003089e-36, 
    2.055969e-20, 5.139921e-21, 2.312965e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, -1.541976e-20, 1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    0, 5.139921e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, -1.798972e-20, 3.083953e-20, 
    -2.569961e-20, -5.139921e-21, -1.541976e-20, -1.28498e-20, -1.28498e-20, 
    1.003089e-36, -1.027984e-20, -7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, -2.055969e-20, 1.798972e-20, -5.139921e-21, 2.055969e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, -1.798972e-20, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, -1.003089e-36, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-20, 2.569961e-21, -2.569961e-21, 
    -1.798972e-20, -5.139921e-21, 1.28498e-20, -2.569961e-21, 5.139921e-21, 
    0, -7.709882e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, -1.28498e-20, 1.541976e-20, -5.139921e-21, 
    -2.569961e-21, 1.28498e-20, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, 1.027984e-20, -1.798972e-20, 
    1.28498e-20, -7.709882e-21, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, 1.28498e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    7.709882e-21, 1.798972e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -1.541976e-20, -2.312965e-20, -5.139921e-21, -7.709882e-21, 
    -2.055969e-20, 7.709882e-21, 7.709882e-21, 1.003089e-36, -5.139921e-21, 
    2.569961e-21, -1.28498e-20, -2.569961e-21, 0, -1.28498e-20, 1.027984e-20, 
    -1.003089e-36, -1.798972e-20, 7.709882e-21, 2.569961e-21, 1.798972e-20, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, -1.541976e-20, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -2.312965e-20, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    1.798972e-20, -2.569961e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -2.569961e-21, 1.003089e-36, -1.28498e-20, -2.569961e-21, 1.798972e-20, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 2.055969e-20, 1.798972e-20, 
    -1.027984e-20, -1.28498e-20, -2.569961e-21, 0, -1.798972e-20, 
    1.541976e-20, 1.003089e-36, 1.28498e-20, -1.003089e-36, 7.709882e-21, 
    -5.139921e-21, 1.28498e-20, -1.798972e-20, 0, 7.709882e-21, 1.541976e-20, 
    5.015443e-37, -7.709882e-21, 2.569961e-21, -1.798972e-20, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, 0, 0, -2.569961e-20, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 1.28498e-20, -7.709882e-21, 
    -7.709882e-21, 7.709882e-21, -1.541976e-20, 0, -7.709882e-21, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 1.003089e-36, 7.709882e-21, 
    7.709882e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, -1.003089e-36, 
    1.798972e-20, 1.003089e-36, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -1.28498e-20, 1.798972e-20, -2.569961e-21, 2.569961e-21, 1.798972e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.541976e-20, 2.312965e-20, 
    -5.139921e-21, -7.709882e-21, 1.003089e-36, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, -1.28498e-20, 1.541976e-20, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, 2.055969e-20, 1.798972e-20, -1.28498e-20, 1.798972e-20, 
    -7.709882e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -1.541976e-20, -5.139921e-21, 
    7.709882e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, -1.541976e-20, 7.709882e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-20, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.541976e-20, 1.798972e-20, 2.569961e-21, 
    -1.541976e-20, 1.541976e-20,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259424e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.25942e-29, 6.259417e-29, 6.259414e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259453e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259466e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259426e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.25944e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259458e-29, 6.259458e-29, 6.259458e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259441e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259413e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.259459e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.259419e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259421e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259461e-29, 6.259463e-29, 
    6.259462e-29, 6.259467e-29, 6.259453e-29, 6.259458e-29, 6.259421e-29, 
    6.259422e-29, 6.259422e-29, 6.259418e-29, 6.259417e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259427e-29, 
    6.259432e-29, 6.259438e-29, 6.259445e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259454e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.259429e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259455e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259455e-29, 6.259458e-29, 6.259461e-29, 6.259463e-29, 6.259469e-29, 
    6.259467e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259429e-29, 
    6.259431e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259443e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.25943e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259432e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.25943e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259455e-29, 6.259457e-29, 6.259455e-29, 
    6.259457e-29, 6.259446e-29, 6.259451e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259456e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.259449e-29, 
    6.259445e-29, 6.259457e-29, 6.259454e-29, 6.259459e-29, 6.259456e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.25944e-29, 
    6.259437e-29, 6.259438e-29, 6.259441e-29, 6.259449e-29, 6.259455e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259444e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259444e-29, 6.259444e-29, 6.259441e-29, 
    6.259439e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259453e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.25946e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.25946e-29, 6.259472e-29, 6.259479e-29, 6.259485e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.194025e-10, 2.203681e-10, 2.201804e-10, 2.209592e-10, 2.205272e-10, 
    2.210371e-10, 2.195983e-10, 2.204065e-10, 2.198905e-10, 2.194894e-10, 
    2.224706e-10, 2.20994e-10, 2.240044e-10, 2.230627e-10, 2.254283e-10, 
    2.238579e-10, 2.25745e-10, 2.25383e-10, 2.264724e-10, 2.261603e-10, 
    2.275538e-10, 2.266164e-10, 2.282761e-10, 2.273299e-10, 2.27478e-10, 
    2.265855e-10, 2.212911e-10, 2.222868e-10, 2.212321e-10, 2.213741e-10, 
    2.213104e-10, 2.205361e-10, 2.201459e-10, 2.193287e-10, 2.194771e-10, 
    2.200773e-10, 2.21438e-10, 2.20976e-10, 2.221401e-10, 2.221138e-10, 
    2.234097e-10, 2.228254e-10, 2.250035e-10, 2.243845e-10, 2.261733e-10, 
    2.257234e-10, 2.261522e-10, 2.260222e-10, 2.261539e-10, 2.254941e-10, 
    2.257768e-10, 2.251962e-10, 2.229349e-10, 2.235995e-10, 2.216173e-10, 
    2.204254e-10, 2.196337e-10, 2.19072e-10, 2.191514e-10, 2.193028e-10, 
    2.200808e-10, 2.208123e-10, 2.213697e-10, 2.217426e-10, 2.2211e-10, 
    2.232222e-10, 2.238108e-10, 2.251287e-10, 2.248908e-10, 2.252938e-10, 
    2.256787e-10, 2.26325e-10, 2.262186e-10, 2.265033e-10, 2.252831e-10, 
    2.260941e-10, 2.247554e-10, 2.251215e-10, 2.2221e-10, 2.211007e-10, 
    2.206292e-10, 2.202165e-10, 2.192124e-10, 2.199058e-10, 2.196325e-10, 
    2.202827e-10, 2.206959e-10, 2.204916e-10, 2.217528e-10, 2.212625e-10, 
    2.238457e-10, 2.22733e-10, 2.256338e-10, 2.249397e-10, 2.258002e-10, 
    2.253611e-10, 2.261134e-10, 2.254363e-10, 2.266093e-10, 2.268647e-10, 
    2.266902e-10, 2.273606e-10, 2.253988e-10, 2.261522e-10, 2.204859e-10, 
    2.205192e-10, 2.206745e-10, 2.199919e-10, 2.199502e-10, 2.193247e-10, 
    2.198812e-10, 2.201182e-10, 2.207199e-10, 2.210758e-10, 2.214141e-10, 
    2.221579e-10, 2.229886e-10, 2.241502e-10, 2.249846e-10, 2.25544e-10, 
    2.25201e-10, 2.255038e-10, 2.251653e-10, 2.250067e-10, 2.26769e-10, 
    2.257794e-10, 2.272642e-10, 2.27182e-10, 2.265101e-10, 2.271913e-10, 
    2.205426e-10, 2.203508e-10, 2.196849e-10, 2.20206e-10, 2.192565e-10, 
    2.19788e-10, 2.200936e-10, 2.212728e-10, 2.215318e-10, 2.21772e-10, 
    2.222464e-10, 2.228553e-10, 2.239234e-10, 2.248527e-10, 2.257011e-10, 
    2.256389e-10, 2.256608e-10, 2.258503e-10, 2.253809e-10, 2.259274e-10, 
    2.260191e-10, 2.257793e-10, 2.27171e-10, 2.267734e-10, 2.271803e-10, 
    2.269214e-10, 2.204131e-10, 2.207359e-10, 2.205615e-10, 2.208894e-10, 
    2.206584e-10, 2.216857e-10, 2.219937e-10, 2.234348e-10, 2.228433e-10, 
    2.237846e-10, 2.229389e-10, 2.230888e-10, 2.238154e-10, 2.229846e-10, 
    2.248015e-10, 2.235698e-10, 2.258577e-10, 2.246277e-10, 2.259348e-10, 
    2.256974e-10, 2.260904e-10, 2.264424e-10, 2.268851e-10, 2.277022e-10, 
    2.27513e-10, 2.281962e-10, 2.21217e-10, 2.216356e-10, 2.215987e-10, 
    2.220368e-10, 2.223607e-10, 2.230629e-10, 2.241891e-10, 2.237656e-10, 
    2.24543e-10, 2.246991e-10, 2.235179e-10, 2.242432e-10, 2.219157e-10, 
    2.222918e-10, 2.220679e-10, 2.2125e-10, 2.238632e-10, 2.225221e-10, 
    2.249984e-10, 2.24272e-10, 2.263922e-10, 2.253378e-10, 2.274088e-10, 
    2.282942e-10, 2.291275e-10, 2.301013e-10, 2.21864e-10, 2.215796e-10, 
    2.220888e-10, 2.227935e-10, 2.234472e-10, 2.243163e-10, 2.244052e-10, 
    2.24568e-10, 2.249897e-10, 2.253443e-10, 2.246195e-10, 2.254332e-10, 
    2.22379e-10, 2.239796e-10, 2.214721e-10, 2.222272e-10, 2.227519e-10, 
    2.225217e-10, 2.237172e-10, 2.239989e-10, 2.251439e-10, 2.24552e-10, 
    2.280757e-10, 2.265167e-10, 2.308427e-10, 2.296338e-10, 2.214802e-10, 
    2.21863e-10, 2.231954e-10, 2.225614e-10, 2.243743e-10, 2.248205e-10, 
    2.251832e-10, 2.25647e-10, 2.25697e-10, 2.259718e-10, 2.255215e-10, 
    2.25954e-10, 2.243181e-10, 2.250491e-10, 2.23043e-10, 2.235313e-10, 
    2.233067e-10, 2.230603e-10, 2.238207e-10, 2.246309e-10, 2.246482e-10, 
    2.24908e-10, 2.256401e-10, 2.243816e-10, 2.28277e-10, 2.258714e-10, 
    2.222805e-10, 2.230178e-10, 2.231231e-10, 2.228375e-10, 2.247758e-10, 
    2.240735e-10, 2.259651e-10, 2.254538e-10, 2.262915e-10, 2.258752e-10, 
    2.25814e-10, 2.252794e-10, 2.249466e-10, 2.241057e-10, 2.234215e-10, 
    2.228789e-10, 2.230051e-10, 2.236011e-10, 2.246805e-10, 2.257016e-10, 
    2.254779e-10, 2.262278e-10, 2.242428e-10, 2.250752e-10, 2.247535e-10, 
    2.255923e-10, 2.237543e-10, 2.253196e-10, 2.233542e-10, 2.235265e-10, 
    2.240595e-10, 2.251317e-10, 2.253688e-10, 2.256221e-10, 2.254658e-10, 
    2.247079e-10, 2.245837e-10, 2.240466e-10, 2.238983e-10, 2.23489e-10, 
    2.231502e-10, 2.234598e-10, 2.237849e-10, 2.247082e-10, 2.255402e-10, 
    2.264474e-10, 2.266694e-10, 2.277293e-10, 2.268665e-10, 2.282904e-10, 
    2.270799e-10, 2.291753e-10, 2.254102e-10, 2.270442e-10, 2.240838e-10, 
    2.244027e-10, 2.249796e-10, 2.263027e-10, 2.255884e-10, 2.264237e-10, 
    2.245788e-10, 2.236216e-10, 2.23374e-10, 2.229119e-10, 2.233845e-10, 
    2.233461e-10, 2.237983e-10, 2.23653e-10, 2.247388e-10, 2.241556e-10, 
    2.258125e-10, 2.264171e-10, 2.281246e-10, 2.291714e-10, 2.302369e-10, 
    2.307073e-10, 2.308505e-10, 2.309103e-10 ;

 SOIL2N_TO_SOIL3N =
  1.567161e-11, 1.574058e-11, 1.572717e-11, 1.57828e-11, 1.575194e-11, 
    1.578837e-11, 1.568559e-11, 1.574332e-11, 1.570647e-11, 1.567782e-11, 
    1.589076e-11, 1.578528e-11, 1.600031e-11, 1.593305e-11, 1.610202e-11, 
    1.598985e-11, 1.612464e-11, 1.609878e-11, 1.61766e-11, 1.615431e-11, 
    1.625384e-11, 1.618689e-11, 1.630544e-11, 1.623785e-11, 1.624842e-11, 
    1.618468e-11, 1.580651e-11, 1.587763e-11, 1.580229e-11, 1.581244e-11, 
    1.580788e-11, 1.575258e-11, 1.572471e-11, 1.566634e-11, 1.567693e-11, 
    1.571981e-11, 1.5817e-11, 1.5784e-11, 1.586715e-11, 1.586527e-11, 
    1.595784e-11, 1.59161e-11, 1.607168e-11, 1.602746e-11, 1.615524e-11, 
    1.61231e-11, 1.615373e-11, 1.614444e-11, 1.615385e-11, 1.610672e-11, 
    1.612691e-11, 1.608544e-11, 1.592392e-11, 1.597139e-11, 1.582981e-11, 
    1.574467e-11, 1.568812e-11, 1.5648e-11, 1.565367e-11, 1.566448e-11, 
    1.572006e-11, 1.577231e-11, 1.581212e-11, 1.583876e-11, 1.5865e-11, 
    1.594444e-11, 1.598648e-11, 1.608062e-11, 1.606363e-11, 1.609241e-11, 
    1.611991e-11, 1.616607e-11, 1.615847e-11, 1.617881e-11, 1.609165e-11, 
    1.614958e-11, 1.605395e-11, 1.608011e-11, 1.587214e-11, 1.57929e-11, 
    1.575923e-11, 1.572975e-11, 1.565803e-11, 1.570756e-11, 1.568803e-11, 
    1.573448e-11, 1.5764e-11, 1.57494e-11, 1.583949e-11, 1.580446e-11, 
    1.598898e-11, 1.59095e-11, 1.61167e-11, 1.606712e-11, 1.612858e-11, 
    1.609722e-11, 1.615096e-11, 1.610259e-11, 1.618638e-11, 1.620462e-11, 
    1.619215e-11, 1.624004e-11, 1.609991e-11, 1.615373e-11, 1.574899e-11, 
    1.575137e-11, 1.576246e-11, 1.571371e-11, 1.571073e-11, 1.566605e-11, 
    1.57058e-11, 1.572273e-11, 1.576571e-11, 1.579113e-11, 1.581529e-11, 
    1.586842e-11, 1.592776e-11, 1.601073e-11, 1.607033e-11, 1.611029e-11, 
    1.608579e-11, 1.610742e-11, 1.608324e-11, 1.60719e-11, 1.619779e-11, 
    1.61271e-11, 1.623316e-11, 1.622729e-11, 1.617929e-11, 1.622795e-11, 
    1.575304e-11, 1.573934e-11, 1.569178e-11, 1.5729e-11, 1.566118e-11, 
    1.569914e-11, 1.572097e-11, 1.58052e-11, 1.58237e-11, 1.584086e-11, 
    1.587475e-11, 1.591824e-11, 1.599453e-11, 1.606091e-11, 1.612151e-11, 
    1.611707e-11, 1.611863e-11, 1.613217e-11, 1.609863e-11, 1.613767e-11, 
    1.614422e-11, 1.612709e-11, 1.62265e-11, 1.61981e-11, 1.622716e-11, 
    1.620867e-11, 1.57438e-11, 1.576685e-11, 1.575439e-11, 1.577781e-11, 
    1.576131e-11, 1.583469e-11, 1.585669e-11, 1.595963e-11, 1.591738e-11, 
    1.598462e-11, 1.592421e-11, 1.593491e-11, 1.598681e-11, 1.592747e-11, 
    1.605725e-11, 1.596927e-11, 1.613269e-11, 1.604484e-11, 1.61382e-11, 
    1.612124e-11, 1.614931e-11, 1.617445e-11, 1.620608e-11, 1.626444e-11, 
    1.625093e-11, 1.629973e-11, 1.580121e-11, 1.583111e-11, 1.582848e-11, 
    1.585977e-11, 1.588291e-11, 1.593306e-11, 1.60135e-11, 1.598325e-11, 
    1.603879e-11, 1.604994e-11, 1.596557e-11, 1.601737e-11, 1.585112e-11, 
    1.587798e-11, 1.586199e-11, 1.580357e-11, 1.599023e-11, 1.589444e-11, 
    1.607132e-11, 1.601943e-11, 1.617087e-11, 1.609556e-11, 1.624349e-11, 
    1.630673e-11, 1.636625e-11, 1.643581e-11, 1.584743e-11, 1.582711e-11, 
    1.586349e-11, 1.591382e-11, 1.596051e-11, 1.602259e-11, 1.602894e-11, 
    1.604057e-11, 1.60707e-11, 1.609602e-11, 1.604425e-11, 1.610237e-11, 
    1.588422e-11, 1.599854e-11, 1.581943e-11, 1.587337e-11, 1.591085e-11, 
    1.589441e-11, 1.59798e-11, 1.599992e-11, 1.608171e-11, 1.603943e-11, 
    1.629112e-11, 1.617977e-11, 1.648876e-11, 1.640241e-11, 1.582001e-11, 
    1.584736e-11, 1.594253e-11, 1.589725e-11, 1.602673e-11, 1.605861e-11, 
    1.608452e-11, 1.611764e-11, 1.612122e-11, 1.614084e-11, 1.610868e-11, 
    1.613957e-11, 1.602272e-11, 1.607494e-11, 1.593164e-11, 1.596652e-11, 
    1.595048e-11, 1.593288e-11, 1.59872e-11, 1.604507e-11, 1.60463e-11, 
    1.606486e-11, 1.611715e-11, 1.602726e-11, 1.63055e-11, 1.613367e-11, 
    1.587717e-11, 1.592985e-11, 1.593737e-11, 1.591696e-11, 1.605541e-11, 
    1.600525e-11, 1.614036e-11, 1.610385e-11, 1.616368e-11, 1.613394e-11, 
    1.612957e-11, 1.609139e-11, 1.606761e-11, 1.600755e-11, 1.595868e-11, 
    1.591992e-11, 1.592893e-11, 1.597151e-11, 1.604861e-11, 1.612154e-11, 
    1.610556e-11, 1.615913e-11, 1.601735e-11, 1.60768e-11, 1.605382e-11, 
    1.611374e-11, 1.598245e-11, 1.609425e-11, 1.595387e-11, 1.596618e-11, 
    1.600425e-11, 1.608083e-11, 1.609777e-11, 1.611586e-11, 1.61047e-11, 
    1.605056e-11, 1.604169e-11, 1.600333e-11, 1.599273e-11, 1.59635e-11, 
    1.59393e-11, 1.596141e-11, 1.598464e-11, 1.605058e-11, 1.611002e-11, 
    1.617481e-11, 1.619067e-11, 1.626638e-11, 1.620475e-11, 1.630646e-11, 
    1.621999e-11, 1.636967e-11, 1.610073e-11, 1.621745e-11, 1.600598e-11, 
    1.602877e-11, 1.606997e-11, 1.616448e-11, 1.611345e-11, 1.617312e-11, 
    1.604134e-11, 1.597297e-11, 1.595528e-11, 1.592228e-11, 1.595604e-11, 
    1.595329e-11, 1.598559e-11, 1.597521e-11, 1.605277e-11, 1.601111e-11, 
    1.612946e-11, 1.617265e-11, 1.629462e-11, 1.636939e-11, 1.644549e-11, 
    1.647909e-11, 1.648932e-11, 1.64936e-11 ;

 SOIL2N_vr =
  1.818769, 1.81877, 1.81877, 1.818771, 1.818771, 1.818771, 1.818769, 
    1.81877, 1.81877, 1.818769, 1.818774, 1.818771, 1.818776, 1.818775, 
    1.818778, 1.818776, 1.818779, 1.818778, 1.81878, 1.818779, 1.818782, 
    1.81878, 1.818783, 1.818781, 1.818781, 1.81878, 1.818772, 1.818773, 
    1.818772, 1.818772, 1.818772, 1.818771, 1.81877, 1.818769, 1.818769, 
    1.81877, 1.818772, 1.818771, 1.818773, 1.818773, 1.818775, 1.818774, 
    1.818778, 1.818777, 1.818779, 1.818779, 1.818779, 1.818779, 1.818779, 
    1.818778, 1.818779, 1.818778, 1.818774, 1.818775, 1.818772, 1.81877, 
    1.818769, 1.818768, 1.818768, 1.818769, 1.81877, 1.818771, 1.818772, 
    1.818772, 1.818773, 1.818775, 1.818776, 1.818778, 1.818777, 1.818778, 
    1.818779, 1.81878, 1.81878, 1.81878, 1.818778, 1.818779, 1.818777, 
    1.818778, 1.818773, 1.818771, 1.818771, 1.81877, 1.818768, 1.81877, 
    1.818769, 1.81877, 1.818771, 1.818771, 1.818772, 1.818772, 1.818776, 
    1.818774, 1.818779, 1.818778, 1.818779, 1.818778, 1.818779, 1.818778, 
    1.81878, 1.818781, 1.81878, 1.818781, 1.818778, 1.818779, 1.81877, 
    1.818771, 1.818771, 1.81877, 1.81877, 1.818769, 1.818769, 1.81877, 
    1.818771, 1.818771, 1.818772, 1.818773, 1.818774, 1.818776, 1.818778, 
    1.818779, 1.818778, 1.818778, 1.818778, 1.818778, 1.81878, 1.818779, 
    1.818781, 1.818781, 1.81878, 1.818781, 1.818771, 1.81877, 1.818769, 
    1.81877, 1.818769, 1.818769, 1.81877, 1.818772, 1.818772, 1.818773, 
    1.818773, 1.818774, 1.818776, 1.818777, 1.818779, 1.818779, 1.818779, 
    1.818779, 1.818778, 1.818779, 1.818779, 1.818779, 1.818781, 1.81878, 
    1.818781, 1.818781, 1.81877, 1.818771, 1.818771, 1.818771, 1.818771, 
    1.818772, 1.818773, 1.818775, 1.818774, 1.818776, 1.818774, 1.818775, 
    1.818776, 1.818774, 1.818777, 1.818775, 1.818779, 1.818777, 1.818779, 
    1.818779, 1.818779, 1.81878, 1.818781, 1.818782, 1.818782, 1.818783, 
    1.818772, 1.818772, 1.818772, 1.818773, 1.818773, 1.818775, 1.818776, 
    1.818776, 1.818777, 1.818777, 1.818775, 1.818776, 1.818773, 1.818773, 
    1.818773, 1.818772, 1.818776, 1.818774, 1.818778, 1.818776, 1.81878, 
    1.818778, 1.818781, 1.818783, 1.818784, 1.818786, 1.818773, 1.818772, 
    1.818773, 1.818774, 1.818775, 1.818776, 1.818777, 1.818777, 1.818778, 
    1.818778, 1.818777, 1.818778, 1.818774, 1.818776, 1.818772, 1.818773, 
    1.818774, 1.818774, 1.818776, 1.818776, 1.818778, 1.818777, 1.818782, 
    1.81878, 1.818787, 1.818785, 1.818772, 1.818773, 1.818775, 1.818774, 
    1.818777, 1.818777, 1.818778, 1.818779, 1.818779, 1.818779, 1.818778, 
    1.818779, 1.818776, 1.818778, 1.818774, 1.818775, 1.818775, 1.818775, 
    1.818776, 1.818777, 1.818777, 1.818777, 1.818779, 1.818777, 1.818783, 
    1.818779, 1.818773, 1.818774, 1.818775, 1.818774, 1.818777, 1.818776, 
    1.818779, 1.818778, 1.81878, 1.818779, 1.818779, 1.818778, 1.818778, 
    1.818776, 1.818775, 1.818774, 1.818774, 1.818775, 1.818777, 1.818779, 
    1.818778, 1.81878, 1.818776, 1.818778, 1.818777, 1.818779, 1.818776, 
    1.818778, 1.818775, 1.818775, 1.818776, 1.818778, 1.818778, 1.818779, 
    1.818778, 1.818777, 1.818777, 1.818776, 1.818776, 1.818775, 1.818775, 
    1.818775, 1.818776, 1.818777, 1.818779, 1.81878, 1.81878, 1.818782, 
    1.818781, 1.818783, 1.818781, 1.818784, 1.818778, 1.818781, 1.818776, 
    1.818777, 1.818778, 1.81878, 1.818779, 1.81878, 1.818777, 1.818775, 
    1.818775, 1.818774, 1.818775, 1.818775, 1.818776, 1.818776, 1.818777, 
    1.818776, 1.818779, 1.81878, 1.818783, 1.818784, 1.818786, 1.818787, 
    1.818787, 1.818787,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818743, 1.818741, 
    1.818746, 1.818743, 1.818747, 1.818746, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818752, 1.81875, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818733, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.818739, 1.818739, 1.818742, 1.818741, 
    1.818745, 1.818744, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818738, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818733, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.818739, 1.818742, 1.818743, 1.818746, 1.818745, 1.818746, 
    1.818747, 1.818748, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818737, 1.818736, 1.818735, 1.818733, 1.818735, 
    1.818734, 1.818735, 1.818736, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 
    1.818749, 1.818749, 1.818749, 1.818751, 1.818746, 1.818748, 1.818736, 
    1.818736, 1.818736, 1.818735, 1.818735, 1.818733, 1.818735, 1.818735, 
    1.818736, 1.818737, 1.818738, 1.818739, 1.818741, 1.818744, 1.818745, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818745, 1.818749, 1.818747, 
    1.81875, 1.81875, 1.818749, 1.81875, 1.818736, 1.818736, 1.818734, 
    1.818735, 1.818733, 1.818734, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818747, 1.818746, 1.818747, 1.818748, 1.818747, 1.81875, 1.818749, 
    1.81875, 1.81875, 1.818736, 1.818736, 1.818736, 1.818737, 1.818736, 
    1.818738, 1.818739, 1.818742, 1.818741, 1.818743, 1.818741, 1.818741, 
    1.818743, 1.818741, 1.818745, 1.818742, 1.818747, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.818749, 1.818751, 1.818751, 1.818752, 
    1.818737, 1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818742, 1.818744, 1.818739, 1.81874, 
    1.818739, 1.818738, 1.818743, 1.81874, 1.818745, 1.818744, 1.818748, 
    1.818746, 1.818751, 1.818753, 1.818754, 1.818756, 1.818739, 1.818738, 
    1.818739, 1.818741, 1.818742, 1.818744, 1.818744, 1.818745, 1.818745, 
    1.818746, 1.818745, 1.818746, 1.81874, 1.818743, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818743, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818755, 1.818738, 1.818739, 1.818742, 1.81874, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818741, 1.818742, 1.818742, 1.818741, 
    1.818743, 1.818745, 1.818745, 1.818745, 1.818747, 1.818744, 1.818752, 
    1.818747, 1.81874, 1.818741, 1.818741, 1.818741, 1.818745, 1.818743, 
    1.818748, 1.818746, 1.818748, 1.818747, 1.818747, 1.818746, 1.818745, 
    1.818744, 1.818742, 1.818741, 1.818741, 1.818743, 1.818745, 1.818747, 
    1.818746, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818742, 1.818743, 1.818746, 1.818746, 1.818747, 
    1.818746, 1.818745, 1.818745, 1.818743, 1.818743, 1.818742, 1.818742, 
    1.818742, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818751, 
    1.818749, 1.818752, 1.81875, 1.818754, 1.818746, 1.81875, 1.818744, 
    1.818744, 1.818745, 1.818748, 1.818747, 1.818748, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818747, 1.818748, 1.818752, 1.818754, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818685, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818683, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818697, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818683, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818687, 1.818686, 1.818685, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818686, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818686, 1.818685, 1.818685, 1.818683, 1.818685, 1.818685, 
    1.818687, 1.818687, 1.818688, 1.81869, 1.818692, 1.818694, 1.818696, 
    1.818698, 1.818697, 1.818697, 1.818697, 1.818696, 1.8187, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818701, 1.818686, 1.818686, 1.818684, 
    1.818685, 1.818683, 1.818684, 1.818685, 1.818688, 1.818688, 1.818689, 
    1.81869, 1.818691, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818698, 1.818699, 1.818698, 1.818701, 1.8187, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818686, 
    1.818689, 1.818689, 1.818693, 1.818691, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818695, 1.818698, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818702, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.81869, 1.818692, 1.818694, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.818699, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818695, 1.818696, 
    1.818697, 1.818695, 1.818697, 1.81869, 1.818694, 1.818688, 1.81869, 
    1.818691, 1.818691, 1.818693, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.818709, 1.818707, 1.818688, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818697, 
    1.818699, 1.818695, 1.818696, 1.818692, 1.818693, 1.818692, 1.818692, 
    1.818694, 1.818695, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818691, 1.818696, 1.818694, 
    1.818699, 1.818697, 1.818699, 1.818698, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818691, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818697, 1.818699, 1.818695, 1.818696, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818697, 1.818696, 1.818695, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818702, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818695, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818694, 1.818698, 1.818699, 1.818703, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818643, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818657, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818643, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818646, 1.818645, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.81866, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818643, 1.818645, 1.818645, 
    1.818647, 1.818647, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818657, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818645, 1.818643, 1.818645, 1.818645, 1.818648, 1.818648, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818646, 
    1.818649, 1.81865, 1.818653, 1.818651, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.81866, 1.818662, 1.818662, 1.818663, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818654, 
    1.818653, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.818659, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.818669, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818658, 1.818657, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818655, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818651, 1.818656, 1.818654, 
    1.818658, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818651, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818656, 1.818656, 1.818658, 1.818653, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818662, 
    1.81866, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818659, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818586, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.81859, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818587, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.818589, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.81859, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.327385e-09, 1.333227e-09, 1.332091e-09, 1.336803e-09, 1.334189e-09, 
    1.337275e-09, 1.32857e-09, 1.333459e-09, 1.330338e-09, 1.327911e-09, 
    1.345947e-09, 1.337013e-09, 1.355227e-09, 1.349529e-09, 1.363841e-09, 
    1.35434e-09, 1.365757e-09, 1.363567e-09, 1.370158e-09, 1.36827e-09, 
    1.3767e-09, 1.37103e-09, 1.38107e-09, 1.375346e-09, 1.376242e-09, 
    1.370842e-09, 1.338811e-09, 1.344835e-09, 1.338454e-09, 1.339313e-09, 
    1.338928e-09, 1.334243e-09, 1.331883e-09, 1.326939e-09, 1.327836e-09, 
    1.331468e-09, 1.3397e-09, 1.336905e-09, 1.343948e-09, 1.343789e-09, 
    1.351629e-09, 1.348094e-09, 1.361271e-09, 1.357526e-09, 1.368349e-09, 
    1.365627e-09, 1.368221e-09, 1.367434e-09, 1.368231e-09, 1.364239e-09, 
    1.365949e-09, 1.362437e-09, 1.348756e-09, 1.352777e-09, 1.340784e-09, 
    1.333574e-09, 1.328784e-09, 1.325385e-09, 1.325866e-09, 1.326782e-09, 
    1.331489e-09, 1.335914e-09, 1.339287e-09, 1.341543e-09, 1.343766e-09, 
    1.350494e-09, 1.354055e-09, 1.362029e-09, 1.36059e-09, 1.363027e-09, 
    1.365356e-09, 1.369266e-09, 1.368622e-09, 1.370345e-09, 1.362963e-09, 
    1.367869e-09, 1.35977e-09, 1.361985e-09, 1.344371e-09, 1.337659e-09, 
    1.334807e-09, 1.33231e-09, 1.326235e-09, 1.33043e-09, 1.328777e-09, 
    1.332711e-09, 1.33521e-09, 1.333974e-09, 1.341604e-09, 1.338638e-09, 
    1.354266e-09, 1.347535e-09, 1.365084e-09, 1.360885e-09, 1.366091e-09, 
    1.363434e-09, 1.367986e-09, 1.36389e-09, 1.370986e-09, 1.372531e-09, 
    1.371475e-09, 1.375532e-09, 1.363663e-09, 1.368221e-09, 1.333939e-09, 
    1.334141e-09, 1.33508e-09, 1.330951e-09, 1.330698e-09, 1.326914e-09, 
    1.330281e-09, 1.331715e-09, 1.335355e-09, 1.337508e-09, 1.339555e-09, 
    1.344055e-09, 1.349081e-09, 1.356108e-09, 1.361157e-09, 1.364541e-09, 
    1.362466e-09, 1.364298e-09, 1.36225e-09, 1.36129e-09, 1.371952e-09, 
    1.365965e-09, 1.374948e-09, 1.374451e-09, 1.370386e-09, 1.374507e-09, 
    1.334283e-09, 1.333122e-09, 1.329094e-09, 1.332246e-09, 1.326502e-09, 
    1.329718e-09, 1.331566e-09, 1.3387e-09, 1.340267e-09, 1.341721e-09, 
    1.344591e-09, 1.348275e-09, 1.354737e-09, 1.360359e-09, 1.365491e-09, 
    1.365115e-09, 1.365248e-09, 1.366394e-09, 1.363554e-09, 1.366861e-09, 
    1.367416e-09, 1.365965e-09, 1.374385e-09, 1.371979e-09, 1.374441e-09, 
    1.372874e-09, 1.333499e-09, 1.335452e-09, 1.334397e-09, 1.336381e-09, 
    1.334983e-09, 1.341198e-09, 1.343062e-09, 1.351781e-09, 1.348202e-09, 
    1.353897e-09, 1.348781e-09, 1.349687e-09, 1.354083e-09, 1.349057e-09, 
    1.360049e-09, 1.352597e-09, 1.366439e-09, 1.358998e-09, 1.366905e-09, 
    1.365469e-09, 1.367847e-09, 1.369976e-09, 1.372655e-09, 1.377598e-09, 
    1.376454e-09, 1.380587e-09, 1.338363e-09, 1.340895e-09, 1.340672e-09, 
    1.343322e-09, 1.345282e-09, 1.34953e-09, 1.356344e-09, 1.353782e-09, 
    1.358485e-09, 1.359429e-09, 1.352284e-09, 1.356671e-09, 1.34259e-09, 
    1.344865e-09, 1.34351e-09, 1.338562e-09, 1.354372e-09, 1.346259e-09, 
    1.361241e-09, 1.356845e-09, 1.369673e-09, 1.363293e-09, 1.375823e-09, 
    1.38118e-09, 1.386221e-09, 1.392113e-09, 1.342277e-09, 1.340556e-09, 
    1.343637e-09, 1.3479e-09, 1.351855e-09, 1.357113e-09, 1.357651e-09, 
    1.358636e-09, 1.361188e-09, 1.363333e-09, 1.358948e-09, 1.363871e-09, 
    1.345393e-09, 1.355076e-09, 1.339906e-09, 1.344474e-09, 1.347649e-09, 
    1.346256e-09, 1.353489e-09, 1.355193e-09, 1.36212e-09, 1.35854e-09, 
    1.379858e-09, 1.370426e-09, 1.396598e-09, 1.389284e-09, 1.339955e-09, 
    1.342271e-09, 1.350332e-09, 1.346497e-09, 1.357464e-09, 1.360164e-09, 
    1.362359e-09, 1.365164e-09, 1.365467e-09, 1.367129e-09, 1.364405e-09, 
    1.367022e-09, 1.357125e-09, 1.361547e-09, 1.34941e-09, 1.352365e-09, 
    1.351006e-09, 1.349515e-09, 1.354115e-09, 1.359017e-09, 1.359122e-09, 
    1.360693e-09, 1.365123e-09, 1.357509e-09, 1.381076e-09, 1.366522e-09, 
    1.344797e-09, 1.349258e-09, 1.349895e-09, 1.348167e-09, 1.359893e-09, 
    1.355644e-09, 1.367089e-09, 1.363996e-09, 1.369063e-09, 1.366545e-09, 
    1.366175e-09, 1.36294e-09, 1.360927e-09, 1.355839e-09, 1.3517e-09, 
    1.348417e-09, 1.349181e-09, 1.352787e-09, 1.359317e-09, 1.365494e-09, 
    1.364141e-09, 1.368678e-09, 1.356669e-09, 1.361705e-09, 1.359759e-09, 
    1.364833e-09, 1.353714e-09, 1.363183e-09, 1.351293e-09, 1.352336e-09, 
    1.35556e-09, 1.362047e-09, 1.363481e-09, 1.365014e-09, 1.364068e-09, 
    1.359483e-09, 1.358731e-09, 1.355482e-09, 1.354585e-09, 1.352109e-09, 
    1.350059e-09, 1.351932e-09, 1.353899e-09, 1.359485e-09, 1.364518e-09, 
    1.370007e-09, 1.37135e-09, 1.377763e-09, 1.372542e-09, 1.381157e-09, 
    1.373833e-09, 1.386511e-09, 1.363732e-09, 1.373618e-09, 1.355707e-09, 
    1.357636e-09, 1.361127e-09, 1.369131e-09, 1.36481e-09, 1.369864e-09, 
    1.358702e-09, 1.352911e-09, 1.351413e-09, 1.348617e-09, 1.351476e-09, 
    1.351244e-09, 1.35398e-09, 1.353101e-09, 1.35967e-09, 1.356141e-09, 
    1.366165e-09, 1.369824e-09, 1.380154e-09, 1.386487e-09, 1.392933e-09, 
    1.395779e-09, 1.396645e-09, 1.397008e-09 ;

 SOIL2_HR_S3 =
  9.481324e-11, 9.52305e-11, 9.514939e-11, 9.548595e-11, 9.529925e-11, 
    9.551963e-11, 9.489783e-11, 9.524707e-11, 9.502412e-11, 9.485079e-11, 
    9.61391e-11, 9.550096e-11, 9.68019e-11, 9.639493e-11, 9.741723e-11, 
    9.673858e-11, 9.755407e-11, 9.739764e-11, 9.786843e-11, 9.773356e-11, 
    9.833574e-11, 9.793068e-11, 9.864789e-11, 9.8239e-11, 9.830297e-11, 
    9.791731e-11, 9.562937e-11, 9.605965e-11, 9.560388e-11, 9.566523e-11, 
    9.56377e-11, 9.530311e-11, 9.51345e-11, 9.478134e-11, 9.484545e-11, 
    9.510483e-11, 9.569283e-11, 9.549322e-11, 9.599625e-11, 9.598489e-11, 
    9.654491e-11, 9.629241e-11, 9.723366e-11, 9.696614e-11, 9.773918e-11, 
    9.754477e-11, 9.773005e-11, 9.767387e-11, 9.773079e-11, 9.744566e-11, 
    9.756782e-11, 9.731693e-11, 9.63397e-11, 9.662691e-11, 9.577032e-11, 
    9.525528e-11, 9.491315e-11, 9.467038e-11, 9.47047e-11, 9.477013e-11, 
    9.510635e-11, 9.542245e-11, 9.566335e-11, 9.582449e-11, 9.598326e-11, 
    9.646387e-11, 9.671822e-11, 9.728775e-11, 9.718496e-11, 9.735909e-11, 
    9.752543e-11, 9.780471e-11, 9.775875e-11, 9.788179e-11, 9.735449e-11, 
    9.770494e-11, 9.712642e-11, 9.728465e-11, 9.602646e-11, 9.554707e-11, 
    9.534334e-11, 9.516498e-11, 9.473109e-11, 9.503073e-11, 9.491261e-11, 
    9.519362e-11, 9.537218e-11, 9.528386e-11, 9.582889e-11, 9.5617e-11, 
    9.67333e-11, 9.625248e-11, 9.750603e-11, 9.720606e-11, 9.757793e-11, 
    9.738817e-11, 9.771331e-11, 9.742069e-11, 9.792758e-11, 9.803796e-11, 
    9.796253e-11, 9.825226e-11, 9.740447e-11, 9.773006e-11, 9.528139e-11, 
    9.529579e-11, 9.536289e-11, 9.506794e-11, 9.504989e-11, 9.477958e-11, 
    9.50201e-11, 9.512253e-11, 9.538252e-11, 9.553631e-11, 9.56825e-11, 
    9.600394e-11, 9.636292e-11, 9.686489e-11, 9.722551e-11, 9.746724e-11, 
    9.731901e-11, 9.744987e-11, 9.730358e-11, 9.723502e-11, 9.79966e-11, 
    9.756897e-11, 9.821059e-11, 9.817509e-11, 9.788471e-11, 9.817908e-11, 
    9.53059e-11, 9.522302e-11, 9.493525e-11, 9.516046e-11, 9.475015e-11, 
    9.497982e-11, 9.511188e-11, 9.562143e-11, 9.573338e-11, 9.583719e-11, 
    9.604222e-11, 9.630533e-11, 9.676691e-11, 9.71685e-11, 9.75351e-11, 
    9.750824e-11, 9.75177e-11, 9.75996e-11, 9.739674e-11, 9.763291e-11, 
    9.767255e-11, 9.756891e-11, 9.817033e-11, 9.799851e-11, 9.817433e-11, 
    9.806245e-11, 9.524996e-11, 9.538943e-11, 9.531406e-11, 9.545578e-11, 
    9.535594e-11, 9.579987e-11, 9.593298e-11, 9.655576e-11, 9.630016e-11, 
    9.670693e-11, 9.634148e-11, 9.640624e-11, 9.672022e-11, 9.636122e-11, 
    9.714637e-11, 9.661408e-11, 9.760279e-11, 9.707126e-11, 9.763609e-11, 
    9.753352e-11, 9.770335e-11, 9.785545e-11, 9.80468e-11, 9.839987e-11, 
    9.831811e-11, 9.861337e-11, 9.559733e-11, 9.577823e-11, 9.576229e-11, 
    9.595159e-11, 9.609159e-11, 9.639503e-11, 9.68817e-11, 9.669869e-11, 
    9.703466e-11, 9.710211e-11, 9.659168e-11, 9.690508e-11, 9.589929e-11, 
    9.60618e-11, 9.596503e-11, 9.561161e-11, 9.674087e-11, 9.616134e-11, 
    9.723147e-11, 9.691752e-11, 9.783376e-11, 9.737811e-11, 9.82731e-11, 
    9.865572e-11, 9.90158e-11, 9.943662e-11, 9.587695e-11, 9.575403e-11, 
    9.59741e-11, 9.62786e-11, 9.65611e-11, 9.693667e-11, 9.697509e-11, 
    9.704546e-11, 9.722771e-11, 9.738094e-11, 9.706771e-11, 9.741936e-11, 
    9.60995e-11, 9.679117e-11, 9.570757e-11, 9.603388e-11, 9.626065e-11, 
    9.616116e-11, 9.667777e-11, 9.679953e-11, 9.729431e-11, 9.703854e-11, 
    9.85613e-11, 9.788759e-11, 9.975702e-11, 9.92346e-11, 9.571108e-11, 
    9.587652e-11, 9.645228e-11, 9.617833e-11, 9.696174e-11, 9.715458e-11, 
    9.731133e-11, 9.751173e-11, 9.753336e-11, 9.765209e-11, 9.745753e-11, 
    9.76444e-11, 9.693747e-11, 9.725338e-11, 9.638645e-11, 9.659747e-11, 
    9.650039e-11, 9.639391e-11, 9.672253e-11, 9.707265e-11, 9.708011e-11, 
    9.719238e-11, 9.750876e-11, 9.696492e-11, 9.864828e-11, 9.76087e-11, 
    9.605691e-11, 9.637557e-11, 9.642107e-11, 9.629763e-11, 9.713525e-11, 
    9.683175e-11, 9.764919e-11, 9.742826e-11, 9.779025e-11, 9.761037e-11, 
    9.758391e-11, 9.735288e-11, 9.720905e-11, 9.684567e-11, 9.655e-11, 
    9.631553e-11, 9.637005e-11, 9.662761e-11, 9.709406e-11, 9.753532e-11, 
    9.743866e-11, 9.776274e-11, 9.690494e-11, 9.726463e-11, 9.712562e-11, 
    9.74881e-11, 9.669383e-11, 9.737024e-11, 9.652094e-11, 9.65954e-11, 
    9.682573e-11, 9.728904e-11, 9.739153e-11, 9.750098e-11, 9.743344e-11, 
    9.71059e-11, 9.705223e-11, 9.682013e-11, 9.675605e-11, 9.657918e-11, 
    9.643276e-11, 9.656655e-11, 9.670705e-11, 9.710603e-11, 9.74656e-11, 
    9.785762e-11, 9.795355e-11, 9.841161e-11, 9.803874e-11, 9.865406e-11, 
    9.813095e-11, 9.903647e-11, 9.740941e-11, 9.811555e-11, 9.683621e-11, 
    9.697403e-11, 9.722333e-11, 9.779508e-11, 9.748639e-11, 9.78474e-11, 
    9.705013e-11, 9.66365e-11, 9.652946e-11, 9.632979e-11, 9.653403e-11, 
    9.651742e-11, 9.671285e-11, 9.665005e-11, 9.711928e-11, 9.686723e-11, 
    9.758325e-11, 9.784454e-11, 9.858243e-11, 9.903479e-11, 9.949523e-11, 
    9.969852e-11, 9.976039e-11, 9.978626e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.617555e-11, 2.629073e-11, 2.626834e-11, 2.636123e-11, 2.63097e-11, 
    2.637053e-11, 2.61989e-11, 2.62953e-11, 2.623376e-11, 2.618592e-11, 
    2.654151e-11, 2.636538e-11, 2.672445e-11, 2.661212e-11, 2.689429e-11, 
    2.670697e-11, 2.693206e-11, 2.688888e-11, 2.701883e-11, 2.69816e-11, 
    2.714781e-11, 2.703601e-11, 2.723397e-11, 2.712111e-11, 2.713877e-11, 
    2.703232e-11, 2.640082e-11, 2.651958e-11, 2.639378e-11, 2.641072e-11, 
    2.640312e-11, 2.631076e-11, 2.626423e-11, 2.616675e-11, 2.618445e-11, 
    2.625604e-11, 2.641833e-11, 2.636324e-11, 2.650208e-11, 2.649895e-11, 
    2.665352e-11, 2.658383e-11, 2.684362e-11, 2.676978e-11, 2.698315e-11, 
    2.692949e-11, 2.698063e-11, 2.696513e-11, 2.698084e-11, 2.690214e-11, 
    2.693586e-11, 2.68666e-11, 2.659688e-11, 2.667615e-11, 2.643972e-11, 
    2.629756e-11, 2.620313e-11, 2.613612e-11, 2.61456e-11, 2.616366e-11, 
    2.625646e-11, 2.63437e-11, 2.64102e-11, 2.645467e-11, 2.64985e-11, 
    2.663115e-11, 2.670136e-11, 2.685855e-11, 2.683018e-11, 2.687824e-11, 
    2.692416e-11, 2.700124e-11, 2.698855e-11, 2.702251e-11, 2.687697e-11, 
    2.69737e-11, 2.681402e-11, 2.68577e-11, 2.651042e-11, 2.63781e-11, 
    2.632187e-11, 2.627264e-11, 2.615288e-11, 2.623558e-11, 2.620298e-11, 
    2.628054e-11, 2.632983e-11, 2.630545e-11, 2.645589e-11, 2.63974e-11, 
    2.670552e-11, 2.65728e-11, 2.69188e-11, 2.683601e-11, 2.693864e-11, 
    2.688627e-11, 2.697601e-11, 2.689524e-11, 2.703515e-11, 2.706562e-11, 
    2.70448e-11, 2.712477e-11, 2.689077e-11, 2.698063e-11, 2.630477e-11, 
    2.630875e-11, 2.632727e-11, 2.624585e-11, 2.624087e-11, 2.616627e-11, 
    2.623265e-11, 2.626092e-11, 2.633268e-11, 2.637513e-11, 2.641548e-11, 
    2.650421e-11, 2.660329e-11, 2.674184e-11, 2.684137e-11, 2.690809e-11, 
    2.686718e-11, 2.69033e-11, 2.686292e-11, 2.6844e-11, 2.70542e-11, 
    2.693617e-11, 2.711327e-11, 2.710347e-11, 2.702332e-11, 2.710457e-11, 
    2.631154e-11, 2.628866e-11, 2.620923e-11, 2.627139e-11, 2.615814e-11, 
    2.622153e-11, 2.625799e-11, 2.639863e-11, 2.642953e-11, 2.645818e-11, 
    2.651477e-11, 2.658739e-11, 2.671479e-11, 2.682564e-11, 2.692683e-11, 
    2.691941e-11, 2.692202e-11, 2.694463e-11, 2.688863e-11, 2.695382e-11, 
    2.696476e-11, 2.693615e-11, 2.710215e-11, 2.705473e-11, 2.710326e-11, 
    2.707238e-11, 2.62961e-11, 2.633459e-11, 2.631379e-11, 2.63529e-11, 
    2.632535e-11, 2.644788e-11, 2.648462e-11, 2.665651e-11, 2.658596e-11, 
    2.669824e-11, 2.659737e-11, 2.661524e-11, 2.670191e-11, 2.660282e-11, 
    2.681953e-11, 2.667261e-11, 2.694551e-11, 2.67988e-11, 2.69547e-11, 
    2.692639e-11, 2.697326e-11, 2.701524e-11, 2.706806e-11, 2.716551e-11, 
    2.714294e-11, 2.722444e-11, 2.639198e-11, 2.64419e-11, 2.643751e-11, 
    2.648976e-11, 2.65284e-11, 2.661215e-11, 2.674648e-11, 2.669596e-11, 
    2.67887e-11, 2.680731e-11, 2.666643e-11, 2.675293e-11, 2.647532e-11, 
    2.652017e-11, 2.649347e-11, 2.639591e-11, 2.670761e-11, 2.654765e-11, 
    2.684302e-11, 2.675637e-11, 2.700926e-11, 2.688349e-11, 2.713052e-11, 
    2.723613e-11, 2.733551e-11, 2.745166e-11, 2.646915e-11, 2.643523e-11, 
    2.649597e-11, 2.658001e-11, 2.665799e-11, 2.676165e-11, 2.677226e-11, 
    2.679168e-11, 2.684198e-11, 2.688427e-11, 2.679782e-11, 2.689488e-11, 
    2.653058e-11, 2.672149e-11, 2.64224e-11, 2.651247e-11, 2.657506e-11, 
    2.65476e-11, 2.669019e-11, 2.67238e-11, 2.686036e-11, 2.678977e-11, 
    2.721007e-11, 2.702411e-11, 2.75401e-11, 2.73959e-11, 2.642337e-11, 
    2.646903e-11, 2.662795e-11, 2.655234e-11, 2.676857e-11, 2.68218e-11, 
    2.686506e-11, 2.692037e-11, 2.692634e-11, 2.695911e-11, 2.690541e-11, 
    2.695699e-11, 2.676187e-11, 2.684907e-11, 2.660978e-11, 2.666803e-11, 
    2.664123e-11, 2.661184e-11, 2.670255e-11, 2.679918e-11, 2.680124e-11, 
    2.683223e-11, 2.691955e-11, 2.676945e-11, 2.723407e-11, 2.694714e-11, 
    2.651883e-11, 2.660678e-11, 2.661934e-11, 2.658527e-11, 2.681646e-11, 
    2.673269e-11, 2.695831e-11, 2.689734e-11, 2.699725e-11, 2.69476e-11, 
    2.69403e-11, 2.687653e-11, 2.683683e-11, 2.673653e-11, 2.665492e-11, 
    2.659021e-11, 2.660526e-11, 2.667635e-11, 2.680509e-11, 2.692688e-11, 
    2.690021e-11, 2.698965e-11, 2.675289e-11, 2.685217e-11, 2.68138e-11, 
    2.691385e-11, 2.669462e-11, 2.688132e-11, 2.66469e-11, 2.666745e-11, 
    2.673103e-11, 2.685891e-11, 2.68872e-11, 2.691741e-11, 2.689876e-11, 
    2.680836e-11, 2.679355e-11, 2.672948e-11, 2.67118e-11, 2.666298e-11, 
    2.662257e-11, 2.665949e-11, 2.669827e-11, 2.68084e-11, 2.690764e-11, 
    2.701584e-11, 2.704232e-11, 2.716875e-11, 2.706584e-11, 2.723567e-11, 
    2.709129e-11, 2.734122e-11, 2.689213e-11, 2.708703e-11, 2.673392e-11, 
    2.677196e-11, 2.684077e-11, 2.699858e-11, 2.691338e-11, 2.701302e-11, 
    2.679297e-11, 2.66788e-11, 2.664926e-11, 2.659414e-11, 2.665052e-11, 
    2.664593e-11, 2.669987e-11, 2.668254e-11, 2.681205e-11, 2.674248e-11, 
    2.694011e-11, 2.701223e-11, 2.72159e-11, 2.734075e-11, 2.746784e-11, 
    2.752395e-11, 2.754103e-11, 2.754817e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, -1.28498e-20, 
    -1.541976e-20, 7.709882e-21, 1.541976e-20, -2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.003089e-36, -2.055969e-20, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -1.798972e-20, 1.28498e-20, -7.709882e-21, -1.28498e-20, 
    1.027984e-20, 1.541976e-20, -1.003089e-36, -2.569961e-21, 1.541976e-20, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 1.003089e-36, -2.569961e-21, 
    5.139921e-21, 0, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, 5.139921e-21, 0, 1.798972e-20, 
    -1.003089e-36, 1.027984e-20, 1.003089e-36, 1.28498e-20, 1.798972e-20, 
    7.709882e-21, -5.139921e-21, 0, 1.541976e-20, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, 1.28498e-20, -1.798972e-20, 
    1.027984e-20, 2.569961e-21, 2.569961e-21, 1.003089e-36, 2.569961e-21, 
    2.569961e-21, -1.28498e-20, 1.027984e-20, -2.569961e-21, 0, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, -1.003089e-36, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, 1.003089e-36, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, 0, 0, 7.709882e-21, -7.709882e-21, 
    -1.28498e-20, 1.28498e-20, 0, -1.027984e-20, -1.28498e-20, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 1.003089e-36, -5.139921e-21, 7.709882e-21, 
    -1.541976e-20, 1.541976e-20, -2.569961e-21, 1.541976e-20, 5.139921e-21, 
    2.569961e-21, 0, 1.003089e-36, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 1.28498e-20, -1.798972e-20, 2.312965e-20, 5.139921e-21, 
    7.709882e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 0, 1.003089e-36, 0, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 1.28498e-20, 1.541976e-20, -5.139921e-21, 1.003089e-36, 
    -1.003089e-36, -2.569961e-21, -1.027984e-20, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.541976e-20, 1.28498e-20, 
    -7.709882e-21, 7.709882e-21, 2.569961e-20, -7.709882e-21, -1.003089e-36, 
    -7.709882e-21, -1.027984e-20, -2.569961e-21, -1.027984e-20, 1.027984e-20, 
    7.709882e-21, -1.28498e-20, -1.28498e-20, -7.709882e-21, -1.541976e-20, 
    -7.709882e-21, -5.139921e-21, -2.055969e-20, 1.28498e-20, 1.541976e-20, 
    -1.003089e-36, 2.569961e-21, -2.569961e-21, -5.139921e-21, 1.798972e-20, 
    1.027984e-20, -1.003089e-36, -7.709882e-21, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, 1.28498e-20, 2.312965e-20, -2.312965e-20, 
    1.28498e-20, -1.28498e-20, 1.003089e-36, -7.709882e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, 1.28498e-20, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -7.709882e-21, -1.28498e-20, -1.798972e-20, 
    -2.569961e-21, -2.569961e-21, -1.798972e-20, 1.027984e-20, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 1.003089e-36, 5.139921e-21, 
    7.709882e-21, 1.003089e-36, 1.28498e-20, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -1.027984e-20, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, 1.541976e-20, -1.003089e-36, 
    2.569961e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 1.003089e-36, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, 1.027984e-20, -1.541976e-20, 1.003089e-36, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 1.28498e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    -5.139921e-21, 0, -7.709882e-21, 5.139921e-21, -7.709882e-21, 0, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 7.709882e-21, 1.28498e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 1.798972e-20, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    0, 2.569961e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -5.139921e-21, 1.541976e-20, 1.003089e-36, -1.541976e-20, 7.709882e-21, 
    1.28498e-20, 1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    1.003089e-36, 0, -5.139921e-21, -7.709882e-21, -1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    1.28498e-20, 5.139921e-21,
  -1.28498e-20, 7.709882e-21, -5.139921e-21, -2.055969e-20, -2.569961e-21, 
    2.569961e-21, -1.003089e-36, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 0, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -2.569961e-21, -1.28498e-20, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -1.28498e-20, 1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 0, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, -1.28498e-20, -1.28498e-20, -7.709882e-21, 0, 
    0, -1.027984e-20, -1.28498e-20, 0, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 0, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 0, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    -7.709882e-21, 0, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 0, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    1.003089e-36, -1.28498e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    -1.541976e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21, 0, 0, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -1.003089e-36, -5.139921e-21, -5.139921e-21, 1.541976e-20, -2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -1.28498e-20, 0, 1.28498e-20, -1.027984e-20, 
    1.28498e-20, 5.139921e-21, 1.28498e-20, 7.709882e-21, -7.709882e-21, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    -1.027984e-20, 1.003089e-36, -5.139921e-21, 5.139921e-21, 1.28498e-20, 
    7.709882e-21, 5.139921e-21, -2.569961e-21, -1.798972e-20, -1.541976e-20, 
    -2.569961e-21, 1.541976e-20, -7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 0, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, 0, -2.569961e-21, 0, 
    1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 1.003089e-36, 
    -7.709882e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, -1.28498e-20, 
    0, 1.027984e-20, 5.139921e-21, 0, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 7.709882e-21, -1.541976e-20, 2.055969e-20, 
    -2.569961e-21, 0, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 7.709882e-21, -1.003089e-36, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 2.055969e-20, 1.28498e-20, -2.569961e-21, 
    1.027984e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, 0, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -5.139921e-21, -7.709882e-21, 
    -1.027984e-20, -7.709882e-21, -1.28498e-20, -1.28498e-20, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, -1.28498e-20, 
    0, 1.027984e-20, 1.798972e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, 1.003089e-36, -5.139921e-21, 1.003089e-36, 
    -1.027984e-20, 2.569961e-21, -1.003089e-36, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, -1.28498e-20, -7.709882e-21, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    1.28498e-20, 2.055969e-20, -1.28498e-20, -1.003089e-36, -7.709882e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, -1.003089e-36, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, 0, 2.569961e-21, 2.569961e-21, 
    -1.003089e-36, 0, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -1.28498e-20, 1.541976e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, 2.055969e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 0, 1.027984e-20, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 0, 0, -2.569961e-21, -5.139921e-21, 
    1.027984e-20, 0, -7.709882e-21, -2.569961e-21, -1.28498e-20, 0,
  2.569961e-21, -5.139921e-21, 1.541976e-20, -2.569961e-21, 1.28498e-20, 
    -1.003089e-36, -1.027984e-20, 2.569961e-21, -5.139921e-21, 0, 
    7.709882e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, -2.055969e-20, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    -1.541976e-20, 0, -2.569961e-21, -1.027984e-20, -2.055969e-20, 
    1.003089e-36, 1.28498e-20, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 1.28498e-20, 0, 2.569961e-21, -1.28498e-20, -2.569961e-21, 
    0, 1.003089e-36, 2.569961e-21, -2.569961e-21, 0, 1.003089e-36, 0, 
    -5.139921e-21, 0, -1.28498e-20, -2.055969e-20, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 1.003089e-36, 1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 0, 2.569961e-21, 5.139921e-21, 7.709882e-21, 
    0, 0, 1.003089e-36, 1.28498e-20, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, 
    1.003089e-36, -1.027984e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, -1.003089e-36, 1.027984e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, 1.28498e-20, 
    2.569961e-21, 1.798972e-20, -1.28498e-20, -1.027984e-20, 7.709882e-21, 0, 
    7.709882e-21, -1.027984e-20, 1.003089e-36, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, 0, -7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -1.003089e-36, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -2.569961e-21, 1.541976e-20, -5.139921e-21, 
    1.28498e-20, 2.569961e-21, 1.28498e-20, -5.139921e-21, 1.28498e-20, 
    1.003089e-36, -1.003089e-36, -2.569961e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.027984e-20, -1.28498e-20, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    1.027984e-20, 1.027984e-20, -7.709882e-21, -1.003089e-36, -5.139921e-21, 
    5.139921e-21, 0, 2.569961e-21, 1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 0, -1.28498e-20, -1.027984e-20, -1.003089e-36, 
    -5.139921e-21, 0, 7.709882e-21, -1.541976e-20, -1.003089e-36, 0, 
    5.139921e-21, -1.027984e-20, -2.312965e-20, -7.709882e-21, -1.003089e-36, 
    2.569961e-21, 0, -1.027984e-20, 7.709882e-21, -2.569961e-21, 
    -1.003089e-36, -1.798972e-20, 2.055969e-20, 1.003089e-36, 1.027984e-20, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 1.003089e-36, 
    -1.027984e-20, -7.709882e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, -1.28498e-20, -5.139921e-21, -5.139921e-21, 0, 
    -1.027984e-20, 1.798972e-20, 1.003089e-36, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 1.003089e-36, 
    5.139921e-21, -1.541976e-20, 1.28498e-20, 1.28498e-20, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, 1.003089e-36, -5.139921e-21, 0, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -7.709882e-21, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, 1.003089e-36, -2.569961e-21, 0, -7.709882e-21, 
    1.027984e-20, -1.28498e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, 1.003089e-36, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 1.798972e-20, 2.569961e-21, 1.003089e-36, 
    1.027984e-20, 2.055969e-20, 1.28498e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 2.569961e-21, 0, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, -1.003089e-36, 
    0, 1.027984e-20, -1.003089e-36, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    0, 1.027984e-20, -2.569961e-21, 1.798972e-20, -5.139921e-21, 
    -1.798972e-20, -1.027984e-20, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    2.569961e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -1.798972e-20, 0, 1.003089e-36, -7.709882e-21, 
    5.139921e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.28498e-20, 0, -1.798972e-20, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 1.28498e-20, 
    1.28498e-20, 5.139921e-21, -2.569961e-21, -1.027984e-20, 7.709882e-21, 0, 
    1.027984e-20, -2.569961e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    1.798972e-20,
  -5.139921e-21, 2.569961e-21, -2.569961e-21, 0, 1.003089e-36, 7.709882e-21, 
    7.709882e-21, 1.027984e-20, 2.312965e-20, 1.28498e-20, 5.139921e-21, 
    1.28498e-20, 7.709882e-21, 2.055969e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, 1.541976e-20, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, 1.003089e-36, -1.541976e-20, 
    7.709882e-21, -1.027984e-20, 1.28498e-20, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.28498e-20, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, 1.798972e-20, 2.569961e-21, 
    1.541976e-20, -7.709882e-21, 5.139921e-21, -7.709882e-21, -1.541976e-20, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, -1.541976e-20, -7.709882e-21, 
    -1.027984e-20, 1.28498e-20, 7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -1.28498e-20, 2.312965e-20, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 0, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -1.003089e-36, -7.709882e-21, -1.798972e-20, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, 1.798972e-20, -5.139921e-21, -5.139921e-21, -1.003089e-36, 
    -1.798972e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -1.027984e-20, 1.28498e-20, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 0, 
    -5.139921e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 0, 
    2.055969e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    1.027984e-20, -2.569961e-21, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    -1.541976e-20, 7.709882e-21, 1.28498e-20, 7.709882e-21, -7.709882e-21, 
    1.027984e-20, 1.28498e-20, 1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 1.798972e-20, 1.541976e-20, -7.709882e-21, -5.139921e-21, 
    1.003089e-36, 1.027984e-20, 2.569961e-21, 1.027984e-20, 0, 1.003089e-36, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, -2.569961e-21, 
    -1.28498e-20, -2.569961e-21, 5.139921e-21, 1.003089e-36, -7.709882e-21, 
    2.569961e-20, -1.541976e-20, -5.139921e-21, 2.569961e-21, 1.541976e-20, 
    0, -2.569961e-21, -1.003089e-36, -7.709882e-21, -2.569961e-21, 0, 
    -2.569961e-21, -7.709882e-21, 1.541976e-20, 2.569961e-21, -2.569961e-21, 
    1.003089e-36, 5.139921e-21, -1.003089e-36, 1.027984e-20, 1.003089e-36, 
    2.055969e-20, -2.055969e-20, 1.003089e-36, -7.709882e-21, -1.798972e-20, 
    1.541976e-20, -1.003089e-36, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, -1.003089e-36, 2.569961e-21, -1.541976e-20, 1.798972e-20, 
    2.055969e-20, -2.569961e-21, 1.003089e-36, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 2.569961e-20, 1.027984e-20, 1.003089e-36, 
    -2.569961e-21, 0, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, -1.003089e-36, -2.055969e-20, 
    0, -2.312965e-20, -1.28498e-20, -1.003089e-36, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.541976e-20, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, 2.569961e-21, -2.826957e-20, 7.709882e-21, 
    1.28498e-20, 2.569961e-21, 1.027984e-20, -2.569961e-21, -1.027984e-20, 
    1.027984e-20, -1.798972e-20, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    2.312965e-20, -1.003089e-36, 1.28498e-20, 5.139921e-21, 1.003089e-36, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, -2.826957e-20, 0, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 1.28498e-20, 2.569961e-21, -1.027984e-20, -7.709882e-21, 
    2.569961e-21, -1.003089e-36, -2.055969e-20, 5.139921e-21, -1.28498e-20, 
    1.541976e-20, -7.709882e-21, -5.139921e-21, 1.28498e-20, 1.28498e-20, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -1.003089e-36, -5.139921e-21, 1.541976e-20, 7.709882e-21, 0, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    1.003089e-36, 5.139921e-21, -5.139921e-21, 2.569961e-21, -2.055969e-20, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, 0, 1.28498e-20, 5.139921e-21, -1.003089e-36, 
    -1.541976e-20, 2.569961e-21, 1.027984e-20, 2.312965e-20, 1.28498e-20, 
    7.709882e-21, 5.139921e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 1.798972e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21,
  1.027984e-20, 7.709882e-21, -5.139921e-21, -5.139921e-21, 1.003089e-36, 
    -2.055969e-20, 7.709882e-21, 2.055969e-20, -1.027984e-20, -2.055969e-20, 
    -1.28498e-20, -5.139921e-21, -1.003089e-36, 2.312965e-20, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 1.541976e-20, -5.139921e-21, 
    -2.312965e-20, -1.798972e-20, 2.569961e-21, -1.28498e-20, -1.28498e-20, 
    -2.569961e-21, 1.027984e-20, -2.055969e-20, -1.003089e-36, 7.709882e-21, 
    2.569961e-21, 1.798972e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, -2.055969e-20, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, 2.055969e-20, -2.569961e-21, 1.798972e-20, -1.027984e-20, 
    -1.798972e-20, 2.569961e-21, -2.569961e-21, 0, 1.28498e-20, 1.027984e-20, 
    -1.798972e-20, 1.003089e-36, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    1.28498e-20, 1.027984e-20, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, 1.003089e-36, 1.027984e-20, -7.709882e-21, 2.312965e-20, 
    7.709882e-21, 2.826957e-20, -1.003089e-36, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, -1.003089e-36, 
    -2.055969e-20, 1.541976e-20, 1.003089e-36, -1.003089e-36, -1.027984e-20, 
    1.003089e-36, -7.709882e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -2.312965e-20, 7.709882e-21, 1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -1.798972e-20, 7.709882e-21, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    -1.798972e-20, 7.709882e-21, 1.027984e-20, 0, 7.709882e-21, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, -1.798972e-20, 1.027984e-20, 
    7.709882e-21, 1.003089e-36, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -3.009266e-36, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 0, 7.709882e-21, -1.027984e-20, -3.009266e-36, 
    1.541976e-20, 1.541976e-20, 2.569961e-21, -7.709882e-21, 5.139921e-21, 0, 
    2.055969e-20, -1.541976e-20, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.798972e-20, 
    -2.569961e-21, -1.541976e-20, -2.569961e-21, 1.027984e-20, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, 3.009266e-36, 1.027984e-20, -5.139921e-21, 
    1.798972e-20, 2.569961e-21, 1.28498e-20, 1.28498e-20, 1.28498e-20, 
    1.027984e-20, -1.541976e-20, -7.709882e-21, -5.139921e-21, 1.003089e-36, 
    -1.003089e-36, 1.027984e-20, 0, -1.003089e-36, 0, 2.055969e-20, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 1.798972e-20, 
    -1.003089e-36, -7.709882e-21, -1.28498e-20, -1.798972e-20, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, 2.312965e-20, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, 1.003089e-36, 1.28498e-20, 1.027984e-20, 2.312965e-20, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, -1.003089e-36, 
    -1.003089e-36, 2.569961e-21, 7.709882e-21, -2.569961e-21, 1.003089e-36, 
    -7.709882e-21, -1.28498e-20, -5.139921e-21, 1.28498e-20, -1.28498e-20, 
    -5.139921e-21, 7.709882e-21, 1.28498e-20, -2.569961e-21, -2.312965e-20, 
    2.569961e-21, -2.569961e-21, 2.569961e-20, -1.003089e-36, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, 1.003089e-36, 1.28498e-20, -1.28498e-20, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, -2.569961e-20, 2.826957e-20, 2.312965e-20, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, -7.709882e-21, 
    -1.027984e-20, 1.541976e-20, -2.569961e-21, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -1.003089e-36, 0, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 1.28498e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, 5.139921e-21, 1.28498e-20, -1.003089e-36, 
    1.003089e-36, -1.798972e-20, 2.569961e-21, 7.709882e-21, -2.312965e-20, 
    -1.28498e-20, -1.027984e-20, 7.709882e-21, 7.709882e-21, -2.312965e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, 1.027984e-20, -1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -2.569961e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    1.541976e-20, -2.055969e-20, -5.139921e-21, 1.027984e-20, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, 1.003089e-36, -1.28498e-20, 
    5.139921e-21, -1.027984e-20, 7.709882e-21, -1.027984e-20, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, -2.826957e-20, 2.569961e-21, 5.139921e-21, 2.055969e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.287991e-12, 5.311258e-12, 5.306735e-12, 5.325501e-12, 5.315091e-12, 
    5.327379e-12, 5.292708e-12, 5.312182e-12, 5.29975e-12, 5.290085e-12, 
    5.361921e-12, 5.326338e-12, 5.398879e-12, 5.376186e-12, 5.43319e-12, 
    5.395348e-12, 5.44082e-12, 5.432097e-12, 5.458349e-12, 5.450828e-12, 
    5.484406e-12, 5.46182e-12, 5.501811e-12, 5.479012e-12, 5.482579e-12, 
    5.461075e-12, 5.333499e-12, 5.357491e-12, 5.332077e-12, 5.335499e-12, 
    5.333963e-12, 5.315306e-12, 5.305904e-12, 5.286212e-12, 5.289787e-12, 
    5.30425e-12, 5.337037e-12, 5.325907e-12, 5.353956e-12, 5.353323e-12, 
    5.384549e-12, 5.37047e-12, 5.422954e-12, 5.408037e-12, 5.451142e-12, 
    5.440302e-12, 5.450633e-12, 5.4475e-12, 5.450674e-12, 5.434775e-12, 
    5.441587e-12, 5.427597e-12, 5.373107e-12, 5.389121e-12, 5.341358e-12, 
    5.312639e-12, 5.293562e-12, 5.280025e-12, 5.281939e-12, 5.285587e-12, 
    5.304335e-12, 5.321961e-12, 5.335393e-12, 5.344379e-12, 5.353231e-12, 
    5.380031e-12, 5.394213e-12, 5.42597e-12, 5.420239e-12, 5.429948e-12, 
    5.439223e-12, 5.454796e-12, 5.452232e-12, 5.459094e-12, 5.429692e-12, 
    5.449233e-12, 5.416974e-12, 5.425797e-12, 5.35564e-12, 5.32891e-12, 
    5.317549e-12, 5.307604e-12, 5.28341e-12, 5.300118e-12, 5.293532e-12, 
    5.309201e-12, 5.319157e-12, 5.314233e-12, 5.344624e-12, 5.332809e-12, 
    5.395054e-12, 5.368243e-12, 5.438141e-12, 5.421415e-12, 5.442151e-12, 
    5.43157e-12, 5.449699e-12, 5.433383e-12, 5.461647e-12, 5.467802e-12, 
    5.463596e-12, 5.479751e-12, 5.432478e-12, 5.450633e-12, 5.314095e-12, 
    5.314898e-12, 5.31864e-12, 5.302193e-12, 5.301187e-12, 5.286114e-12, 
    5.299526e-12, 5.305237e-12, 5.319734e-12, 5.32831e-12, 5.336462e-12, 
    5.354385e-12, 5.374402e-12, 5.402392e-12, 5.4225e-12, 5.435978e-12, 
    5.427713e-12, 5.43501e-12, 5.426853e-12, 5.42303e-12, 5.465496e-12, 
    5.441651e-12, 5.477428e-12, 5.475448e-12, 5.459257e-12, 5.475671e-12, 
    5.315462e-12, 5.31084e-12, 5.294795e-12, 5.307352e-12, 5.284473e-12, 
    5.29728e-12, 5.304643e-12, 5.333056e-12, 5.339298e-12, 5.345087e-12, 
    5.356519e-12, 5.37119e-12, 5.396928e-12, 5.419321e-12, 5.439763e-12, 
    5.438265e-12, 5.438792e-12, 5.443359e-12, 5.432047e-12, 5.445216e-12, 
    5.447426e-12, 5.441648e-12, 5.475183e-12, 5.465602e-12, 5.475406e-12, 
    5.469168e-12, 5.312343e-12, 5.320119e-12, 5.315917e-12, 5.323819e-12, 
    5.318252e-12, 5.343006e-12, 5.350428e-12, 5.385154e-12, 5.370902e-12, 
    5.393584e-12, 5.373206e-12, 5.376817e-12, 5.394325e-12, 5.374307e-12, 
    5.418087e-12, 5.388406e-12, 5.443537e-12, 5.413899e-12, 5.445394e-12, 
    5.439674e-12, 5.449144e-12, 5.457625e-12, 5.468294e-12, 5.487982e-12, 
    5.483423e-12, 5.499887e-12, 5.331712e-12, 5.341799e-12, 5.34091e-12, 
    5.351466e-12, 5.359272e-12, 5.376192e-12, 5.403329e-12, 5.393124e-12, 
    5.411858e-12, 5.415619e-12, 5.387157e-12, 5.404632e-12, 5.348549e-12, 
    5.357611e-12, 5.352215e-12, 5.332508e-12, 5.395476e-12, 5.363161e-12, 
    5.422832e-12, 5.405326e-12, 5.456416e-12, 5.431009e-12, 5.480913e-12, 
    5.502248e-12, 5.522325e-12, 5.54579e-12, 5.347303e-12, 5.34045e-12, 
    5.352721e-12, 5.3697e-12, 5.385452e-12, 5.406394e-12, 5.408536e-12, 
    5.41246e-12, 5.422622e-12, 5.431166e-12, 5.413701e-12, 5.433308e-12, 
    5.359713e-12, 5.398281e-12, 5.337859e-12, 5.356054e-12, 5.368699e-12, 
    5.363152e-12, 5.391958e-12, 5.398747e-12, 5.426336e-12, 5.412074e-12, 
    5.496983e-12, 5.459417e-12, 5.563655e-12, 5.534526e-12, 5.338055e-12, 
    5.347279e-12, 5.379384e-12, 5.364109e-12, 5.407792e-12, 5.418545e-12, 
    5.427285e-12, 5.438459e-12, 5.439665e-12, 5.446285e-12, 5.435437e-12, 
    5.445857e-12, 5.406439e-12, 5.424054e-12, 5.375714e-12, 5.38748e-12, 
    5.382067e-12, 5.37613e-12, 5.394454e-12, 5.413976e-12, 5.414392e-12, 
    5.420652e-12, 5.438294e-12, 5.407969e-12, 5.501832e-12, 5.443866e-12, 
    5.357338e-12, 5.375107e-12, 5.377644e-12, 5.370761e-12, 5.417467e-12, 
    5.400544e-12, 5.446124e-12, 5.433805e-12, 5.453989e-12, 5.44396e-12, 
    5.442484e-12, 5.429602e-12, 5.421582e-12, 5.40132e-12, 5.384833e-12, 
    5.371759e-12, 5.374799e-12, 5.38916e-12, 5.41517e-12, 5.439774e-12, 
    5.434385e-12, 5.452455e-12, 5.404625e-12, 5.424681e-12, 5.41693e-12, 
    5.437142e-12, 5.392853e-12, 5.43057e-12, 5.383213e-12, 5.387365e-12, 
    5.400208e-12, 5.426042e-12, 5.431757e-12, 5.43786e-12, 5.434094e-12, 
    5.41583e-12, 5.412838e-12, 5.399895e-12, 5.396322e-12, 5.38646e-12, 
    5.378296e-12, 5.385756e-12, 5.39359e-12, 5.415837e-12, 5.435887e-12, 
    5.457746e-12, 5.463095e-12, 5.488636e-12, 5.467846e-12, 5.502156e-12, 
    5.472987e-12, 5.523478e-12, 5.432754e-12, 5.472128e-12, 5.400792e-12, 
    5.408477e-12, 5.422378e-12, 5.454259e-12, 5.437047e-12, 5.457176e-12, 
    5.412721e-12, 5.389657e-12, 5.383688e-12, 5.372554e-12, 5.383942e-12, 
    5.383017e-12, 5.393914e-12, 5.390412e-12, 5.416576e-12, 5.402522e-12, 
    5.442447e-12, 5.457017e-12, 5.498161e-12, 5.523384e-12, 5.549059e-12, 
    5.560394e-12, 5.563844e-12, 5.565286e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.199234e-11, 3.213311e-11, 3.210575e-11, 3.221928e-11, 3.21563e-11, 
    3.223065e-11, 3.202088e-11, 3.21387e-11, 3.206349e-11, 3.200501e-11, 
    3.243962e-11, 3.222435e-11, 3.266322e-11, 3.252593e-11, 3.28708e-11, 
    3.264185e-11, 3.291696e-11, 3.286419e-11, 3.302301e-11, 3.297751e-11, 
    3.318066e-11, 3.304401e-11, 3.328596e-11, 3.314802e-11, 3.31696e-11, 
    3.30395e-11, 3.226767e-11, 3.241282e-11, 3.225907e-11, 3.227977e-11, 
    3.227048e-11, 3.21576e-11, 3.210072e-11, 3.198158e-11, 3.200321e-11, 
    3.209071e-11, 3.228907e-11, 3.222174e-11, 3.239143e-11, 3.23876e-11, 
    3.257652e-11, 3.249134e-11, 3.280887e-11, 3.271862e-11, 3.297941e-11, 
    3.291382e-11, 3.297633e-11, 3.295738e-11, 3.297658e-11, 3.288039e-11, 
    3.29216e-11, 3.283696e-11, 3.25073e-11, 3.260419e-11, 3.231522e-11, 
    3.214147e-11, 3.202605e-11, 3.194415e-11, 3.195573e-11, 3.19778e-11, 
    3.209123e-11, 3.219786e-11, 3.227913e-11, 3.233349e-11, 3.238705e-11, 
    3.254919e-11, 3.263499e-11, 3.282712e-11, 3.279245e-11, 3.285119e-11, 
    3.29073e-11, 3.300151e-11, 3.298601e-11, 3.302751e-11, 3.284964e-11, 
    3.296786e-11, 3.277269e-11, 3.282607e-11, 3.240163e-11, 3.22399e-11, 
    3.217118e-11, 3.2111e-11, 3.196463e-11, 3.206571e-11, 3.202587e-11, 
    3.212066e-11, 3.21809e-11, 3.215111e-11, 3.233497e-11, 3.226349e-11, 
    3.264008e-11, 3.247787e-11, 3.290076e-11, 3.279956e-11, 3.292501e-11, 
    3.2861e-11, 3.297068e-11, 3.287197e-11, 3.304296e-11, 3.30802e-11, 
    3.305475e-11, 3.315249e-11, 3.286649e-11, 3.297633e-11, 3.215028e-11, 
    3.215513e-11, 3.217777e-11, 3.207827e-11, 3.207218e-11, 3.198099e-11, 
    3.206213e-11, 3.209668e-11, 3.218439e-11, 3.223627e-11, 3.228559e-11, 
    3.239403e-11, 3.251513e-11, 3.268447e-11, 3.280612e-11, 3.288767e-11, 
    3.283766e-11, 3.288181e-11, 3.283246e-11, 3.280933e-11, 3.306625e-11, 
    3.292198e-11, 3.313844e-11, 3.312646e-11, 3.30285e-11, 3.312781e-11, 
    3.215855e-11, 3.213058e-11, 3.203351e-11, 3.210948e-11, 3.197106e-11, 
    3.204854e-11, 3.209309e-11, 3.226499e-11, 3.230275e-11, 3.233777e-11, 
    3.240694e-11, 3.24957e-11, 3.265141e-11, 3.278689e-11, 3.291056e-11, 
    3.29015e-11, 3.290469e-11, 3.293232e-11, 3.286389e-11, 3.294356e-11, 
    3.295693e-11, 3.292197e-11, 3.312485e-11, 3.306689e-11, 3.31262e-11, 
    3.308846e-11, 3.213967e-11, 3.218672e-11, 3.21613e-11, 3.22091e-11, 
    3.217543e-11, 3.232519e-11, 3.237009e-11, 3.258019e-11, 3.249396e-11, 
    3.263118e-11, 3.25079e-11, 3.252974e-11, 3.263567e-11, 3.251456e-11, 
    3.277943e-11, 3.259986e-11, 3.29334e-11, 3.275409e-11, 3.294463e-11, 
    3.291003e-11, 3.296732e-11, 3.301863e-11, 3.308318e-11, 3.320229e-11, 
    3.317471e-11, 3.327431e-11, 3.225686e-11, 3.231788e-11, 3.231251e-11, 
    3.237637e-11, 3.24236e-11, 3.252596e-11, 3.269014e-11, 3.26284e-11, 
    3.274174e-11, 3.276449e-11, 3.25923e-11, 3.269803e-11, 3.235872e-11, 
    3.241355e-11, 3.23809e-11, 3.226167e-11, 3.264263e-11, 3.244712e-11, 
    3.280813e-11, 3.270222e-11, 3.301132e-11, 3.28576e-11, 3.315952e-11, 
    3.32886e-11, 3.341007e-11, 3.355203e-11, 3.235119e-11, 3.230972e-11, 
    3.238396e-11, 3.248668e-11, 3.258199e-11, 3.270869e-11, 3.272165e-11, 
    3.274538e-11, 3.280686e-11, 3.285856e-11, 3.275289e-11, 3.287151e-11, 
    3.242627e-11, 3.26596e-11, 3.229405e-11, 3.240413e-11, 3.248063e-11, 
    3.244707e-11, 3.262134e-11, 3.266242e-11, 3.282933e-11, 3.274305e-11, 
    3.325674e-11, 3.302947e-11, 3.366012e-11, 3.348388e-11, 3.229524e-11, 
    3.235104e-11, 3.254527e-11, 3.245286e-11, 3.271714e-11, 3.278219e-11, 
    3.283507e-11, 3.290268e-11, 3.290997e-11, 3.295003e-11, 3.288439e-11, 
    3.294743e-11, 3.270895e-11, 3.281552e-11, 3.252307e-11, 3.259425e-11, 
    3.256151e-11, 3.252559e-11, 3.263645e-11, 3.275456e-11, 3.275707e-11, 
    3.279495e-11, 3.290168e-11, 3.271821e-11, 3.328609e-11, 3.293539e-11, 
    3.24119e-11, 3.25194e-11, 3.253475e-11, 3.249311e-11, 3.277567e-11, 
    3.267329e-11, 3.294905e-11, 3.287452e-11, 3.299663e-11, 3.293596e-11, 
    3.292703e-11, 3.284909e-11, 3.280057e-11, 3.267799e-11, 3.257824e-11, 
    3.249914e-11, 3.251753e-11, 3.260442e-11, 3.276178e-11, 3.291064e-11, 
    3.287803e-11, 3.298736e-11, 3.269798e-11, 3.281932e-11, 3.277242e-11, 
    3.289471e-11, 3.262676e-11, 3.285494e-11, 3.256843e-11, 3.259356e-11, 
    3.267126e-11, 3.282756e-11, 3.286213e-11, 3.289905e-11, 3.287627e-11, 
    3.276577e-11, 3.274767e-11, 3.266937e-11, 3.264775e-11, 3.258809e-11, 
    3.253869e-11, 3.258382e-11, 3.263122e-11, 3.276582e-11, 3.288712e-11, 
    3.301936e-11, 3.305172e-11, 3.320625e-11, 3.308047e-11, 3.328804e-11, 
    3.311157e-11, 3.341704e-11, 3.286816e-11, 3.310638e-11, 3.267479e-11, 
    3.272129e-11, 3.280539e-11, 3.299827e-11, 3.289413e-11, 3.301591e-11, 
    3.274696e-11, 3.260742e-11, 3.257131e-11, 3.250395e-11, 3.257285e-11, 
    3.256725e-11, 3.263318e-11, 3.261199e-11, 3.277029e-11, 3.268526e-11, 
    3.29268e-11, 3.301495e-11, 3.326388e-11, 3.341647e-11, 3.357181e-11, 
    3.364038e-11, 3.366125e-11, 3.366998e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.356892e-08, 6.384848e-08, 6.379413e-08, 6.401962e-08, 6.389453e-08, 
    6.404218e-08, 6.362559e-08, 6.385958e-08, 6.37102e-08, 6.359408e-08, 
    6.445721e-08, 6.402967e-08, 6.490126e-08, 6.462861e-08, 6.531352e-08, 
    6.485884e-08, 6.54052e-08, 6.530039e-08, 6.561581e-08, 6.552545e-08, 
    6.592889e-08, 6.565751e-08, 6.613801e-08, 6.586408e-08, 6.590693e-08, 
    6.564856e-08, 6.41157e-08, 6.440398e-08, 6.409863e-08, 6.413973e-08, 
    6.412129e-08, 6.389712e-08, 6.378416e-08, 6.354755e-08, 6.35905e-08, 
    6.376428e-08, 6.415822e-08, 6.402449e-08, 6.436151e-08, 6.43539e-08, 
    6.472909e-08, 6.455993e-08, 6.519053e-08, 6.50113e-08, 6.552921e-08, 
    6.539896e-08, 6.55231e-08, 6.548546e-08, 6.552359e-08, 6.533256e-08, 
    6.541441e-08, 6.524632e-08, 6.459161e-08, 6.478403e-08, 6.421014e-08, 
    6.386507e-08, 6.363586e-08, 6.347321e-08, 6.34962e-08, 6.354004e-08, 
    6.37653e-08, 6.397708e-08, 6.413847e-08, 6.424643e-08, 6.43528e-08, 
    6.46748e-08, 6.484521e-08, 6.522678e-08, 6.515791e-08, 6.527457e-08, 
    6.538601e-08, 6.557312e-08, 6.554232e-08, 6.562475e-08, 6.527149e-08, 
    6.550627e-08, 6.511868e-08, 6.522469e-08, 6.438174e-08, 6.406056e-08, 
    6.392407e-08, 6.380458e-08, 6.351388e-08, 6.371463e-08, 6.36355e-08, 
    6.382376e-08, 6.394339e-08, 6.388422e-08, 6.424938e-08, 6.410742e-08, 
    6.485531e-08, 6.453317e-08, 6.537302e-08, 6.517205e-08, 6.542118e-08, 
    6.529405e-08, 6.551188e-08, 6.531584e-08, 6.565543e-08, 6.572938e-08, 
    6.567885e-08, 6.587296e-08, 6.530497e-08, 6.55231e-08, 6.388257e-08, 
    6.389222e-08, 6.393717e-08, 6.373956e-08, 6.372747e-08, 6.354637e-08, 
    6.370751e-08, 6.377613e-08, 6.395032e-08, 6.405336e-08, 6.415131e-08, 
    6.436666e-08, 6.460716e-08, 6.494347e-08, 6.518507e-08, 6.534702e-08, 
    6.524771e-08, 6.533539e-08, 6.523738e-08, 6.519144e-08, 6.570168e-08, 
    6.541517e-08, 6.584504e-08, 6.582125e-08, 6.562671e-08, 6.582393e-08, 
    6.389899e-08, 6.384346e-08, 6.365067e-08, 6.380154e-08, 6.352665e-08, 
    6.368052e-08, 6.376901e-08, 6.411039e-08, 6.418539e-08, 6.425494e-08, 
    6.43923e-08, 6.456858e-08, 6.487782e-08, 6.514688e-08, 6.539249e-08, 
    6.537449e-08, 6.538083e-08, 6.54357e-08, 6.529979e-08, 6.545802e-08, 
    6.548457e-08, 6.541514e-08, 6.581807e-08, 6.570296e-08, 6.582075e-08, 
    6.574579e-08, 6.386151e-08, 6.395495e-08, 6.390446e-08, 6.39994e-08, 
    6.393252e-08, 6.422994e-08, 6.431911e-08, 6.473636e-08, 6.456511e-08, 
    6.483764e-08, 6.45928e-08, 6.463618e-08, 6.484655e-08, 6.460603e-08, 
    6.513206e-08, 6.477543e-08, 6.543784e-08, 6.508173e-08, 6.546015e-08, 
    6.539143e-08, 6.55052e-08, 6.560711e-08, 6.573531e-08, 6.597185e-08, 
    6.591708e-08, 6.611489e-08, 6.409424e-08, 6.421543e-08, 6.420476e-08, 
    6.433159e-08, 6.442539e-08, 6.462868e-08, 6.495473e-08, 6.483211e-08, 
    6.505721e-08, 6.51024e-08, 6.476043e-08, 6.497039e-08, 6.429654e-08, 
    6.440542e-08, 6.434059e-08, 6.41038e-08, 6.486038e-08, 6.447211e-08, 
    6.518906e-08, 6.497873e-08, 6.559258e-08, 6.528731e-08, 6.588692e-08, 
    6.614327e-08, 6.638449e-08, 6.666644e-08, 6.428157e-08, 6.419923e-08, 
    6.434667e-08, 6.455067e-08, 6.473994e-08, 6.499156e-08, 6.50173e-08, 
    6.506445e-08, 6.518654e-08, 6.528921e-08, 6.507936e-08, 6.531494e-08, 
    6.443068e-08, 6.489408e-08, 6.41681e-08, 6.438672e-08, 6.453865e-08, 
    6.447199e-08, 6.48181e-08, 6.489968e-08, 6.523117e-08, 6.505981e-08, 
    6.608001e-08, 6.562864e-08, 6.688109e-08, 6.653109e-08, 6.417046e-08, 
    6.428129e-08, 6.466703e-08, 6.448349e-08, 6.500836e-08, 6.513755e-08, 
    6.524257e-08, 6.537682e-08, 6.539132e-08, 6.547086e-08, 6.534052e-08, 
    6.546571e-08, 6.49921e-08, 6.520374e-08, 6.462293e-08, 6.47643e-08, 
    6.469926e-08, 6.462793e-08, 6.484809e-08, 6.508266e-08, 6.508766e-08, 
    6.516288e-08, 6.537484e-08, 6.501048e-08, 6.613828e-08, 6.54418e-08, 
    6.440214e-08, 6.461564e-08, 6.464612e-08, 6.456342e-08, 6.51246e-08, 
    6.492127e-08, 6.546892e-08, 6.532091e-08, 6.556343e-08, 6.544292e-08, 
    6.542518e-08, 6.527041e-08, 6.517404e-08, 6.493059e-08, 6.47325e-08, 
    6.457542e-08, 6.461194e-08, 6.478449e-08, 6.509701e-08, 6.539263e-08, 
    6.532787e-08, 6.5545e-08, 6.49703e-08, 6.521128e-08, 6.511815e-08, 
    6.5361e-08, 6.482886e-08, 6.528204e-08, 6.471303e-08, 6.476292e-08, 
    6.491723e-08, 6.522764e-08, 6.52963e-08, 6.536963e-08, 6.532438e-08, 
    6.510494e-08, 6.506898e-08, 6.491348e-08, 6.487055e-08, 6.475205e-08, 
    6.465395e-08, 6.474359e-08, 6.483771e-08, 6.510503e-08, 6.534592e-08, 
    6.560856e-08, 6.567284e-08, 6.597972e-08, 6.572991e-08, 6.614216e-08, 
    6.579169e-08, 6.639835e-08, 6.530828e-08, 6.578136e-08, 6.492425e-08, 
    6.501659e-08, 6.518361e-08, 6.556667e-08, 6.535986e-08, 6.560172e-08, 
    6.506757e-08, 6.479046e-08, 6.471874e-08, 6.458497e-08, 6.47218e-08, 
    6.471067e-08, 6.484161e-08, 6.479953e-08, 6.51139e-08, 6.494503e-08, 
    6.542474e-08, 6.55998e-08, 6.609416e-08, 6.639722e-08, 6.67057e-08, 
    6.684189e-08, 6.688335e-08, 6.690068e-08 ;

 SOILC_LOSS =
  6.356892e-08, 6.384848e-08, 6.379413e-08, 6.401962e-08, 6.389453e-08, 
    6.404218e-08, 6.362559e-08, 6.385958e-08, 6.37102e-08, 6.359408e-08, 
    6.445721e-08, 6.402967e-08, 6.490126e-08, 6.462861e-08, 6.531352e-08, 
    6.485884e-08, 6.54052e-08, 6.530039e-08, 6.561581e-08, 6.552545e-08, 
    6.592889e-08, 6.565751e-08, 6.613801e-08, 6.586408e-08, 6.590693e-08, 
    6.564856e-08, 6.41157e-08, 6.440398e-08, 6.409863e-08, 6.413973e-08, 
    6.412129e-08, 6.389712e-08, 6.378416e-08, 6.354755e-08, 6.35905e-08, 
    6.376428e-08, 6.415822e-08, 6.402449e-08, 6.436151e-08, 6.43539e-08, 
    6.472909e-08, 6.455993e-08, 6.519053e-08, 6.50113e-08, 6.552921e-08, 
    6.539896e-08, 6.55231e-08, 6.548546e-08, 6.552359e-08, 6.533256e-08, 
    6.541441e-08, 6.524632e-08, 6.459161e-08, 6.478403e-08, 6.421014e-08, 
    6.386507e-08, 6.363586e-08, 6.347321e-08, 6.34962e-08, 6.354004e-08, 
    6.37653e-08, 6.397708e-08, 6.413847e-08, 6.424643e-08, 6.43528e-08, 
    6.46748e-08, 6.484521e-08, 6.522678e-08, 6.515791e-08, 6.527457e-08, 
    6.538601e-08, 6.557312e-08, 6.554232e-08, 6.562475e-08, 6.527149e-08, 
    6.550627e-08, 6.511868e-08, 6.522469e-08, 6.438174e-08, 6.406056e-08, 
    6.392407e-08, 6.380458e-08, 6.351388e-08, 6.371463e-08, 6.36355e-08, 
    6.382376e-08, 6.394339e-08, 6.388422e-08, 6.424938e-08, 6.410742e-08, 
    6.485531e-08, 6.453317e-08, 6.537302e-08, 6.517205e-08, 6.542118e-08, 
    6.529405e-08, 6.551188e-08, 6.531584e-08, 6.565543e-08, 6.572938e-08, 
    6.567885e-08, 6.587296e-08, 6.530497e-08, 6.55231e-08, 6.388257e-08, 
    6.389222e-08, 6.393717e-08, 6.373956e-08, 6.372747e-08, 6.354637e-08, 
    6.370751e-08, 6.377613e-08, 6.395032e-08, 6.405336e-08, 6.415131e-08, 
    6.436666e-08, 6.460716e-08, 6.494347e-08, 6.518507e-08, 6.534702e-08, 
    6.524771e-08, 6.533539e-08, 6.523738e-08, 6.519144e-08, 6.570168e-08, 
    6.541517e-08, 6.584504e-08, 6.582125e-08, 6.562671e-08, 6.582393e-08, 
    6.389899e-08, 6.384346e-08, 6.365067e-08, 6.380154e-08, 6.352665e-08, 
    6.368052e-08, 6.376901e-08, 6.411039e-08, 6.418539e-08, 6.425494e-08, 
    6.43923e-08, 6.456858e-08, 6.487782e-08, 6.514688e-08, 6.539249e-08, 
    6.537449e-08, 6.538083e-08, 6.54357e-08, 6.529979e-08, 6.545802e-08, 
    6.548457e-08, 6.541514e-08, 6.581807e-08, 6.570296e-08, 6.582075e-08, 
    6.574579e-08, 6.386151e-08, 6.395495e-08, 6.390446e-08, 6.39994e-08, 
    6.393252e-08, 6.422994e-08, 6.431911e-08, 6.473636e-08, 6.456511e-08, 
    6.483764e-08, 6.45928e-08, 6.463618e-08, 6.484655e-08, 6.460603e-08, 
    6.513206e-08, 6.477543e-08, 6.543784e-08, 6.508173e-08, 6.546015e-08, 
    6.539143e-08, 6.55052e-08, 6.560711e-08, 6.573531e-08, 6.597185e-08, 
    6.591708e-08, 6.611489e-08, 6.409424e-08, 6.421543e-08, 6.420476e-08, 
    6.433159e-08, 6.442539e-08, 6.462868e-08, 6.495473e-08, 6.483211e-08, 
    6.505721e-08, 6.51024e-08, 6.476043e-08, 6.497039e-08, 6.429654e-08, 
    6.440542e-08, 6.434059e-08, 6.41038e-08, 6.486038e-08, 6.447211e-08, 
    6.518906e-08, 6.497873e-08, 6.559258e-08, 6.528731e-08, 6.588692e-08, 
    6.614327e-08, 6.638449e-08, 6.666644e-08, 6.428157e-08, 6.419923e-08, 
    6.434667e-08, 6.455067e-08, 6.473994e-08, 6.499156e-08, 6.50173e-08, 
    6.506445e-08, 6.518654e-08, 6.528921e-08, 6.507936e-08, 6.531494e-08, 
    6.443068e-08, 6.489408e-08, 6.41681e-08, 6.438672e-08, 6.453865e-08, 
    6.447199e-08, 6.48181e-08, 6.489968e-08, 6.523117e-08, 6.505981e-08, 
    6.608001e-08, 6.562864e-08, 6.688109e-08, 6.653109e-08, 6.417046e-08, 
    6.428129e-08, 6.466703e-08, 6.448349e-08, 6.500836e-08, 6.513755e-08, 
    6.524257e-08, 6.537682e-08, 6.539132e-08, 6.547086e-08, 6.534052e-08, 
    6.546571e-08, 6.49921e-08, 6.520374e-08, 6.462293e-08, 6.47643e-08, 
    6.469926e-08, 6.462793e-08, 6.484809e-08, 6.508266e-08, 6.508766e-08, 
    6.516288e-08, 6.537484e-08, 6.501048e-08, 6.613828e-08, 6.54418e-08, 
    6.440214e-08, 6.461564e-08, 6.464612e-08, 6.456342e-08, 6.51246e-08, 
    6.492127e-08, 6.546892e-08, 6.532091e-08, 6.556343e-08, 6.544292e-08, 
    6.542518e-08, 6.527041e-08, 6.517404e-08, 6.493059e-08, 6.47325e-08, 
    6.457542e-08, 6.461194e-08, 6.478449e-08, 6.509701e-08, 6.539263e-08, 
    6.532787e-08, 6.5545e-08, 6.49703e-08, 6.521128e-08, 6.511815e-08, 
    6.5361e-08, 6.482886e-08, 6.528204e-08, 6.471303e-08, 6.476292e-08, 
    6.491723e-08, 6.522764e-08, 6.52963e-08, 6.536963e-08, 6.532438e-08, 
    6.510494e-08, 6.506898e-08, 6.491348e-08, 6.487055e-08, 6.475205e-08, 
    6.465395e-08, 6.474359e-08, 6.483771e-08, 6.510503e-08, 6.534592e-08, 
    6.560856e-08, 6.567284e-08, 6.597972e-08, 6.572991e-08, 6.614216e-08, 
    6.579169e-08, 6.639835e-08, 6.530828e-08, 6.578136e-08, 6.492425e-08, 
    6.501659e-08, 6.518361e-08, 6.556667e-08, 6.535986e-08, 6.560172e-08, 
    6.506757e-08, 6.479046e-08, 6.471874e-08, 6.458497e-08, 6.47218e-08, 
    6.471067e-08, 6.484161e-08, 6.479953e-08, 6.51139e-08, 6.494503e-08, 
    6.542474e-08, 6.55998e-08, 6.609416e-08, 6.639722e-08, 6.67057e-08, 
    6.684189e-08, 6.688335e-08, 6.690068e-08 ;

 SOILICE =
  56.54166, 56.73485, 56.69727, 56.85336, 56.76675, 56.86901, 56.58081, 
    56.7425, 56.63926, 56.55907, 57.1572, 56.86034, 57.46719, 57.27683, 
    57.75607, 57.43749, 57.82048, 57.74693, 57.96872, 57.90511, 58.18938, 
    57.99809, 58.33728, 58.14369, 58.17392, 57.99178, 56.92005, 57.12015, 
    56.90819, 56.93669, 56.92392, 56.76852, 56.69029, 56.52696, 56.5566, 
    56.6766, 56.94951, 56.85679, 57.09084, 57.08554, 57.34695, 57.22897, 
    57.66984, 57.54427, 57.90777, 57.81617, 57.90345, 57.87698, 57.9038, 
    57.76951, 57.82701, 57.70898, 57.25104, 57.3853, 56.98558, 56.74623, 
    56.58788, 56.47569, 56.49154, 56.52175, 56.6773, 56.82393, 56.93586, 
    57.01083, 57.08478, 57.30892, 57.428, 57.69522, 57.64698, 57.72877, 
    57.80707, 57.93864, 57.91698, 57.97499, 57.72665, 57.89158, 57.6195, 
    57.69381, 57.10466, 56.88181, 56.78709, 56.70448, 56.50372, 56.64228, 
    56.58762, 56.71779, 56.80059, 56.75964, 57.01288, 56.91431, 57.43506, 
    57.21029, 57.79793, 57.65688, 57.83179, 57.7425, 57.89554, 57.75779, 
    57.99661, 58.04869, 58.01309, 58.15001, 57.75016, 57.90343, 56.75848, 
    56.76515, 56.7963, 56.65951, 56.65116, 56.52614, 56.6374, 56.68481, 
    56.80541, 56.8768, 56.94476, 57.09439, 57.26185, 57.49675, 57.66602, 
    57.77969, 57.70998, 57.77152, 57.70272, 57.67051, 58.02916, 57.82753, 
    58.1303, 58.11353, 57.97636, 58.11541, 56.76985, 56.73143, 56.59812, 
    56.70242, 56.51254, 56.61873, 56.67985, 56.91631, 56.96843, 57.01672, 
    57.11225, 57.235, 57.45084, 57.63921, 57.81164, 57.79899, 57.80344, 
    57.84199, 57.74651, 57.85768, 57.87633, 57.82754, 58.11127, 58.03011, 
    58.11317, 58.06031, 56.74392, 56.8086, 56.77364, 56.83939, 56.79304, 
    56.99929, 57.06125, 57.35196, 57.23257, 57.42275, 57.25188, 57.28212, 
    57.42886, 57.26112, 57.62877, 57.37922, 57.84349, 57.59345, 57.85918, 
    57.81089, 57.89088, 57.96257, 58.05291, 58.2198, 58.18113, 58.32096, 
    56.90517, 56.98925, 56.98189, 57.07001, 57.13525, 57.27691, 57.50465, 
    57.41894, 57.57642, 57.60806, 57.36887, 57.51559, 57.04562, 57.12129, 
    57.07626, 56.91177, 57.43862, 57.16772, 57.66881, 57.52146, 57.95234, 
    57.73769, 58.15984, 58.34093, 58.51197, 58.7121, 57.03523, 56.97805, 
    57.08052, 57.22245, 57.35453, 57.53043, 57.54848, 57.58147, 57.66707, 
    57.73909, 57.59187, 57.75716, 57.13877, 57.46221, 56.9564, 57.10826, 
    57.2141, 57.1677, 57.40916, 57.46618, 57.69831, 57.57825, 58.29616, 
    57.97766, 58.86497, 58.61593, 56.95807, 57.03506, 57.30362, 57.17572, 
    57.54221, 57.63269, 57.70637, 57.80059, 57.8108, 57.8667, 57.77512, 
    57.8631, 57.53081, 57.67912, 57.27292, 57.37155, 57.32617, 57.2764, 
    57.43012, 57.59417, 57.59775, 57.65043, 57.79894, 57.5437, 58.33723, 
    57.84604, 57.11911, 57.26773, 57.28907, 57.23143, 57.62362, 57.48125, 
    57.86535, 57.76135, 57.93184, 57.84706, 57.8346, 57.7259, 57.65829, 
    57.48776, 57.34933, 57.23979, 57.26525, 57.38564, 57.60424, 57.8117, 
    57.76619, 57.91887, 57.51558, 57.68438, 57.61906, 57.7895, 57.41665, 
    57.73381, 57.33578, 57.37061, 57.47843, 57.69579, 57.74407, 57.79553, 
    57.76379, 57.60981, 57.58464, 57.47583, 57.44577, 57.36303, 57.29456, 
    57.35709, 57.42281, 57.6099, 57.77888, 57.96358, 58.00888, 58.22523, 
    58.04897, 58.33997, 58.09235, 58.52158, 57.75234, 58.08522, 57.48336, 
    57.54798, 57.66493, 57.93401, 57.7887, 57.95871, 57.58366, 57.38976, 
    57.33976, 57.24643, 57.3419, 57.33413, 57.42559, 57.39619, 57.61612, 
    57.49791, 57.83427, 57.95738, 58.30627, 58.52091, 58.74014, 58.83709, 
    58.86662, 58.87897,
  78.1883, 78.48907, 78.43057, 78.67358, 78.53878, 78.69795, 78.24929, 
    78.50095, 78.34027, 78.21546, 79.13866, 78.68446, 79.60855, 79.32022, 
    80.04643, 79.5635, 80.14414, 80.03271, 80.36906, 80.2726, 80.70355, 
    80.41361, 80.92805, 80.63436, 80.68015, 80.40402, 78.77749, 79.08253, 
    78.75902, 78.80337, 78.78351, 78.54149, 78.41962, 78.16549, 78.21162, 
    78.39836, 78.82333, 78.679, 79.03854, 79.03053, 79.42648, 79.24775, 
    79.91583, 79.72555, 80.27662, 80.13771, 80.27006, 80.22993, 80.27058, 
    80.06694, 80.15412, 79.97519, 79.28115, 79.48454, 78.87906, 78.50666, 
    78.26028, 78.08567, 78.11033, 78.15733, 78.39945, 78.62782, 78.80215, 
    78.91736, 79.02937, 79.36861, 79.54916, 79.95424, 79.88122, 80.00512, 
    80.12391, 80.3234, 80.29057, 80.37852, 80.00199, 80.252, 79.83959, 
    79.95219, 79.05906, 78.71795, 78.57031, 78.44179, 78.12929, 78.34495, 
    78.25986, 78.46255, 78.59148, 78.52773, 78.92046, 78.76856, 79.55987, 
    79.21938, 80.11005, 79.89622, 80.1614, 80.02603, 80.25803, 80.04921, 
    80.41133, 80.49026, 80.4363, 80.64402, 80.03763, 80.26997, 78.5259, 
    78.53629, 78.58479, 78.37176, 78.35878, 78.16419, 78.33738, 78.41117, 
    78.59901, 78.71015, 78.81598, 79.04388, 79.29748, 79.65341, 79.91006, 
    80.08242, 79.97675, 80.07003, 79.96572, 79.91691, 80.46062, 80.15489, 
    80.61412, 80.58868, 80.38058, 80.59155, 78.5436, 78.4838, 78.27622, 
    78.43863, 78.14303, 78.3083, 78.4034, 78.77161, 78.85287, 78.92624, 
    79.07095, 79.25688, 79.58387, 79.86938, 80.13086, 80.11169, 80.11843, 
    80.17685, 80.0321, 80.20064, 80.22888, 80.15495, 80.58527, 80.46215, 
    80.58813, 80.50798, 78.50325, 78.60395, 78.54951, 78.65187, 78.5797, 
    78.89976, 78.99357, 79.43396, 79.25317, 79.54127, 79.28246, 79.32822, 
    79.55035, 79.29649, 79.85346, 79.47521, 80.17912, 79.79984, 80.20292, 
    80.12972, 80.25102, 80.3597, 80.49673, 80.74982, 80.69119, 80.90334, 
    78.75433, 78.8846, 78.87354, 79.00699, 79.10577, 79.3204, 79.66545, 
    79.5356, 79.77428, 79.82221, 79.45974, 79.68199, 78.96998, 79.08451, 
    79.01641, 78.76458, 79.5653, 79.15485, 79.91427, 79.69094, 80.34417, 
    80.01862, 80.6589, 80.93346, 81.19324, 81.49686, 78.95428, 78.86772, 
    79.02291, 79.23776, 79.43797, 79.70452, 79.73192, 79.78191, 79.91169, 
    80.02087, 79.79758, 80.04826, 79.1108, 79.60107, 78.83409, 79.06476, 
    79.22515, 79.15491, 79.52081, 79.60719, 79.95896, 79.77705, 80.8655, 
    80.38246, 81.72913, 81.35091, 78.83673, 78.95406, 79.36076, 79.16707, 
    79.72242, 79.85954, 79.97128, 80.11404, 80.12959, 80.2143, 80.07549, 
    80.20887, 79.70509, 79.92992, 79.31437, 79.46375, 79.39505, 79.31964, 
    79.55255, 79.80105, 79.8066, 79.88638, 80.11111, 79.72469, 80.92757, 
    80.18259, 79.08136, 79.30632, 79.33879, 79.2515, 79.84577, 79.63, 
    80.21227, 80.05462, 80.31312, 80.18456, 80.16565, 80.00086, 79.89834, 
    79.63984, 79.43008, 79.26418, 79.30275, 79.48508, 79.81632, 80.13088, 
    80.06186, 80.29346, 79.68204, 79.93784, 79.83881, 80.09726, 79.5321, 
    80.01244, 79.40961, 79.46236, 79.62572, 79.95505, 80.02841, 80.10638, 
    80.0583, 79.82479, 79.78669, 79.62181, 79.57622, 79.4509, 79.34715, 
    79.44188, 79.5414, 79.82498, 80.08112, 80.36121, 80.42996, 80.75784, 
    80.49053, 80.93169, 80.55602, 81.20747, 80.0407, 80.54545, 79.63325, 
    79.73117, 79.90829, 80.31624, 80.09605, 80.35373, 79.78522, 79.49126, 
    79.41563, 79.27422, 79.41887, 79.4071, 79.54569, 79.50115, 79.83442, 
    79.65527, 80.16512, 80.35175, 80.881, 81.20667, 81.53962, 81.68682, 
    81.73169, 81.75044,
  118.5267, 119.0832, 118.9749, 119.4248, 119.1751, 119.4699, 118.6394, 
    119.1053, 118.8077, 118.5768, 120.3015, 119.4449, 121.1961, 120.6463, 
    122.0309, 121.1104, 122.2134, 122.0043, 122.628, 122.45, 123.2462, 
    122.7102, 123.6604, 123.118, 123.2028, 122.6926, 119.617, 120.1946, 
    119.5828, 119.665, 119.6281, 119.1802, 118.955, 118.4843, 118.5696, 
    118.9154, 119.702, 119.4346, 120.1095, 120.0942, 120.8487, 120.5081, 
    121.7815, 121.4186, 122.4574, 122.2012, 122.4454, 122.3713, 122.4464, 
    122.0696, 122.2315, 121.8946, 120.5719, 120.9595, 119.806, 119.1162, 
    118.6598, 118.3366, 118.3823, 118.4693, 118.9174, 119.3399, 119.6625, 
    119.8787, 120.092, 120.7393, 121.0829, 121.8549, 121.7154, 121.9519, 
    122.1757, 122.5439, 122.4832, 122.6456, 121.9457, 122.4122, 121.6359, 
    121.8508, 120.15, 119.5067, 119.234, 118.9957, 118.4174, 118.8165, 
    118.6591, 119.034, 119.2726, 119.1545, 119.8846, 119.6004, 121.1033, 
    120.4543, 122.1502, 121.744, 122.2449, 121.9915, 122.4233, 122.0357, 
    122.7061, 122.852, 122.7523, 123.1356, 122.0136, 122.4454, 119.1512, 
    119.1705, 119.2602, 118.8662, 118.8421, 118.4819, 118.8024, 118.939, 
    119.2865, 119.4923, 119.6882, 120.1198, 120.6031, 121.2814, 121.7704, 
    122.099, 121.8975, 122.0754, 121.8765, 121.7833, 122.7973, 122.233, 
    123.0805, 123.0335, 122.6495, 123.0387, 119.184, 119.0732, 118.6893, 
    118.9897, 118.4428, 118.7487, 118.9248, 119.6063, 119.7565, 119.8958, 
    120.1713, 120.5255, 121.1488, 121.693, 122.1885, 122.1531, 122.1655, 
    122.2734, 122.0031, 122.3173, 122.3695, 122.233, 123.0272, 122.7999, 
    123.0325, 122.8844, 119.1092, 119.2957, 119.1949, 119.3845, 119.2509, 
    119.8456, 120.0244, 120.8634, 120.5186, 121.0677, 120.5743, 120.6616, 
    121.0856, 120.6009, 121.6629, 120.9421, 122.2776, 121.561, 122.3215, 
    122.1864, 122.4102, 122.6109, 122.8637, 123.3312, 123.2229, 123.6146, 
    119.5741, 119.8166, 119.7953, 120.0495, 120.2377, 120.6465, 121.3042, 
    121.0566, 121.5115, 121.6029, 120.9119, 121.3358, 119.9792, 120.1976, 
    120.0675, 119.5932, 121.1136, 120.3315, 121.7785, 121.3527, 122.5822, 
    121.9777, 123.1632, 123.6708, 124.1501, 124.7117, 119.9492, 119.7842, 
    120.0797, 120.4895, 120.8706, 121.3787, 121.4307, 121.5261, 121.7734, 
    121.9816, 121.5563, 122.0339, 120.2482, 121.1816, 119.7218, 120.16, 
    120.4653, 120.3313, 121.0283, 121.193, 121.8639, 121.5167, 123.5454, 
    122.6532, 125.1407, 124.4418, 119.7266, 119.9486, 120.7237, 120.3544, 
    121.4126, 121.6741, 121.887, 122.1576, 122.1861, 122.3426, 122.0858, 
    122.3325, 121.3797, 121.8083, 120.6349, 120.9197, 120.7887, 120.645, 
    121.0888, 121.5629, 121.5731, 121.7254, 122.1535, 121.4169, 123.6608, 
    122.2852, 120.1911, 120.6202, 120.6816, 120.5152, 121.6479, 121.2366, 
    122.3388, 122.046, 122.5248, 122.2876, 122.2527, 121.9435, 121.7481, 
    121.2554, 120.8556, 120.5393, 120.6128, 120.9605, 121.592, 122.1887, 
    122.0601, 122.4885, 121.3357, 121.8235, 121.6348, 122.1266, 121.05, 
    121.9669, 120.8164, 120.917, 121.2284, 121.8567, 121.996, 122.1435, 
    122.053, 121.6081, 121.5353, 121.2208, 121.1341, 120.8951, 120.6974, 
    120.878, 121.0678, 121.6083, 122.0968, 122.6137, 122.7405, 123.3467, 
    122.853, 123.6685, 122.9748, 124.1774, 122.0203, 122.9545, 121.2426, 
    121.4293, 121.7674, 122.5311, 122.1243, 122.6002, 121.5324, 120.9725, 
    120.8279, 120.5585, 120.8341, 120.8116, 121.0757, 120.9908, 121.6262, 
    121.2846, 122.2518, 122.5964, 123.5735, 124.1753, 124.7902, 125.0623, 
    125.1452, 125.1799,
  187.3257, 188.3278, 188.1326, 188.9433, 188.4933, 189.0246, 187.5285, 
    188.3677, 187.8316, 187.4157, 190.5242, 188.9795, 192.1386, 191.146, 
    193.6468, 191.9839, 193.9758, 193.5986, 194.7247, 194.4031, 195.8423, 
    194.8732, 196.5915, 195.6105, 195.7637, 194.8413, 189.2895, 190.3314, 
    189.228, 189.3762, 189.3096, 188.5026, 188.0969, 187.2492, 187.4029, 
    188.0256, 189.4429, 188.9608, 190.1774, 190.1499, 191.5113, 190.8966, 
    193.1959, 192.5402, 194.4165, 193.9536, 194.3947, 194.2609, 194.3965, 
    193.7167, 194.0085, 193.4003, 191.0116, 191.7113, 189.6303, 188.3875, 
    187.5653, 186.9835, 187.0657, 187.2224, 188.0292, 188.7901, 189.3716, 
    189.7613, 190.146, 191.314, 191.9342, 193.3287, 193.0764, 193.5039, 
    193.9077, 194.5727, 194.4631, 194.7566, 193.4926, 194.3349, 192.9328, 
    193.321, 190.2509, 189.0908, 188.5995, 188.1702, 187.1289, 187.8475, 
    187.564, 188.239, 188.6689, 188.4562, 189.772, 189.2596, 191.971, 
    190.7995, 193.8615, 193.1282, 194.0325, 193.5753, 194.3549, 193.6553, 
    194.8658, 195.1295, 194.9493, 195.6422, 193.6154, 194.3948, 188.4502, 
    188.4849, 188.6465, 187.9369, 187.8935, 187.245, 187.822, 188.0681, 
    188.6938, 189.0648, 189.4179, 190.1961, 191.0681, 192.2926, 193.1759, 
    193.7693, 193.4054, 193.727, 193.3675, 193.1992, 195.0307, 194.0112, 
    195.5424, 195.4574, 194.7635, 195.467, 188.5093, 188.3097, 187.6183, 
    188.1592, 187.1745, 187.7253, 188.0425, 189.2704, 189.5409, 189.7921, 
    190.2889, 190.928, 192.0531, 193.0361, 193.9306, 193.8668, 193.8893, 
    194.0841, 193.5964, 194.1634, 194.2578, 194.0111, 195.446, 195.0352, 
    195.4556, 195.188, 188.3746, 188.7105, 188.5289, 188.8705, 188.6298, 
    189.7018, 190.0241, 191.5378, 190.9154, 191.9066, 191.0159, 191.1735, 
    191.9391, 191.0639, 192.9818, 191.6801, 194.0917, 192.7978, 194.171, 
    193.9269, 194.3311, 194.6937, 195.1506, 195.996, 195.7999, 196.5085, 
    189.2121, 189.6494, 189.6108, 190.0692, 190.4088, 191.1462, 192.3336, 
    191.8864, 192.708, 192.8732, 191.6253, 192.3909, 189.9425, 190.3365, 
    190.1018, 189.2466, 191.9895, 190.5781, 193.1905, 192.4213, 194.642, 
    193.5506, 195.6921, 196.6104, 197.4775, 198.4949, 189.8884, 189.5909, 
    190.1237, 190.863, 191.5508, 192.4681, 192.5621, 192.7345, 193.1813, 
    193.5576, 192.789, 193.652, 190.4281, 192.1124, 189.4785, 190.2688, 
    190.8194, 190.5776, 191.8354, 192.1327, 193.3448, 192.7175, 196.3835, 
    194.7704, 199.2722, 198.006, 189.487, 189.8873, 191.2856, 190.6193, 
    192.5294, 193.0019, 193.3866, 193.8751, 193.9265, 194.209, 193.7458, 
    194.1907, 192.4701, 193.2443, 191.1253, 191.6395, 191.4028, 191.1435, 
    191.9447, 192.8011, 192.8194, 193.0946, 193.8682, 192.5372, 196.5926, 
    194.1059, 190.3246, 191.0989, 191.2096, 190.9093, 192.9545, 192.2115, 
    194.2021, 193.6739, 194.5382, 194.1097, 194.0468, 193.4886, 193.1355, 
    192.2455, 191.5237, 190.9528, 191.0854, 191.713, 192.8536, 193.9312, 
    193.6995, 194.4726, 192.3905, 193.2719, 192.9309, 193.8189, 191.8746, 
    193.5314, 191.4529, 191.6344, 192.1968, 193.3319, 193.5836, 193.8495, 
    193.6866, 192.8826, 192.7511, 192.1831, 192.0265, 191.5949, 191.2381, 
    191.5641, 191.9069, 192.8829, 193.7654, 194.6989, 194.9278, 196.0242, 
    195.1315, 196.6065, 195.3521, 197.5275, 193.6276, 195.3151, 192.2224, 
    192.5595, 193.1706, 194.5498, 193.8148, 194.6745, 192.7459, 191.7347, 
    191.4736, 190.9875, 191.4848, 191.4443, 191.921, 191.7677, 192.9153, 
    192.2982, 194.0452, 194.6677, 196.4342, 197.5234, 198.6369, 199.1301, 
    199.2803, 199.3432,
  314.8267, 316.5648, 316.2261, 317.6333, 316.8519, 317.7744, 315.1783, 
    316.634, 315.7039, 314.9827, 320.3815, 317.6962, 323.1932, 321.4637, 
    325.825, 322.9236, 326.413, 325.7408, 327.7677, 327.1858, 329.7831, 
    328.0367, 331.0962, 329.372, 329.6455, 327.9789, 318.2347, 320.0461, 
    318.1277, 318.3853, 318.2697, 316.8681, 316.1642, 314.6942, 314.9605, 
    316.0403, 318.5012, 317.6637, 319.7782, 319.7303, 322.1, 321.0295, 
    325.0375, 323.8935, 327.2101, 326.3729, 327.1707, 326.9286, 327.1739, 
    325.947, 326.4721, 325.3944, 321.2297, 322.4484, 318.8269, 316.6684, 
    315.242, 314.2337, 314.3761, 314.6477, 316.0467, 317.3673, 318.3773, 
    319.0547, 319.7234, 321.7563, 322.8369, 325.2694, 324.829, 325.5754, 
    326.2897, 327.4927, 327.2944, 327.8255, 325.5555, 327.0625, 324.5784, 
    325.256, 319.906, 317.8894, 317.0365, 316.2912, 314.4856, 315.7315, 
    315.2398, 316.4107, 317.1569, 316.7876, 319.0732, 318.1828, 322.9011, 
    320.8605, 326.2063, 324.9193, 326.5155, 325.7001, 327.0986, 325.8397, 
    328.0233, 328.5007, 328.1744, 329.4294, 325.77, 327.1708, 316.7773, 
    316.8375, 317.118, 315.8865, 315.8113, 314.6869, 315.6872, 316.1141, 
    317.2002, 317.8443, 318.4578, 319.8107, 321.3282, 323.4616, 325.0026, 
    326.0396, 325.4033, 325.965, 325.3372, 325.0433, 328.3218, 326.477, 
    329.2487, 329.0947, 327.8382, 329.112, 316.8798, 316.5334, 315.334, 
    316.2723, 314.5646, 315.5195, 316.0698, 318.2015, 318.6715, 319.1082, 
    319.9721, 321.0842, 323.0441, 324.7586, 326.3313, 326.2158, 326.2565, 
    326.6088, 325.7368, 326.7522, 326.9229, 326.4767, 329.074, 328.33, 
    329.0914, 328.6067, 316.6459, 317.2291, 316.9138, 317.5069, 317.089, 
    318.9513, 319.5116, 322.1462, 321.0623, 322.7888, 321.2372, 321.5117, 
    322.8455, 321.3208, 324.6639, 322.394, 326.6225, 324.3428, 326.7659, 
    326.3245, 327.0556, 327.7117, 328.5389, 330.0524, 329.7089, 330.9507, 
    318.1002, 318.8602, 318.7931, 319.59, 320.1805, 321.4641, 323.5332, 
    322.7536, 324.1861, 324.4745, 322.2986, 323.633, 319.3696, 320.0549, 
    319.6466, 318.1602, 322.9332, 320.4752, 325.0282, 323.686, 327.6181, 
    325.657, 329.5199, 331.1294, 332.6507, 334.4381, 319.2755, 318.7583, 
    319.6848, 320.9711, 322.1687, 323.7677, 323.9317, 324.2323, 325.012, 
    325.669, 324.3275, 325.8339, 320.2142, 323.1474, 318.5631, 319.9371, 
    320.8951, 320.4744, 322.6646, 323.1829, 325.2975, 324.2027, 330.7316, 
    327.8507, 335.8051, 333.5789, 318.5779, 319.2737, 321.7069, 320.5469, 
    323.8747, 324.6989, 325.3704, 326.2309, 326.3238, 326.8348, 325.9979, 
    326.8016, 323.7711, 325.122, 321.4277, 322.3232, 321.9109, 321.4594, 
    322.855, 324.3486, 324.3804, 324.8608, 326.2186, 323.8882, 331.0983, 
    326.6484, 320.0341, 321.3818, 321.5745, 321.0515, 324.6162, 323.3203, 
    326.8223, 325.8722, 327.4303, 326.6552, 326.5413, 325.5486, 324.9321, 
    323.3796, 322.1216, 321.1273, 321.3582, 322.4514, 324.4402, 326.3323, 
    325.9169, 327.3116, 323.6323, 325.1703, 324.5751, 326.1293, 322.7329, 
    325.6235, 321.9981, 322.3144, 323.2946, 325.275, 325.7144, 326.1847, 
    325.8944, 324.4908, 324.2613, 323.2707, 322.9978, 322.2455, 321.6241, 
    322.1918, 322.7892, 324.4913, 326.0326, 327.7211, 328.1355, 330.1019, 
    328.5043, 331.1227, 328.904, 332.7387, 325.7915, 328.8369, 323.3392, 
    323.9271, 324.9934, 327.4513, 326.1219, 327.6771, 324.2523, 322.4892, 
    322.0344, 321.1877, 322.0537, 321.9832, 322.8138, 322.5467, 324.5479, 
    323.4715, 326.5385, 327.6647, 330.8204, 332.7313, 334.6876, 335.555, 
    335.8195, 335.9301,
  523.2241, 526.4968, 525.8586, 528.5126, 527.0382, 528.7791, 523.8855, 
    526.6274, 524.8749, 523.5175, 533.7101, 528.6313, 539.0477, 535.7621, 
    544.0626, 538.535, 545.1855, 543.9017, 547.7762, 546.6627, 551.6569, 
    548.2911, 554.2677, 550.8506, 551.3835, 548.1806, 529.6483, 533.0747, 
    529.4462, 529.9329, 529.7144, 527.0687, 525.7418, 522.9748, 523.4758, 
    525.5085, 530.152, 528.5699, 532.5674, 532.4767, 536.97, 534.9384, 
    542.5602, 540.3803, 546.7092, 545.1089, 546.6339, 546.1709, 546.64, 
    544.2954, 545.2984, 543.2408, 535.3182, 537.6318, 530.7676, 526.6922, 
    524.0054, 522.1091, 522.3767, 522.8873, 525.5204, 528.0105, 529.9178, 
    531.1983, 532.4637, 536.3174, 538.3702, 543.0025, 542.1626, 543.5862, 
    544.9501, 547.2499, 546.8705, 547.8868, 543.5483, 546.427, 541.6849, 
    542.9769, 532.8095, 528.9961, 527.3863, 525.9812, 522.5826, 524.9268, 
    524.0012, 526.2063, 527.6135, 526.9169, 531.2334, 529.5502, 538.4922, 
    534.618, 544.7908, 542.3348, 545.3814, 543.8241, 546.496, 544.0906, 
    548.2656, 549.1801, 548.5549, 550.9608, 543.9576, 546.634, 526.8975, 
    527.011, 527.5402, 525.2188, 525.0771, 522.9611, 524.8434, 525.6475, 
    527.6951, 528.9109, 530.0699, 532.6289, 535.5049, 539.5583, 542.4936, 
    544.4723, 543.2579, 544.3299, 543.1317, 542.5712, 548.8373, 545.3079, 
    550.614, 550.3186, 547.9111, 550.3519, 527.0907, 526.4377, 524.1785, 
    525.9455, 522.7313, 524.5276, 525.564, 529.5856, 530.4739, 531.2995, 
    532.9346, 535.0421, 538.7641, 542.0284, 545.0295, 544.8088, 544.8865, 
    545.5597, 543.8943, 545.8337, 546.1602, 545.3073, 550.2791, 548.8529, 
    550.3123, 549.3831, 526.6498, 527.7496, 527.155, 528.2739, 527.4854, 
    531.0027, 532.0629, 537.0577, 535.0006, 538.2787, 535.3324, 535.8531, 
    538.3866, 535.491, 541.848, 537.5285, 545.5859, 541.2361, 545.8599, 
    545.0165, 546.4137, 547.6691, 549.2532, 552.1918, 551.5095, 553.9781, 
    529.3943, 530.8304, 530.7036, 532.2111, 533.3294, 535.7628, 539.6946, 
    538.2119, 540.9376, 541.4869, 537.3472, 539.8845, 531.7941, 533.0914, 
    532.3184, 529.5075, 538.5534, 533.8877, 542.5423, 539.9854, 547.4899, 
    543.7419, 551.1345, 554.3337, 557.2768, 560.7276, 531.6161, 530.6379, 
    532.3906, 534.8277, 537.1005, 540.1409, 540.4531, 541.0255, 542.5115, 
    543.7649, 541.2069, 544.0797, 533.3932, 538.9606, 530.2689, 532.8683, 
    534.6836, 533.8861, 538.0427, 539.0281, 543.056, 540.9691, 553.5422, 
    547.935, 563.3732, 559.0676, 530.2968, 531.6126, 536.2236, 534.0236, 
    540.3445, 541.9147, 543.195, 544.8376, 545.0151, 545.9916, 544.3926, 
    545.9282, 540.1475, 542.7213, 535.6938, 537.394, 536.611, 535.7538, 
    538.4047, 541.2471, 541.3077, 542.2232, 544.8141, 540.3704, 554.2719, 
    545.6353, 533.052, 535.6067, 535.9724, 534.9802, 541.757, 539.2894, 
    545.9677, 544.1526, 547.1304, 545.6483, 545.4306, 543.5351, 542.3592, 
    539.4023, 537.011, 535.1239, 535.562, 537.6375, 541.4215, 545.0314, 
    544.2381, 546.9034, 539.8832, 542.8134, 541.6786, 544.6436, 538.1726, 
    543.678, 536.7766, 537.3773, 539.2405, 543.0131, 543.8516, 544.7493, 
    544.1951, 541.5179, 541.0807, 539.1951, 538.6761, 537.2463, 536.0663, 
    537.1445, 538.2795, 541.5189, 544.459, 547.687, 548.4805, 552.2903, 
    549.187, 554.3205, 549.953, 557.4465, 543.9987, 549.8245, 539.3254, 
    540.4444, 542.476, 547.1707, 544.6296, 547.6027, 541.0635, 537.7094, 
    536.8453, 535.2385, 536.8821, 536.7482, 538.3264, 537.8186, 541.6268, 
    539.5771, 545.4252, 547.5791, 553.7189, 557.4323, 561.21, 562.8888, 
    563.401, 563.6154,
  947.1252, 953.998, 952.6549, 958.2488, 955.1384, 958.8117, 948.5112, 
    954.2729, 950.5876, 947.7399, 969.1228, 958.4996, 980.1627, 973.3557, 
    990.624, 979.098, 992.9788, 990.2872, 998.4282, 996.0831, 1006.636, 
    999.5141, 1012.19, 1004.926, 1006.056, 999.2809, 960.6497, 967.8149, 
    960.2222, 961.2521, 960.7896, 955.2027, 952.4093, 946.603, 947.6523, 
    951.9189, 961.7158, 958.3699, 966.7717, 966.5853, 975.8538, 971.6547, 
    987.4808, 982.934, 996.1807, 992.818, 996.0224, 995.0486, 996.0351, 
    991.1119, 993.2156, 988.9039, 972.4387, 977.2248, 963.0202, 954.4094, 
    948.7628, 944.7917, 945.3513, 946.4199, 951.944, 957.1887, 961.22, 
    963.9335, 966.5585, 974.5035, 978.756, 988.4053, 986.6502, 989.6265, 
    992.4846, 997.3192, 996.5203, 998.6613, 989.5472, 995.5871, 985.6532, 
    988.3517, 967.2695, 959.2704, 955.8721, 952.9129, 945.782, 950.6966, 
    948.754, 953.3865, 956.351, 954.8827, 964.0079, 960.4421, 979.0092, 
    970.9939, 992.1504, 987.0099, 993.39, 990.1246, 995.7322, 990.6827, 
    999.4601, 1001.391, 1000.071, 1005.16, 990.4042, 996.0226, 954.8417, 
    955.0809, 956.1964, 951.31, 951.0124, 946.5743, 950.5213, 952.211, 
    956.5232, 959.0905, 961.5421, 966.8981, 972.8243, 981.2239, 987.3416, 
    991.4827, 988.9394, 991.1841, 988.6755, 987.5037, 1000.667, 993.2355, 
    1004.425, 1003.799, 998.7124, 1003.87, 955.2489, 953.8735, 949.1257, 
    952.8378, 946.0931, 949.8585, 952.0355, 960.517, 962.3976, 964.1481, 
    967.5267, 971.8688, 979.5736, 986.37, 992.6512, 992.1884, 992.3513, 
    993.7643, 990.2716, 994.3398, 995.0259, 993.2343, 1003.716, 1000.7, 
    1003.786, 1001.82, 954.3201, 956.6383, 955.3845, 957.7448, 956.0811, 
    963.5187, 965.735, 976.0355, 971.7831, 978.5663, 972.468, 973.5436, 
    978.7901, 972.7956, 985.9934, 977.0107, 993.8193, 984.717, 994.395, 
    992.6239, 995.5592, 998.2023, 1001.546, 1007.772, 1006.324, 1011.573, 
    960.1123, 963.1534, 962.8846, 966.0395, 968.339, 973.3571, 981.5072, 
    978.4274, 984.0947, 985.24, 976.6351, 981.9022, 965.1832, 967.8492, 
    966.2599, 960.3519, 979.1362, 969.4886, 987.4434, 982.1121, 997.8247, 
    989.9525, 1005.528, 1012.331, 1018.812, 1026.49, 964.8176, 962.7454, 
    966.4084, 971.4264, 976.1241, 982.4358, 983.0856, 984.2781, 987.379, 
    990.0006, 984.6562, 990.6598, 968.4703, 979.9818, 961.9636, 967.3903, 
    971.1291, 969.4853, 978.0765, 980.1221, 988.5173, 984.1605, 1010.644, 
    998.7629, 1032.29, 1022.79, 962.0225, 964.8105, 974.3096, 969.7685, 
    982.8596, 986.1326, 988.808, 992.2487, 992.6211, 994.6717, 991.3157, 
    994.5385, 982.4493, 987.8174, 973.2145, 976.732, 975.1108, 973.3385, 
    978.8276, 984.74, 984.8663, 986.7768, 992.1995, 982.9133, 1012.199, 
    993.9232, 967.7681, 973.0344, 973.79, 971.741, 985.8036, 980.6649, 
    994.6215, 990.8128, 997.0675, 993.9503, 993.4932, 989.5195, 987.0609, 
    980.8995, 975.9388, 972.0376, 972.9421, 977.2364, 985.1036, 992.6552, 
    990.9918, 996.5895, 981.8994, 988.0099, 985.6401, 991.8417, 978.346, 
    989.8188, 975.4534, 976.6972, 980.5634, 988.4275, 990.1821, 992.0635, 
    990.9017, 985.3047, 984.3931, 980.4689, 979.3909, 976.4261, 973.9844, 
    976.215, 978.5679, 985.3068, 991.4548, 998.2401, 999.9137, 1007.982, 
    1001.406, 1012.302, 1003.026, 1019.188, 990.4902, 1002.754, 980.7397, 
    983.0674, 987.3049, 997.1524, 991.8124, 998.0624, 984.3574, 977.3856, 
    975.5958, 972.2741, 975.6719, 975.3947, 978.665, 977.6119, 985.532, 
    981.2628, 993.4819, 998.0126, 1011.02, 1019.156, 1027.567, 1031.239, 
    1032.351, 1032.816,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.786, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.368, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.288, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.251, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.495, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.375, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.824, 1995.068, 1990.795, 2007.356, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.699, 1840.855, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.442, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.949, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.384, 1967.079, 1965.616, 1966.131, 
    1970.605, 1959.577, 1972.433, 1974.615, 1968.925, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.141, 1901.946, 1923.064, 1904.062, 1907.391, 
    1923.767, 1905.075, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.774, 1874.989, 1884.356, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.877, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.029, 2079.234, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.519, 1872.306, 1888.469, 
    1899.93, 1894.878, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.747, 
    1936.524, 1946.646, 1954.988, 1965.806, 1966.984, 1973.488, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.672, 
    1971.109, 1889.623, 1905.814, 1908.155, 1901.817, 1945.625, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.572, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.084, 1963.301, 1984.896, 1990.287, 2016.644, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.429, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.07, 1944.782, 
    1931.565, 1969.709, 1984.166, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.539419, 4.557943, 4.554338, 4.56931, 4.560999, 4.57081, 4.543169, 
    4.558681, 4.548774, 4.541083, 4.598465, 4.569978, 4.628177, 4.609915, 
    4.65588, 4.625333, 4.662055, 4.654995, 4.676262, 4.670163, 4.69744, 
    4.679079, 4.711618, 4.69305, 4.695952, 4.678474, 4.575699, 4.594913, 
    4.574563, 4.577299, 4.576071, 4.561172, 4.553677, 4.538004, 4.540846, 
    4.552358, 4.578529, 4.569633, 4.592074, 4.591566, 4.616639, 4.605322, 
    4.647602, 4.635558, 4.670417, 4.661634, 4.670005, 4.667465, 4.670038, 
    4.657161, 4.662675, 4.651355, 4.607441, 4.620318, 4.581986, 4.559046, 
    4.543849, 4.533088, 4.534608, 4.537508, 4.552426, 4.566481, 4.577213, 
    4.584403, 4.591493, 4.613008, 4.624419, 4.650041, 4.645408, 4.653257, 
    4.660761, 4.67338, 4.671301, 4.676867, 4.653049, 4.66887, 4.642771, 
    4.6499, 4.593429, 4.572031, 4.562963, 4.55503, 4.535778, 4.549067, 
    4.543825, 4.556302, 4.564244, 4.560315, 4.584599, 4.575148, 4.625095, 
    4.603535, 4.659885, 4.646358, 4.663131, 4.654567, 4.669249, 4.656034, 
    4.678939, 4.683938, 4.680522, 4.69365, 4.655303, 4.670005, 4.560205, 
    4.560845, 4.56383, 4.55072, 4.549918, 4.537926, 4.548595, 4.553144, 
    4.564703, 4.571552, 4.578068, 4.592418, 4.608482, 4.631007, 4.647235, 
    4.658134, 4.651448, 4.657351, 4.650753, 4.647663, 4.682065, 4.662727, 
    4.691761, 4.690151, 4.677, 4.690332, 4.561295, 4.557609, 4.544829, 
    4.554829, 4.536622, 4.546808, 4.552672, 4.575346, 4.580337, 4.58497, 
    4.594129, 4.605901, 4.626604, 4.644668, 4.661198, 4.659985, 4.660412, 
    4.66411, 4.654954, 4.665615, 4.667406, 4.662724, 4.689935, 4.68215, 
    4.690116, 4.685046, 4.558807, 4.565011, 4.561658, 4.567966, 4.563522, 
    4.583306, 4.589249, 4.617127, 4.60567, 4.623911, 4.60752, 4.610422, 
    4.62451, 4.608404, 4.643672, 4.619744, 4.664254, 4.640291, 4.665759, 
    4.661126, 4.668797, 4.675676, 4.684337, 4.700349, 4.696638, 4.710049, 
    4.574271, 4.582339, 4.581627, 4.590079, 4.596337, 4.609919, 4.631762, 
    4.623539, 4.638641, 4.641677, 4.618736, 4.632813, 4.587743, 4.595006, 
    4.59068, 4.574908, 4.625435, 4.599457, 4.647503, 4.633372, 4.674695, 
    4.654115, 4.694596, 4.711977, 4.728366, 4.747574, 4.586745, 4.581258, 
    4.591084, 4.604705, 4.617365, 4.634233, 4.635961, 4.639127, 4.647333, 
    4.654241, 4.64013, 4.655974, 4.596694, 4.627694, 4.579186, 4.593758, 
    4.603901, 4.599448, 4.6226, 4.628068, 4.650336, 4.638815, 4.707684, 
    4.677131, 4.762229, 4.738348, 4.579343, 4.586725, 4.612485, 4.600216, 
    4.635361, 4.64404, 4.651102, 4.660143, 4.661119, 4.666481, 4.657696, 
    4.666134, 4.63427, 4.64849, 4.609535, 4.618997, 4.614642, 4.609869, 
    4.62461, 4.640352, 4.640687, 4.645743, 4.660014, 4.635503, 4.711641, 
    4.664526, 4.594785, 4.609049, 4.611086, 4.605556, 4.643169, 4.629517, 
    4.66635, 4.656376, 4.672726, 4.664597, 4.663402, 4.652976, 4.646493, 
    4.630143, 4.616867, 4.606358, 4.608799, 4.620349, 4.641316, 4.661208, 
    4.656846, 4.671482, 4.632806, 4.648999, 4.642736, 4.659076, 4.623322, 
    4.653763, 4.615563, 4.618903, 4.629246, 4.6501, 4.654718, 4.659658, 
    4.656609, 4.641849, 4.639432, 4.628994, 4.626116, 4.618176, 4.61161, 
    4.617609, 4.623915, 4.641854, 4.658061, 4.675774, 4.680115, 4.700885, 
    4.683976, 4.711905, 4.688157, 4.729313, 4.655529, 4.687456, 4.629716, 
    4.635913, 4.647138, 4.672947, 4.658999, 4.675313, 4.639338, 4.620749, 
    4.615945, 4.606997, 4.61615, 4.615405, 4.624175, 4.621356, 4.64245, 
    4.631111, 4.663372, 4.675183, 4.708642, 4.729234, 4.750251, 4.75955, 
    4.762383, 4.763567,
  5.632068, 5.65533, 5.650802, 5.669606, 5.659168, 5.67149, 5.636777, 
    5.656256, 5.643815, 5.634158, 5.706233, 5.670445, 5.743571, 5.72062, 
    5.778398, 5.739996, 5.786162, 5.777284, 5.804028, 5.796357, 5.830667, 
    5.807571, 5.848504, 5.825143, 5.828794, 5.80681, 5.677631, 5.701769, 
    5.676204, 5.679641, 5.678098, 5.659384, 5.649972, 5.630291, 5.63386, 
    5.648316, 5.681187, 5.670011, 5.698202, 5.697564, 5.729069, 5.714849, 
    5.76799, 5.752849, 5.796677, 5.785633, 5.796158, 5.792965, 5.7962, 
    5.780008, 5.786942, 5.772707, 5.717511, 5.733694, 5.685529, 5.656715, 
    5.637631, 5.62412, 5.626028, 5.629669, 5.648401, 5.666053, 5.679533, 
    5.688564, 5.697473, 5.724506, 5.738847, 5.771056, 5.765232, 5.775099, 
    5.784535, 5.800404, 5.79779, 5.804789, 5.774837, 5.794732, 5.761916, 
    5.770878, 5.699905, 5.673024, 5.661634, 5.651672, 5.627496, 5.644184, 
    5.637601, 5.653269, 5.663243, 5.658308, 5.688811, 5.676939, 5.739698, 
    5.712603, 5.783433, 5.766427, 5.787515, 5.776747, 5.795208, 5.778591, 
    5.807395, 5.813682, 5.809385, 5.825899, 5.777671, 5.796159, 5.65817, 
    5.658975, 5.662724, 5.646259, 5.645252, 5.630194, 5.64359, 5.649303, 
    5.66382, 5.672422, 5.680607, 5.698635, 5.718819, 5.747128, 5.767528, 
    5.781232, 5.772825, 5.780247, 5.771951, 5.768066, 5.811326, 5.787007, 
    5.823522, 5.821496, 5.804956, 5.821725, 5.65954, 5.654911, 5.638862, 
    5.651418, 5.628556, 5.641346, 5.64871, 5.677188, 5.683457, 5.689278, 
    5.700784, 5.715576, 5.741594, 5.7643, 5.785084, 5.783559, 5.784096, 
    5.788746, 5.777233, 5.790638, 5.792891, 5.787003, 5.821225, 5.811433, 
    5.821454, 5.815076, 5.656415, 5.664207, 5.659996, 5.667917, 5.662336, 
    5.687187, 5.694653, 5.729682, 5.715285, 5.738209, 5.71761, 5.721257, 
    5.738962, 5.718721, 5.763048, 5.732972, 5.788927, 5.758799, 5.790819, 
    5.784994, 5.79464, 5.80329, 5.814184, 5.834326, 5.829658, 5.846529, 
    5.675837, 5.685972, 5.685078, 5.695695, 5.703558, 5.720624, 5.748077, 
    5.737742, 5.756724, 5.76054, 5.731705, 5.749399, 5.692761, 5.701886, 
    5.69645, 5.676637, 5.740125, 5.707479, 5.767866, 5.750101, 5.802057, 
    5.776178, 5.827089, 5.848955, 5.869579, 5.893755, 5.691507, 5.684615, 
    5.696959, 5.714073, 5.729982, 5.751184, 5.753356, 5.757336, 5.767652, 
    5.776337, 5.758596, 5.778515, 5.704007, 5.742964, 5.682012, 5.700318, 
    5.713063, 5.707468, 5.736561, 5.743434, 5.771427, 5.756943, 5.843554, 
    5.805121, 5.912204, 5.882141, 5.682208, 5.691483, 5.72385, 5.708433, 
    5.7526, 5.763511, 5.77239, 5.783757, 5.784984, 5.791728, 5.780681, 
    5.791291, 5.751229, 5.769107, 5.720141, 5.732032, 5.726559, 5.720562, 
    5.739088, 5.758875, 5.759296, 5.765652, 5.783596, 5.75278, 5.848533, 
    5.789269, 5.701609, 5.719531, 5.722091, 5.715142, 5.762417, 5.745255, 
    5.791563, 5.779021, 5.799581, 5.789358, 5.787855, 5.774745, 5.766596, 
    5.746041, 5.729356, 5.716149, 5.719218, 5.733733, 5.760087, 5.785097, 
    5.779612, 5.798016, 5.74939, 5.769745, 5.761872, 5.782416, 5.737468, 
    5.775736, 5.727717, 5.731915, 5.744915, 5.77113, 5.776937, 5.783147, 
    5.779314, 5.760756, 5.757719, 5.744598, 5.74098, 5.731, 5.722749, 
    5.730289, 5.738214, 5.760763, 5.78114, 5.803414, 5.808873, 5.835001, 
    5.813729, 5.848865, 5.818989, 5.870771, 5.777955, 5.818107, 5.745506, 
    5.753295, 5.767406, 5.799859, 5.782319, 5.802834, 5.7576, 5.734235, 
    5.728198, 5.716952, 5.728455, 5.727519, 5.738541, 5.734997, 5.761513, 
    5.747259, 5.787818, 5.802671, 5.84476, 5.870671, 5.897125, 5.908832, 
    5.912398, 5.913889,
  8.097889, 8.132088, 8.125429, 8.153082, 8.137732, 8.155853, 8.104812, 
    8.13345, 8.115157, 8.100961, 8.206968, 8.154317, 8.261936, 8.228145, 
    8.313236, 8.256673, 8.324678, 8.311596, 8.35101, 8.339704, 8.390287, 
    8.356234, 8.416598, 8.382143, 8.387527, 8.355112, 8.164887, 8.200399, 
    8.162787, 8.167843, 8.165573, 8.13805, 8.12421, 8.095278, 8.100523, 
    8.121776, 8.170116, 8.153678, 8.195151, 8.194213, 8.240583, 8.21965, 
    8.297902, 8.2756, 8.340176, 8.323898, 8.339411, 8.334704, 8.339472, 
    8.31561, 8.325827, 8.304853, 8.223568, 8.247392, 8.176505, 8.134126, 
    8.106067, 8.086206, 8.089011, 8.094362, 8.1219, 8.147858, 8.167686, 
    8.180971, 8.194078, 8.233866, 8.25498, 8.30242, 8.293839, 8.308377, 
    8.32228, 8.345668, 8.341814, 8.352133, 8.307991, 8.337308, 8.288955, 
    8.302158, 8.197658, 8.15811, 8.141358, 8.126709, 8.091169, 8.1157, 
    8.106023, 8.129058, 8.143723, 8.136467, 8.181334, 8.163868, 8.256232, 
    8.216345, 8.320658, 8.295599, 8.326672, 8.310804, 8.338009, 8.313521, 
    8.355974, 8.365242, 8.358908, 8.383257, 8.312166, 8.339412, 8.136264, 
    8.137447, 8.142961, 8.11875, 8.11727, 8.095135, 8.114827, 8.123226, 
    8.144574, 8.157225, 8.169265, 8.195787, 8.225493, 8.267175, 8.297222, 
    8.317412, 8.305026, 8.315961, 8.303739, 8.298015, 8.36177, 8.325923, 
    8.379751, 8.376764, 8.352378, 8.377101, 8.138278, 8.131471, 8.107876, 
    8.126336, 8.092727, 8.111527, 8.122355, 8.164235, 8.173457, 8.18202, 
    8.19895, 8.22072, 8.259025, 8.292467, 8.323089, 8.320842, 8.321633, 
    8.328486, 8.311521, 8.331274, 8.334595, 8.325917, 8.376365, 8.361928, 
    8.376701, 8.367298, 8.133683, 8.145142, 8.138948, 8.150599, 8.14239, 
    8.178944, 8.189929, 8.241487, 8.220292, 8.254041, 8.223714, 8.229082, 
    8.255149, 8.225349, 8.290623, 8.246329, 8.328753, 8.284363, 8.331541, 
    8.322956, 8.337173, 8.349923, 8.365983, 8.395685, 8.388799, 8.413684, 
    8.162248, 8.177156, 8.175841, 8.191463, 8.203032, 8.228151, 8.268572, 
    8.253352, 8.281307, 8.286929, 8.244465, 8.270519, 8.187145, 8.200572, 
    8.192574, 8.163424, 8.256861, 8.208803, 8.29772, 8.271553, 8.348104, 
    8.309966, 8.385011, 8.417263, 8.447694, 8.48338, 8.185301, 8.175159, 
    8.193322, 8.218509, 8.241927, 8.273148, 8.276346, 8.282207, 8.297404, 
    8.3102, 8.284064, 8.31341, 8.203693, 8.261042, 8.17133, 8.198265, 
    8.217021, 8.208786, 8.251614, 8.261735, 8.302967, 8.281631, 8.409296, 
    8.352622, 8.510624, 8.466235, 8.171619, 8.185265, 8.2329, 8.210207, 
    8.275234, 8.291305, 8.304385, 8.321135, 8.322943, 8.332881, 8.316601, 
    8.332236, 8.273214, 8.299548, 8.227441, 8.244946, 8.236888, 8.228059, 
    8.255334, 8.284476, 8.285095, 8.294459, 8.320896, 8.275498, 8.41664, 
    8.329257, 8.200164, 8.226542, 8.23031, 8.220081, 8.289693, 8.264416, 
    8.332638, 8.314155, 8.344455, 8.329388, 8.327172, 8.307856, 8.295849, 
    8.265574, 8.241006, 8.221564, 8.226081, 8.247449, 8.286261, 8.323108, 
    8.315026, 8.342149, 8.270505, 8.300488, 8.288891, 8.319158, 8.25295, 
    8.309315, 8.238593, 8.244773, 8.263915, 8.302528, 8.311085, 8.320235, 
    8.314587, 8.287247, 8.282773, 8.263448, 8.258121, 8.243427, 8.231279, 
    8.242378, 8.254048, 8.287256, 8.317277, 8.350105, 8.358153, 8.39668, 
    8.365313, 8.41713, 8.373068, 8.449453, 8.312585, 8.371766, 8.264785, 
    8.276257, 8.297042, 8.344864, 8.319016, 8.34925, 8.282598, 8.248189, 
    8.239301, 8.222746, 8.239679, 8.238301, 8.254529, 8.249311, 8.288361, 
    8.267366, 8.327118, 8.34901, 8.411075, 8.449306, 8.488356, 8.505643, 
    8.51091, 8.513112,
  12.66457, 12.72003, 12.70923, 12.7541, 12.72919, 12.7586, 12.6758, 
    12.72224, 12.69257, 12.66955, 12.8416, 12.75611, 12.93095, 12.87601, 
    13.01443, 12.92239, 13.03306, 13.01176, 13.07595, 13.05753, 13.13997, 
    13.08446, 13.18288, 13.12669, 13.13547, 13.08263, 12.77326, 12.83093, 
    12.76985, 12.77806, 12.77438, 12.72971, 12.70726, 12.66034, 12.66884, 
    12.70331, 12.78175, 12.75507, 12.82241, 12.82088, 12.89623, 12.86221, 
    12.98947, 12.95318, 13.0583, 13.03179, 13.05705, 13.04939, 13.05715, 
    13.01829, 13.03493, 13.00078, 12.86858, 12.9073, 12.79212, 12.72334, 
    12.67783, 12.64563, 12.65018, 12.65885, 12.70351, 12.74562, 12.77781, 
    12.79938, 12.82066, 12.88531, 12.91964, 12.99682, 12.98286, 13.00652, 
    13.02915, 13.06725, 13.06097, 13.07778, 13.00589, 13.05363, 12.97491, 
    12.9964, 12.82648, 12.76226, 12.73508, 12.71131, 12.65368, 12.69345, 
    12.67776, 12.71512, 12.73891, 12.72714, 12.79997, 12.77161, 12.92168, 
    12.85684, 13.02651, 12.98572, 13.03631, 13.01047, 13.05477, 13.01489, 
    13.08404, 13.09914, 13.08882, 13.12851, 13.01269, 13.05706, 12.72681, 
    12.72873, 12.73768, 12.6984, 12.696, 12.66011, 12.69204, 12.70566, 
    12.74029, 12.76083, 12.78037, 12.82344, 12.87171, 12.93947, 12.98836, 
    13.02123, 13.00107, 13.01887, 12.99897, 12.98965, 13.09348, 13.03509, 
    13.12279, 13.11792, 13.07818, 13.11847, 12.73008, 12.71903, 12.68077, 
    12.7107, 12.6562, 12.68669, 12.70425, 12.7722, 12.78718, 12.80108, 
    12.82858, 12.86395, 12.92622, 12.98062, 13.03047, 13.02681, 13.0281, 
    13.03926, 13.01164, 13.0438, 13.04921, 13.03508, 13.11727, 13.09374, 
    13.11782, 13.10249, 12.72262, 12.74122, 12.73117, 12.75007, 12.73675, 
    12.79608, 12.81392, 12.8977, 12.86325, 12.91811, 12.86881, 12.87754, 
    12.91992, 12.87147, 12.97762, 12.90557, 13.0397, 12.96744, 13.04424, 
    13.03026, 13.05341, 13.07418, 13.10035, 13.14877, 13.13754, 13.17813, 
    12.76898, 12.79318, 12.79105, 12.81642, 12.83521, 12.87603, 12.94175, 
    12.917, 12.96247, 12.97161, 12.90254, 12.94491, 12.8094, 12.83121, 
    12.81822, 12.77089, 12.9227, 12.84458, 12.98917, 12.9466, 13.07122, 
    13.00911, 13.13137, 13.18397, 13.23363, 13.29191, 12.80641, 12.78994, 
    12.81944, 12.86035, 12.89842, 12.94919, 12.95439, 12.96393, 12.98866, 
    13.00949, 12.96695, 13.01471, 12.83628, 12.9295, 12.78372, 12.82746, 
    12.85794, 12.84456, 12.91417, 12.93063, 12.99771, 12.96299, 13.17097, 
    13.07858, 13.33643, 13.2639, 12.78419, 12.80635, 12.88374, 12.84686, 
    12.95258, 12.97873, 13.00002, 13.02729, 13.03023, 13.04642, 13.01991, 
    13.04537, 12.9493, 12.99215, 12.87487, 12.90333, 12.89023, 12.87587, 
    12.92022, 12.96762, 12.96863, 12.98387, 13.0269, 12.95301, 13.18295, 
    13.04052, 12.83055, 12.87341, 12.87953, 12.86291, 12.97611, 12.93499, 
    13.04602, 13.01593, 13.06527, 13.04073, 13.03712, 13.00567, 12.98613, 
    12.93687, 12.89692, 12.86532, 12.87266, 12.9074, 12.97052, 13.0305, 
    13.01734, 13.06151, 12.94489, 12.99368, 12.9748, 13.02407, 12.91634, 
    13.00805, 12.893, 12.90304, 12.93417, 12.997, 13.01093, 13.02583, 
    13.01663, 12.97213, 12.96485, 12.93341, 12.92475, 12.90086, 12.88111, 
    12.89915, 12.91813, 12.97215, 13.02101, 13.07448, 13.08759, 13.15039, 
    13.09926, 13.18375, 13.1119, 13.2365, 13.01337, 13.10977, 12.93559, 
    12.95425, 12.98807, 13.06594, 13.02384, 13.07308, 12.96456, 12.9086, 
    12.89415, 12.86724, 12.89476, 12.89252, 12.91891, 12.91042, 12.97394, 
    12.93979, 13.03703, 13.07269, 13.17387, 13.23626, 13.30004, 13.32829, 
    13.33689, 13.34049,
  20.59555, 20.6916, 20.67289, 20.75065, 20.70747, 20.75845, 20.61498, 
    20.69543, 20.64403, 20.60417, 20.90253, 20.75413, 21.05791, 20.96234, 
    21.20336, 21.04301, 21.23585, 21.1987, 21.31072, 21.27856, 21.4226, 
    21.32558, 21.49769, 21.39938, 21.41473, 21.32239, 20.78389, 20.88399, 
    20.77798, 20.79221, 20.78582, 20.70836, 20.66946, 20.58822, 20.60294, 
    20.66262, 20.79862, 20.75233, 20.86918, 20.86654, 20.9975, 20.93834, 
    21.15984, 21.09661, 21.2799, 21.23364, 21.27773, 21.26435, 21.2779, 
    21.2101, 21.23912, 21.17956, 20.9494, 21.01675, 20.81661, 20.69733, 
    20.6185, 20.56278, 20.57064, 20.58566, 20.66297, 20.73595, 20.79177, 
    20.8292, 20.86616, 20.9785, 21.03822, 21.17266, 21.14831, 21.18956, 
    21.22904, 21.29552, 21.28456, 21.31391, 21.18847, 21.27175, 21.13446, 
    21.17191, 20.87625, 20.7648, 20.71767, 20.67648, 20.5767, 20.64555, 
    20.61838, 20.68308, 20.72432, 20.70391, 20.83022, 20.78102, 21.04177, 
    20.929, 21.22443, 21.15331, 21.24152, 21.19645, 21.27374, 21.20417, 
    21.32484, 21.35123, 21.3332, 21.40255, 21.20032, 21.27773, 20.70334, 
    20.70667, 20.72218, 20.65412, 20.64996, 20.58782, 20.6431, 20.66669, 
    20.72671, 20.76231, 20.79622, 20.87098, 20.95484, 21.07274, 21.15791, 
    21.21522, 21.18005, 21.21109, 21.1764, 21.16016, 21.34134, 21.23939, 
    21.39256, 21.38405, 21.31461, 21.38501, 20.70901, 20.68987, 20.62358, 
    20.67544, 20.58107, 20.63383, 20.66425, 20.78205, 20.80803, 20.83216, 
    20.8799, 20.94136, 21.04967, 21.14442, 21.23134, 21.22495, 21.2272, 
    21.24667, 21.19848, 21.2546, 21.26403, 21.23937, 21.38291, 21.34179, 
    21.38387, 21.35708, 20.69608, 20.72831, 20.71089, 20.74366, 20.72057, 
    20.82349, 20.85446, 21.00005, 20.94015, 21.03556, 20.94982, 20.96498, 
    21.0387, 20.95444, 21.13919, 21.01375, 21.24743, 21.12144, 21.25536, 
    21.23096, 21.27136, 21.30763, 21.35334, 21.43799, 21.41836, 21.48936, 
    20.77645, 20.81845, 20.81474, 20.85878, 20.89142, 20.96235, 21.0767, 
    21.03362, 21.11278, 21.12872, 21.00847, 21.08222, 20.84661, 20.88448, 
    20.86192, 20.77977, 21.04355, 20.90771, 21.15932, 21.08515, 21.30245, 
    21.19407, 21.40755, 21.49958, 21.58658, 21.68879, 20.84141, 20.81282, 
    20.86403, 20.93511, 21.0013, 21.08966, 21.09872, 21.11534, 21.15843, 
    21.19474, 21.1206, 21.20385, 20.89328, 21.05538, 20.80204, 20.87797, 
    20.93091, 20.90766, 21.0287, 21.05734, 21.17421, 21.1137, 21.47684, 
    21.3153, 21.76696, 21.63965, 20.80285, 20.8413, 20.97577, 20.91167, 
    21.09557, 21.14113, 21.17823, 21.22579, 21.23092, 21.25916, 21.21291, 
    21.25733, 21.08985, 21.16451, 20.96035, 21.00983, 20.98705, 20.96209, 
    21.03922, 21.12177, 21.12352, 21.15007, 21.22511, 21.09632, 21.4978, 
    21.24886, 20.88333, 20.95781, 20.96846, 20.93955, 21.13655, 21.06493, 
    21.25847, 21.20596, 21.29207, 21.24924, 21.24294, 21.18808, 21.15401, 
    21.06821, 20.99869, 20.94374, 20.9565, 21.01691, 21.12682, 21.23139, 
    21.20844, 21.28551, 21.08218, 21.16718, 21.13428, 21.22017, 21.03248, 
    21.19222, 20.99187, 21.00935, 21.06351, 21.17296, 21.19725, 21.22323, 
    21.20719, 21.12962, 21.11694, 21.06219, 21.04711, 21.00554, 20.97119, 
    21.00257, 21.03559, 21.12965, 21.21483, 21.30814, 21.33105, 21.44083, 
    21.35143, 21.4992, 21.37352, 21.59161, 21.20151, 21.36981, 21.06598, 
    21.09847, 21.1574, 21.29324, 21.21977, 21.30571, 21.11644, 21.01901, 
    20.99387, 20.94708, 20.99494, 20.99104, 21.03695, 21.02218, 21.13278, 
    21.07329, 21.24279, 21.30503, 21.48191, 21.59119, 21.70305, 21.75266, 
    21.76778, 21.77411,
  34.63898, 34.81974, 34.78448, 34.93107, 34.84964, 34.94579, 34.67551, 
    34.82695, 34.73016, 34.65519, 35.21814, 34.93763, 35.51294, 35.33147, 
    35.78992, 35.48462, 35.85194, 35.78104, 35.99503, 35.93353, 36.20937, 
    36.02347, 36.35357, 36.16483, 36.19426, 36.01736, 34.9938, 35.18304, 
    34.98264, 35.00952, 34.99745, 34.85132, 34.77803, 34.62521, 34.65288, 
    34.76515, 35.02161, 34.93423, 35.15502, 35.15001, 35.39818, 35.28597, 
    35.70694, 35.58654, 35.93609, 35.84771, 35.93194, 35.90636, 35.93227, 
    35.80278, 35.85817, 35.74453, 35.30695, 35.43474, 35.05562, 34.83053, 
    34.68213, 34.5774, 34.59218, 34.62038, 34.76581, 34.90334, 35.00868, 
    35.07941, 35.1493, 35.36214, 35.47552, 35.73137, 35.68498, 35.7636, 
    35.83894, 35.96596, 35.945, 36.00114, 35.76151, 35.92051, 35.6586, 
    35.72995, 35.1684, 34.95778, 34.86886, 34.79126, 34.60355, 34.73302, 
    34.6819, 34.80369, 34.88141, 34.84294, 35.08134, 34.98838, 35.48226, 
    35.26828, 35.83014, 35.69449, 35.86276, 35.77674, 35.92432, 35.79146, 
    36.02205, 36.07257, 36.03804, 36.17092, 35.78412, 35.93194, 34.84186, 
    34.84813, 34.87736, 34.74915, 34.74133, 34.62445, 34.72841, 34.77283, 
    34.88592, 34.95307, 35.01708, 35.15842, 35.31726, 35.54114, 35.70326, 
    35.81255, 35.74547, 35.80468, 35.7385, 35.70755, 36.05363, 35.8587, 
    36.15176, 36.13545, 36.00248, 36.13729, 34.85254, 34.81647, 34.69169, 
    34.78928, 34.61176, 34.71098, 34.76822, 34.99033, 35.03939, 35.085, 
    35.1753, 35.2917, 35.49728, 35.67757, 35.84332, 35.83113, 35.83543, 
    35.8726, 35.78062, 35.88774, 35.90577, 35.85867, 36.13327, 36.05449, 
    36.1351, 36.08378, 34.82819, 34.88893, 34.85609, 34.91788, 34.87434, 
    35.0686, 35.12716, 35.40303, 35.28941, 35.47047, 35.30774, 35.33649, 
    35.47643, 35.3165, 35.6676, 35.42903, 35.87405, 35.6338, 35.88919, 
    35.8426, 35.91978, 35.98911, 36.07661, 36.23891, 36.20123, 36.33757, 
    34.97977, 35.05909, 35.05208, 35.13534, 35.19711, 35.33151, 35.54867, 
    35.46677, 35.61732, 35.64766, 35.41902, 35.55915, 35.11231, 35.18396, 
    35.14127, 34.98602, 35.48564, 35.22794, 35.70595, 35.56473, 35.97921, 
    35.77221, 36.18051, 36.35721, 36.52464, 36.72184, 35.10248, 35.04845, 
    35.14526, 35.27986, 35.4054, 35.57332, 35.59056, 35.62218, 35.70425, 
    35.77348, 35.63219, 35.79086, 35.20063, 35.50813, 35.02807, 35.17164, 
    35.2719, 35.22786, 35.45743, 35.51186, 35.73433, 35.61906, 36.31349, 
    36.0038, 36.87302, 36.62698, 35.02961, 35.10229, 35.35696, 35.23545, 
    35.58456, 35.67129, 35.742, 35.83272, 35.84253, 35.89646, 35.80815, 
    35.89296, 35.57368, 35.71584, 35.3277, 35.4216, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63776, 35.68833, 35.83143, 35.58599, 36.35379, 
    35.87679, 35.18179, 35.32288, 35.34308, 35.28828, 35.66258, 35.52629, 
    35.89514, 35.79489, 35.95936, 35.87749, 35.86547, 35.76078, 35.69584, 
    35.53252, 35.40045, 35.29622, 35.32042, 35.43505, 35.64405, 35.84343, 
    35.79961, 35.94682, 35.55908, 35.72092, 35.65825, 35.82201, 35.4646, 
    35.76868, 35.3875, 35.42068, 35.52359, 35.73195, 35.77826, 35.82785, 
    35.79724, 35.64937, 35.62523, 35.52108, 35.49241, 35.41345, 35.34827, 
    35.40782, 35.47051, 35.64943, 35.81181, 35.9901, 36.03392, 36.24435, 
    36.07294, 36.35648, 36.11526, 36.53433, 35.78639, 36.10815, 35.52828, 
    35.59008, 35.70229, 35.96159, 35.82123, 35.98545, 35.62428, 35.43902, 
    35.3913, 35.30255, 35.39333, 35.38593, 35.4731, 35.44505, 35.65539, 
    35.54218, 35.86518, 35.98414, 36.32325, 36.53352, 36.7494, 36.84534, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34589, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59598, 62.19373, 
    63.21417, 62.53307, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73952, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13967, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47564, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13955, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25315, 61.48349, 
    61.63854, 61.79207, 62.26156, 62.51286, 63.08306, 62.97935, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.6428, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73633, 63.85044, 63.77242, 64.07315, 63.20119, 63.5332, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36182, 61.5019, 61.81213, 62.16233, 62.65869, 63.02021, 
    63.26492, 63.11462, 63.24727, 63.09903, 63.02979, 63.80764, 63.36849, 
    64.02972, 63.99276, 63.69214, 63.99692, 61.14231, 61.06372, 60.79243, 
    61.00454, 60.61915, 60.8343, 60.95869, 61.44333, 61.55079, 61.65081, 
    61.84928, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31625, 
    63.39974, 63.19335, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18986, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40972, 63.40299, 62.86511, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59398, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49344, 62.82833, 62.89602, 62.38752, 62.69877, 61.71079, 61.86834, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.09491, 64.49689, 64.87986, 65.33361, 61.68919, 61.57066, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86152, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75535, 62.94876, 63.10686, 63.31018, 63.33219, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29745, 62.19272, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86355, 62.17475, 62.2194, 62.09832, 62.92932, 62.62566, 
    63.4504, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00362, 
    62.63952, 62.34638, 62.11584, 62.16929, 62.42306, 62.88795, 63.3342, 
    63.23591, 63.5667, 62.69861, 63.0597, 62.91965, 63.28613, 62.48863, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26327, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65374, 62.84386, 62.43187, 
    62.3261, 62.12982, 62.33061, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38306, 63.65079, 64.41946, 64.90024, 65.39728, 65.61928, 
    65.68716, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7406, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02024528, -0.01991452, -0.01997837, -0.0197149, -0.0198606, -0.01968874, 
    -0.02017776, -0.01990149, -0.02007739, -0.02021528, -0.01921416, 
    -0.01970324, -0.01872008, -0.01902185, -0.0182736, -0.01876668, 
    -0.01817589, -0.01828766, -0.01795356, -0.0180486, -0.01762841, 
    -0.01790988, -0.01741482, -0.01769521, -0.01765101, -0.01791925, 
    -0.01960378, -0.01927432, -0.01962348, -0.01957608, -0.01959734, 
    -0.01985757, -0.01999009, -0.02027082, -0.02021955, -0.02001352, 
    -0.01955481, -0.01970926, -0.01932255, -0.0193312, -0.01891004, 
    -0.01909869, -0.01840561, -0.0185998, -0.01804462, -0.01818253, 
    -0.01805107, -0.01809083, -0.01805055, -0.01825327, -0.01816612, 
    -0.01834561, -0.0190632, -0.01884921, -0.01949521, -0.01989503, 
    -0.02016555, -0.02035988, -0.02033229, -0.02027979, -0.02001232, 
    -0.01976433, -0.01957756, -0.01945367, -0.01933244, -0.01897032, 
    -0.01878169, -0.01836659, -0.01844079, -0.0183153, -0.01819631, 
    -0.01799838, -0.01803081, -0.01794417, -0.01831862, -0.01806882, 
    -0.0184832, -0.01836884, -0.01929951, -0.01966747, -0.01982605, 
    -0.01996607, -0.0203111, -0.02007215, -0.02016598, -0.01994354, 
    -0.01980356, -0.01987266, -0.0194503, -0.01961334, -0.01877058, 
    -0.0191287, -0.01821015, -0.01842554, -0.01815893, -0.01829445, 
    -0.0180629, -0.01827115, -0.01791205, -0.01783486, -0.01788757, 
    -0.01768605, -0.01828277, -0.01805106, -0.0198746, -0.01986331, 
    -0.01981081, -0.02004269, -0.02005697, -0.02027223, -0.02008058, 
    -0.01999956, -0.01979548, -0.01967581, -0.01956278, -0.0193167, 
    -0.01904579, -0.01867385, -0.01841149, -0.01823785, -0.01834412, 
    -0.01825027, -0.01835521, -0.01840463, -0.01786373, -0.0181653, 
    -0.01771488, -0.01773949, -0.01794211, -0.01773672, -0.01985539, 
    -0.01992042, -0.02014796, -0.01996966, -0.02029582, -0.02011253, 
    -0.02000794, -0.01960989, -0.01952361, -0.01944393, -0.01928763, 
    -0.01908899, -0.01874583, -0.01845269, -0.01818942, -0.01820857, 
    -0.01820183, -0.01814352, -0.01828831, -0.01811987, -0.01809175, 
    -0.01816535, -0.01774279, -0.01786241, -0.01774001, -0.0178178, 
    -0.01989926, -0.01979009, -0.019849, -0.01973837, -0.01981623, 
    -0.01947251, -0.01937071, -0.01890196, -0.01909287, -0.01879003, 
    -0.01906188, -0.0190134, -0.0187802, -0.01904709, -0.0184687, 
    -0.01885868, -0.01814125, -0.01852318, -0.0181176, -0.01819055, 
    -0.01806996, -0.01796268, -0.01782871, -0.01758431, -0.01764059, 
    -0.01743831, -0.01962855, -0.01948913, -0.01950139, -0.01935655, 
    -0.01925017, -0.01902179, -0.01866154, -0.01879614, -0.01854985, 
    -0.01850082, -0.01887533, -0.01864441, -0.01939644, -0.01927274, 
    -0.0193463, -0.0196175, -0.018765, -0.0191974, -0.01840718, -0.01863532, 
    -0.01797793, -0.01830165, -0.01767164, -0.01740947, -0.01716666, 
    -0.01688746, -0.01941352, -0.01950774, -0.01933941, -0.01910905, 
    -0.01889802, -0.01862131, -0.01859326, -0.01854199, -0.01840991, 
    -0.01829964, -0.01852579, -0.01827211, -0.01924413, -0.01872798, 
    -0.01954346, -0.01929392, -0.01912256, -0.01919755, -0.0188116, 
    -0.01872185, -0.01836187, -0.01854703, -0.01747376, -0.01794007, 
    -0.01667824, -0.01702086, -0.01954076, -0.01941385, -0.01897901, 
    -0.01918459, -0.01860301, -0.01846278, -0.01834964, -0.01820608, 
    -0.01819067, -0.01810626, -0.0182448, -0.01811172, -0.01862073, 
    -0.01839138, -0.0190282, -0.01887103, -0.01894317, -0.01902262, 
    -0.01877855, -0.0185222, -0.0185168, -0.01843542, -0.01820811, 
    -0.01860069, -0.01741448, -0.01813698, -0.01927648, -0.01903632, 
    -0.01900232, -0.01909478, -0.01847679, -0.01869817, -0.01810832, 
    -0.01826573, -0.01800859, -0.01813587, -0.01815468, -0.01831978, 
    -0.01842338, -0.01868795, -0.01890626, -0.01908134, -0.01904048, 
    -0.01884869, -0.01850665, -0.01818926, -0.01825827, -0.01802799, 
    -0.01864453, -0.01838325, -0.01848375, -0.01822295, -0.01879973, 
    -0.01830724, -0.01892788, -0.01887257, -0.0187026, -0.01836565, 
    -0.01829205, -0.01821375, -0.01826203, -0.01849806, -0.01853706, 
    -0.01870672, -0.01875384, -0.0188846, -0.01899359, -0.01889398, 
    -0.01878996, -0.01849797, -0.01823901, -0.01796115, -0.01789386, 
    -0.01757621, -0.01783428, -0.01741054, -0.01777002, -0.01715276, 
    -0.01827918, -0.01778078, -0.01869491, -0.01859404, -0.01841304, 
    -0.01800514, -0.01822416, -0.01796832, -0.01853859, -0.01884209, 
    -0.01892153, -0.01907064, -0.01891814, -0.0189305, -0.01878569, 
    -0.0188321, -0.01848836, -0.01867215, -0.01815514, -0.01797033, 
    -0.01745938, -0.01715393, -0.016849, -0.01671624, -0.01667606, -0.01665929,
  -0.05398342, -0.05294037, -0.05314149, -0.05231233, -0.05277063, 
    -0.05223012, -0.05377026, -0.05289936, -0.05345362, -0.0538887, 
    -0.0507418, -0.05227568, -0.04919917, -0.05014054, -0.04781123, 
    -0.04934436, -0.04750828, -0.04785486, -0.04682, -0.04711403, 
    -0.04581604, -0.04668495, -0.04515833, -0.04602204, -0.04588573, 
    -0.0467139, -0.05196321, -0.05093011, -0.05202508, -0.05187624, 
    -0.051943, -0.05276108, -0.05317841, -0.0540641, -0.05390218, 
    -0.05325226, -0.05180946, -0.05229462, -0.0510812, -0.05110827, 
    -0.04979146, -0.05038068, -0.04822098, -0.04882469, -0.04710172, 
    -0.04752886, -0.04712167, -0.04724476, -0.04712007, -0.04774819, 
    -0.04747799, -0.04803471, -0.05026975, -0.04960166, -0.05162242, 
    -0.05287901, -0.05373173, -0.05434553, -0.05425831, -0.05409242, 
    -0.05324848, -0.05246776, -0.05188088, -0.05149215, -0.05111216, 
    -0.0499796, -0.04939116, -0.04809982, -0.04833029, -0.04794062, 
    -0.04757158, -0.04695864, -0.04705896, -0.04679095, -0.04795092, 
    -0.04717662, -0.04846207, -0.04810683, -0.05100899, -0.05216328, 
    -0.0526619, -0.05310276, -0.05419134, -0.05343708, -0.05373307, 
    -0.05303178, -0.05259114, -0.05280861, -0.05148157, -0.05199324, 
    -0.04935652, -0.0504745, -0.04761447, -0.0482829, -0.04745573, 
    -0.04787594, -0.04715829, -0.04780365, -0.04669164, -0.04645312, 
    -0.04661597, -0.0459938, -0.04783969, -0.04712164, -0.05281469, 
    -0.05277916, -0.05261396, -0.05334419, -0.05338923, -0.05406853, 
    -0.05346368, -0.05320825, -0.05256574, -0.05218949, -0.05183448, 
    -0.05106285, -0.05021534, -0.04905518, -0.04823926, -0.04770038, 
    -0.04803008, -0.04773887, -0.04806451, -0.04821797, -0.04654232, 
    -0.04747546, -0.04608274, -0.04615868, -0.04678458, -0.04615011, 
    -0.05275422, -0.05295897, -0.05367622, -0.05311404, -0.05414306, 
    -0.05356445, -0.05323468, -0.05198241, -0.05171155, -0.05146161, 
    -0.05097179, -0.05035034, -0.04927941, -0.04836726, -0.04755022, 
    -0.04760959, -0.04758868, -0.04740797, -0.04785688, -0.0473347, 
    -0.04724763, -0.04747561, -0.04616885, -0.04653825, -0.04616029, 
    -0.04640042, -0.05289233, -0.05254878, -0.05273412, -0.05238614, 
    -0.05263101, -0.05155123, -0.05123207, -0.04976623, -0.05036248, 
    -0.04941716, -0.05026562, -0.05011414, -0.04938649, -0.0502194, 
    -0.04841701, -0.04963122, -0.04740096, -0.04858637, -0.0473277, 
    -0.04755372, -0.04718015, -0.04684818, -0.04643412, -0.04568016, 
    -0.0458536, -0.04523061, -0.05204101, -0.05160338, -0.05164182, 
    -0.05118769, -0.05085453, -0.05014035, -0.04901686, -0.04943621, 
    -0.04866932, -0.04851686, -0.04968315, -0.04896353, -0.05131272, 
    -0.05092518, -0.0511556, -0.0520063, -0.04933915, -0.05068937, 
    -0.04822589, -0.04893523, -0.04689535, -0.04789826, -0.04594936, 
    -0.04514188, -0.04439595, -0.04354046, -0.05136625, -0.05166174, 
    -0.05113399, -0.05041305, -0.04975394, -0.04889164, -0.04880435, 
    -0.04864485, -0.04823436, -0.04789202, -0.04859447, -0.04780662, 
    -0.0508356, -0.04922378, -0.05177386, -0.05099151, -0.05045528, 
    -0.05068984, -0.0494844, -0.0492047, -0.04808518, -0.04866054, 
    -0.0453397, -0.04677828, -0.04290105, -0.04394891, -0.05176539, 
    -0.0513673, -0.05000674, -0.0506493, -0.04883468, -0.04839861, 
    -0.04804722, -0.04760185, -0.04755408, -0.04729256, -0.04772191, 
    -0.04730946, -0.04888982, -0.0481768, -0.0501604, -0.04966974, 
    -0.04989485, -0.05014296, -0.04938137, -0.04858331, -0.04856652, 
    -0.04831359, -0.04760814, -0.04882747, -0.04515729, -0.0473877, 
    -0.05093689, -0.05018574, -0.05007954, -0.05036845, -0.04844214, 
    -0.04913094, -0.04729893, -0.04778683, -0.0469902, -0.04738428, 
    -0.04744254, -0.04795452, -0.04827619, -0.04909911, -0.04977965, 
    -0.05032645, -0.05019875, -0.04960006, -0.04853496, -0.04754971, 
    -0.04776369, -0.04705025, -0.04896391, -0.04815157, -0.0484638, 
    -0.04765415, -0.04944738, -0.0479156, -0.04984713, -0.04967456, 
    -0.04914472, -0.04809691, -0.04786848, -0.04762563, -0.04777535, 
    -0.04850826, -0.04862952, -0.04915755, -0.04930435, -0.04971208, 
    -0.05005229, -0.04974133, -0.04941694, -0.048508, -0.04770397, 
    -0.04684346, -0.04663543, -0.04565518, -0.04645132, -0.04514516, 
    -0.0462529, -0.04435328, -0.04782855, -0.04628612, -0.04912079, 
    -0.04880678, -0.04824409, -0.04697954, -0.04765792, -0.04686563, 
    -0.04863428, -0.04957948, -0.04982732, -0.05029301, -0.04981673, 
    -0.04985529, -0.04940363, -0.04954831, -0.04847813, -0.04904991, 
    -0.04744398, -0.04687186, -0.04529544, -0.04435688, -0.04342283, 
    -0.04301708, -0.0428944, -0.04284322,
  -0.07871159, -0.0770606, -0.07737876, -0.07606762, -0.07679213, 
    -0.07593769, -0.07837401, -0.07699572, -0.07787271, -0.07856157, 
    -0.07358827, -0.07600968, -0.07115836, -0.07264054, -0.06897684, 
    -0.07138684, -0.06850127, -0.06904534, -0.06742165, -0.06788272, 
    -0.06584895, -0.06720995, -0.06482, -0.06617143, -0.06595804, 
    -0.06725533, -0.07551599, -0.07388527, -0.07561374, -0.07537863, 
    -0.07548407, -0.07677703, -0.07743717, -0.07883939, -0.07858291, 
    -0.07755403, -0.07527316, -0.07603963, -0.07412359, -0.07416631, 
    -0.07209067, -0.07301896, -0.0696204, -0.07056932, -0.06786341, 
    -0.06853357, -0.06789471, -0.06808779, -0.06789219, -0.06887786, 
    -0.06845374, -0.06932779, -0.07284413, -0.07179184, -0.07497781, 
    -0.07696354, -0.07831299, -0.0792853, -0.07914709, -0.07888426, 
    -0.07754805, -0.07631329, -0.07538595, -0.07477215, -0.07417245, 
    -0.07238701, -0.07146049, -0.06943006, -0.06979214, -0.06918001, 
    -0.06860062, -0.06763902, -0.06779635, -0.06737611, -0.06919619, 
    -0.06798089, -0.06999924, -0.06944107, -0.07400969, -0.07583208, 
    -0.0766202, -0.07731747, -0.07904097, -0.07784652, -0.07831512, 
    -0.07720519, -0.07650832, -0.07685219, -0.07475544, -0.07556343, 
    -0.07140596, -0.07316684, -0.06866794, -0.06971768, -0.0684188, 
    -0.06907845, -0.06795215, -0.06896494, -0.06722044, -0.06684665, 
    -0.06710184, -0.06612722, -0.06902152, -0.06789466, -0.07686181, 
    -0.07680561, -0.0765444, -0.0776995, -0.07777078, -0.07884641, 
    -0.07788863, -0.07748438, -0.07646817, -0.07587349, -0.07531266, 
    -0.07409465, -0.0727584, -0.07093184, -0.06964912, -0.0688028, 
    -0.06932051, -0.06886323, -0.06937461, -0.06961567, -0.06698641, 
    -0.06844977, -0.06626649, -0.0663854, -0.06736613, -0.06637199, 
    -0.07676619, -0.07709, -0.0782251, -0.07733532, -0.07896448, -0.07804814, 
    -0.07752621, -0.07554632, -0.07511854, -0.07472393, -0.07395101, 
    -0.07297114, -0.07128462, -0.06985024, -0.0685671, -0.06866028, 
    -0.06862746, -0.06834386, -0.06904851, -0.0682289, -0.06809229, -0.06845, 
    -0.06640134, -0.06698004, -0.06638793, -0.06676406, -0.0769846, 
    -0.07644135, -0.07673439, -0.07618427, -0.07657136, -0.07486542, 
    -0.07436167, -0.07205095, -0.07299027, -0.07150141, -0.07283762, 
    -0.07259894, -0.07145315, -0.07276479, -0.06992844, -0.07183836, 
    -0.06833287, -0.07019462, -0.0682179, -0.0685726, -0.06798644, 
    -0.06746583, -0.06681687, -0.06563628, -0.06590774, -0.06493301, 
    -0.0756389, -0.07494774, -0.07500844, -0.07429162, -0.07376605, 
    -0.07264024, -0.07087156, -0.07153139, -0.07032502, -0.07008536, 
    -0.07192013, -0.07078768, -0.07448892, -0.07387748, -0.07424098, 
    -0.07558407, -0.07137863, -0.07350559, -0.06962811, -0.07074317, 
    -0.0675398, -0.06911349, -0.06605764, -0.06479426, -0.06362867, 
    -0.06229363, -0.07457342, -0.07503989, -0.07420689, -0.07306998, 
    -0.07203159, -0.07067461, -0.07053733, -0.07028656, -0.06964142, 
    -0.0691037, -0.07020736, -0.06896959, -0.0737362, -0.07119709, 
    -0.07521693, -0.07398211, -0.07313655, -0.07350634, -0.07160723, 
    -0.07116706, -0.06940706, -0.07031122, -0.06510364, -0.06735626, 
    -0.06129704, -0.06293081, -0.07520355, -0.07457507, -0.07242975, 
    -0.07344241, -0.07058503, -0.06989951, -0.06934743, -0.06864814, 
    -0.06857315, -0.06816277, -0.06883659, -0.06818929, -0.07067174, 
    -0.06955099, -0.07267182, -0.07189901, -0.0722535, -0.07264435, 
    -0.07144507, -0.07018981, -0.07016341, -0.06976591, -0.06865802, 
    -0.0705737, -0.06481837, -0.06831207, -0.07389595, -0.07271175, 
    -0.07254443, -0.07299968, -0.06996793, -0.07105102, -0.06817277, 
    -0.06893852, -0.06768852, -0.06830668, -0.06839811, -0.06920184, 
    -0.06970714, -0.07100094, -0.07207208, -0.07293349, -0.07273225, 
    -0.07178931, -0.07011382, -0.06856629, -0.06890219, -0.06778269, 
    -0.07078827, -0.06951135, -0.07000197, -0.06873023, -0.07154897, 
    -0.06914073, -0.07217835, -0.0719066, -0.07107269, -0.0694255, 
    -0.06906672, -0.06868546, -0.06892049, -0.07007185, -0.07026245, 
    -0.07109288, -0.07132387, -0.07196568, -0.0725015, -0.07201174, 
    -0.07150106, -0.07007143, -0.06880843, -0.06745843, -0.06713233, 
    -0.06559718, -0.06684383, -0.06479941, -0.06653298, -0.06356204, 
    -0.06900404, -0.06658502, -0.07103504, -0.07054116, -0.06965671, 
    -0.06767181, -0.06873615, -0.06749319, -0.07026994, -0.07175691, 
    -0.07214715, -0.07288078, -0.07213047, -0.0721912, -0.07148012, 
    -0.07170784, -0.07002448, -0.07092354, -0.06840037, -0.06750296, 
    -0.0650344, -0.06356765, -0.0621102, -0.06147781, -0.06128668, -0.06120696,
  -0.08618353, -0.0842735, -0.08464148, -0.08312541, -0.08396304, 
    -0.08297522, -0.08579287, -0.08419849, -0.08521286, -0.08600992, 
    -0.08026101, -0.08305844, -0.07745697, -0.07916696, -0.07494242, 
    -0.07772048, -0.07439461, -0.07502132, -0.07315152, -0.07368232, 
    -0.07134197, -0.07290785, -0.07015889, -0.0717129, -0.07146744, 
    -0.07296007, -0.08248783, -0.08060396, -0.08260079, -0.08232908, 
    -0.08245093, -0.08394559, -0.08470905, -0.08633144, -0.08603462, 
    -0.08484421, -0.0822072, -0.08309304, -0.08087918, -0.08092851, 
    -0.07853243, -0.07960374, -0.07568394, -0.07677773, -0.07366008, 
    -0.07443181, -0.07369612, -0.07391844, -0.07369323, -0.07482839, 
    -0.07433987, -0.07534675, -0.07940194, -0.07818765, -0.08186594, 
    -0.08416127, -0.08572227, -0.08684757, -0.08668758, -0.08638337, 
    -0.0848373, -0.0834094, -0.08233754, -0.08162832, -0.0809356, 
    -0.07887438, -0.07780544, -0.0754646, -0.07588185, -0.07517648, 
    -0.07450905, -0.07340176, -0.07358288, -0.0730991, -0.07519512, 
    -0.07379536, -0.07612054, -0.07547727, -0.08074766, -0.08285315, 
    -0.08376425, -0.08457059, -0.08656476, -0.08518257, -0.08572473, 
    -0.08444072, -0.08363488, -0.08403249, -0.08160902, -0.08254265, 
    -0.07774254, -0.07977445, -0.07458659, -0.07579604, -0.07429963, 
    -0.07505946, -0.07376226, -0.0749287, -0.07291993, -0.07248975, 
    -0.07278343, -0.07166203, -0.07499389, -0.07369606, -0.08404363, 
    -0.08397864, -0.08367661, -0.0850125, -0.08509495, -0.08633956, 
    -0.08523127, -0.08476365, -0.08358847, -0.082901, -0.08225285, 
    -0.08084576, -0.07930299, -0.07719573, -0.07571703, -0.07474191, 
    -0.07533836, -0.07481153, -0.07540069, -0.07567848, -0.07265059, 
    -0.07433529, -0.07182224, -0.07195904, -0.07308761, -0.07194361, 
    -0.08393304, -0.0843075, -0.08562057, -0.08459123, -0.08647622, 
    -0.08541583, -0.08481203, -0.08252288, -0.08202854, -0.08157262, 
    -0.08067986, -0.07954855, -0.07760258, -0.07594881, -0.07447042, 
    -0.07457776, -0.07453995, -0.07421333, -0.07502498, -0.07408093, 
    -0.07392362, -0.07433556, -0.07197738, -0.07264325, -0.07196195, 
    -0.07239471, -0.08418562, -0.08355746, -0.08389629, -0.08326024, 
    -0.08370777, -0.08173609, -0.08115415, -0.07848661, -0.07957062, 
    -0.07785264, -0.07939442, -0.07911895, -0.07779697, -0.07931036, 
    -0.07603894, -0.07824133, -0.07420066, -0.07634577, -0.07406828, 
    -0.07447676, -0.07380173, -0.07320238, -0.07245548, -0.07109739, 
    -0.07140958, -0.0702888, -0.08262987, -0.08183119, -0.08190132, 
    -0.08107325, -0.08046628, -0.07916661, -0.07712622, -0.07788721, 
    -0.07649608, -0.07621981, -0.07833566, -0.0770295, -0.08130115, 
    -0.08059496, -0.08101476, -0.0825665, -0.07771101, -0.08016554, 
    -0.07569281, -0.07697817, -0.07328752, -0.07509984, -0.071582, 
    -0.07012932, -0.06878996, -0.06725702, -0.08139875, -0.08193766, 
    -0.08097538, -0.07966264, -0.07846425, -0.07689912, -0.07674085, 
    -0.07645173, -0.07570814, -0.07508856, -0.07636044, -0.07493407, 
    -0.08043182, -0.07750163, -0.08214223, -0.08071579, -0.07973947, 
    -0.0801664, -0.07797469, -0.07746699, -0.0754381, -0.07648017, 
    -0.07048496, -0.07307626, -0.06611346, -0.0679885, -0.08212677, 
    -0.08140066, -0.07892369, -0.08009259, -0.07679583, -0.0760056, 
    -0.07536939, -0.07456377, -0.0744774, -0.07400478, -0.07478085, 
    -0.07403532, -0.07689582, -0.07560394, -0.07920305, -0.07831129, 
    -0.07872031, -0.07917135, -0.07778764, -0.07634022, -0.07630979, 
    -0.07585162, -0.07457517, -0.07678276, -0.07015704, -0.07417673, 
    -0.08061627, -0.07924915, -0.07905604, -0.07958148, -0.07608445, 
    -0.07733316, -0.07401629, -0.07489827, -0.07345873, -0.07417051, 
    -0.07427581, -0.07520163, -0.07578389, -0.07727542, -0.07851098, 
    -0.07950508, -0.07927281, -0.07818474, -0.07625262, -0.07446951, 
    -0.07485642, -0.07356714, -0.07703017, -0.07555827, -0.07612369, 
    -0.07465833, -0.07790749, -0.07513124, -0.07863358, -0.07832004, 
    -0.07735816, -0.07545934, -0.07504596, -0.07460676, -0.0748775, 
    -0.07620424, -0.07642395, -0.07738144, -0.07764784, -0.07838821, 
    -0.07900649, -0.07844135, -0.07785223, -0.07620376, -0.07474841, 
    -0.07319386, -0.07281852, -0.07105244, -0.07248651, -0.07013524, 
    -0.07212885, -0.06871345, -0.07497375, -0.07218871, -0.07731474, 
    -0.07674526, -0.07572578, -0.0734395, -0.07466515, -0.07323388, 
    -0.07643259, -0.07814737, -0.0785976, -0.07944424, -0.07857835, 
    -0.07864843, -0.07782806, -0.07809075, -0.07614964, -0.07718616, 
    -0.0742784, -0.07324512, -0.07040535, -0.06871987, -0.06704648, 
    -0.06632084, -0.06610158, -0.06601012,
  -0.06731972, -0.06577227, -0.0660704, -0.06484209, -0.06552075, 
    -0.06472041, -0.06700323, -0.0657115, -0.06653332, -0.06717907, 
    -0.06252129, -0.06478783, -0.06024929, -0.06163482, -0.05821183, 
    -0.0604628, -0.05776796, -0.05827576, -0.05676073, -0.05719081, 
    -0.05529455, -0.0565633, -0.05433598, -0.05559509, -0.05539621, 
    -0.05660561, -0.06432551, -0.06279916, -0.06441703, -0.0641969, 
    -0.06429562, -0.0655066, -0.06612515, -0.06743955, -0.06719907, 
    -0.06623466, -0.06409815, -0.06481587, -0.06302214, -0.06306212, 
    -0.06112069, -0.06198873, -0.05881266, -0.05969892, -0.0571728, 
    -0.05779811, -0.057202, -0.05738214, -0.05719966, -0.05811944, 
    -0.0577236, -0.05853945, -0.06182522, -0.06084133, -0.06382165, 
    -0.06568135, -0.06694603, -0.06785769, -0.06772807, -0.06748162, 
    -0.06622905, -0.06507218, -0.06420375, -0.06362913, -0.06306786, 
    -0.06139776, -0.06053164, -0.05863494, -0.05897303, -0.05840148, 
    -0.05786068, -0.05696348, -0.05711024, -0.05671826, -0.05841659, 
    -0.05728241, -0.05916642, -0.0586452, -0.06291559, -0.0646215, 
    -0.06535969, -0.06601297, -0.06762857, -0.06650878, -0.06694803, 
    -0.06590775, -0.06525487, -0.06557701, -0.06361348, -0.06436993, 
    -0.06048068, -0.06212704, -0.05792351, -0.05890349, -0.057691, 
    -0.05830666, -0.05725559, -0.05820071, -0.05657308, -0.05622452, 
    -0.05646248, -0.05555387, -0.05825353, -0.05720196, -0.06558603, 
    -0.06553338, -0.06528867, -0.06637099, -0.0664378, -0.06744613, 
    -0.06654824, -0.06616939, -0.06521726, -0.06466027, -0.06413513, 
    -0.06299507, -0.06174504, -0.06003762, -0.05883947, -0.05804937, 
    -0.05853265, -0.05810577, -0.05858315, -0.05880823, -0.05635485, 
    -0.05771989, -0.05568368, -0.05579452, -0.05670895, -0.05578202, 
    -0.06549644, -0.06579982, -0.06686363, -0.06602969, -0.06755684, 
    -0.06669776, -0.06620858, -0.06435392, -0.06395339, -0.063584, 
    -0.06286065, -0.061944, -0.06036728, -0.05902728, -0.05782939, 
    -0.05791636, -0.05788573, -0.05762107, -0.05827872, -0.0575138, 
    -0.05738633, -0.05772012, -0.05580938, -0.0563489, -0.05579688, 
    -0.05614753, -0.06570107, -0.06519213, -0.06546666, -0.06495133, 
    -0.06531393, -0.06371644, -0.06324495, -0.06108357, -0.06196189, 
    -0.06056988, -0.06181912, -0.06159592, -0.06052478, -0.06175101, 
    -0.05910031, -0.06088483, -0.05761081, -0.05934892, -0.05750354, 
    -0.05783452, -0.05728757, -0.05680194, -0.05619676, -0.05509638, 
    -0.05534933, -0.05444123, -0.06444059, -0.0637935, -0.06385031, 
    -0.06317939, -0.0626876, -0.06163454, -0.05998129, -0.06059789, 
    -0.05947071, -0.05924686, -0.06096126, -0.05990292, -0.06336404, 
    -0.06279185, -0.063132, -0.06438926, -0.06045513, -0.06244392, 
    -0.05881985, -0.05986134, -0.05687093, -0.05833939, -0.05548903, 
    -0.05431202, -0.05322686, -0.05198491, -0.06344312, -0.06387976, 
    -0.06310008, -0.06203645, -0.06106545, -0.05979728, -0.05966904, 
    -0.05943478, -0.05883227, -0.05833025, -0.05936081, -0.05820506, 
    -0.06265968, -0.06028548, -0.0640455, -0.06288976, -0.06209871, 
    -0.06244462, -0.06066878, -0.06025741, -0.05861346, -0.05945782, 
    -0.05460017, -0.05669975, -0.05105847, -0.05257753, -0.06403298, 
    -0.06344467, -0.06143772, -0.06238481, -0.05971359, -0.0590733, 
    -0.05855779, -0.05790503, -0.05783505, -0.0574521, -0.05808092, 
    -0.05747684, -0.05979461, -0.05874784, -0.06166407, -0.06094152, 
    -0.06127292, -0.06163839, -0.06051722, -0.05934442, -0.05931976, 
    -0.05894853, -0.05791427, -0.059703, -0.05433448, -0.05759142, 
    -0.06280913, -0.06170142, -0.06154495, -0.06197069, -0.05913718, 
    -0.06014897, -0.05746142, -0.05817606, -0.05700965, -0.05758638, 
    -0.0576717, -0.05842186, -0.05889364, -0.06010218, -0.06110331, 
    -0.06190878, -0.06172059, -0.06083897, -0.05927344, -0.05782865, 
    -0.05814216, -0.05709749, -0.05990347, -0.05871083, -0.05916898, 
    -0.05798164, -0.06061433, -0.05836483, -0.06120266, -0.0609486, 
    -0.06016922, -0.05863068, -0.05829572, -0.05793986, -0.05815923, 
    -0.05923424, -0.05941227, -0.06018809, -0.06040395, -0.06100384, 
    -0.0615048, -0.06104689, -0.06056955, -0.05923385, -0.05805463, 
    -0.05679503, -0.05649091, -0.05505996, -0.05622191, -0.05431683, 
    -0.05593212, -0.05316487, -0.05823722, -0.05598062, -0.06013404, 
    -0.05967261, -0.05884656, -0.05699407, -0.05798717, -0.05682747, 
    -0.05941926, -0.06080869, -0.06117349, -0.06185949, -0.0611579, 
    -0.06121468, -0.06054997, -0.06076282, -0.05919, -0.06002986, -0.0576738, 
    -0.05683658, -0.05453567, -0.05317008, -0.05181434, -0.05122647, 
    -0.05104885, -0.05097476,
  -0.06391447, -0.06222167, -0.06254755, -0.06120564, -0.06194681, 
    -0.06107282, -0.06356799, -0.06215525, -0.06305381, -0.06376047, 
    -0.05867587, -0.06114641, -0.05620678, -0.0577116, -0.0539992, 
    -0.05643849, -0.05351913, -0.05406837, -0.05243094, -0.05289539, 
    -0.05084988, -0.05221782, -0.04981819, -0.05117367, -0.05095939, 
    -0.05226349, -0.06064191, -0.05897837, -0.06074176, -0.06050161, 
    -0.06060929, -0.06193136, -0.06260741, -0.06404569, -0.06378238, 
    -0.06272715, -0.0603939, -0.06117702, -0.05922118, -0.05926472, 
    -0.05715287, -0.05809643, -0.05464952, -0.05560982, -0.05287593, 
    -0.05355173, -0.05290747, -0.0531021, -0.05290494, -0.05389925, 
    -0.05347117, -0.05435374, -0.05791861, -0.05684945, -0.06009239, 
    -0.0621223, -0.06350539, -0.0645037, -0.0643617, -0.06409176, 
    -0.06272102, -0.06145686, -0.06050908, -0.05988252, -0.05927098, 
    -0.05745393, -0.05651321, -0.0544571, -0.0548232, -0.05420442, 
    -0.05361939, -0.05264986, -0.05280836, -0.05238508, -0.05422076, 
    -0.05299434, -0.0550327, -0.05446822, -0.05910514, -0.06096487, 
    -0.06177086, -0.06248477, -0.0642527, -0.06302696, -0.06350757, 
    -0.06236975, -0.06165637, -0.06200828, -0.05986547, -0.06069036, 
    -0.05645789, -0.05824688, -0.05368733, -0.05474789, -0.05343593, 
    -0.05410181, -0.05296537, -0.05398717, -0.05222838, -0.0518523, 
    -0.05210903, -0.05112926, -0.05404432, -0.05290742, -0.06201814, 
    -0.06196061, -0.06169329, -0.06287625, -0.06294932, -0.06405289, 
    -0.06307013, -0.06265578, -0.0616153, -0.06100719, -0.06043423, 
    -0.05919169, -0.05783143, -0.05597714, -0.05467856, -0.05382345, 
    -0.05434638, -0.05388446, -0.05440104, -0.05464473, -0.0519929, 
    -0.05346717, -0.05126915, -0.05138862, -0.05237504, -0.05137515, 
    -0.06192025, -0.06225177, -0.06341521, -0.06250305, -0.06417414, 
    -0.0632337, -0.06269864, -0.06067289, -0.06023603, -0.05983333, 
    -0.05904532, -0.05804779, -0.05633481, -0.05488197, -0.05358555, 
    -0.0536796, -0.05364647, -0.05336033, -0.05407158, -0.05324438, 
    -0.05310663, -0.0534674, -0.05140464, -0.05198648, -0.05139116, 
    -0.05176925, -0.06214385, -0.06158786, -0.06188772, -0.06132491, 
    -0.06172087, -0.0599777, -0.05946387, -0.05711254, -0.05806725, 
    -0.05655472, -0.05791198, -0.05766932, -0.05650576, -0.05783793, 
    -0.05496107, -0.05689669, -0.05334923, -0.05523045, -0.0532333, 
    -0.0535911, -0.05299992, -0.05247543, -0.05182235, -0.05063646, 
    -0.05090889, -0.04993139, -0.06076746, -0.0600617, -0.06012364, 
    -0.05939246, -0.0588569, -0.05771129, -0.05591604, -0.05658513, 
    -0.05536243, -0.05511985, -0.05697969, -0.05583104, -0.05959363, 
    -0.05897041, -0.05934083, -0.06071145, -0.05643016, -0.05859167, 
    -0.05465731, -0.05578594, -0.05254991, -0.05413722, -0.0510594, 
    -0.04979242, -0.04862646, -0.04729465, -0.0596798, -0.06015574, 
    -0.05930608, -0.05814834, -0.05709287, -0.05571648, -0.05557742, 
    -0.05532349, -0.05467076, -0.05412732, -0.05524332, -0.05399187, 
    -0.05882651, -0.05624605, -0.06033648, -0.05907702, -0.05821606, 
    -0.05859243, -0.05666208, -0.05621559, -0.05443386, -0.05534846, 
    -0.05010237, -0.05236511, -0.04630303, -0.0479298, -0.06032282, 
    -0.05968149, -0.05749736, -0.05852734, -0.05562573, -0.05493181, 
    -0.05437359, -0.05366734, -0.05359167, -0.0531777, -0.05385758, 
    -0.05320444, -0.05571358, -0.05457934, -0.0577434, -0.05695825, 
    -0.05731827, -0.05771548, -0.05649755, -0.05522557, -0.05519884, 
    -0.05479667, -0.05367734, -0.05561425, -0.04981658, -0.05332828, 
    -0.05898922, -0.05778401, -0.05761391, -0.05807681, -0.05500102, 
    -0.05609794, -0.05318778, -0.0539605, -0.05269971, -0.05332283, 
    -0.05341506, -0.05422647, -0.05473723, -0.05604718, -0.05713399, 
    -0.05800949, -0.05780485, -0.05684688, -0.05514865, -0.05358475, 
    -0.05392382, -0.05279458, -0.05583163, -0.05453927, -0.05503546, 
    -0.05375019, -0.05660297, -0.05416476, -0.05724192, -0.05696595, 
    -0.05611991, -0.05445249, -0.05408997, -0.05370501, -0.05394229, 
    -0.05510618, -0.05529909, -0.05614038, -0.05637461, -0.05702594, 
    -0.05757027, -0.05707271, -0.05655436, -0.05510575, -0.05382914, 
    -0.05246797, -0.05213971, -0.05059725, -0.05184948, -0.04979759, 
    -0.05153696, -0.04855993, -0.05402667, -0.05158925, -0.05608174, 
    -0.0555813, -0.05468624, -0.05268289, -0.05375617, -0.05250299, 
    -0.05530667, -0.056814, -0.05721024, -0.05795588, -0.05719329, 
    -0.05725498, -0.0565331, -0.05676418, -0.05505824, -0.05596872, 
    -0.05341733, -0.05251282, -0.05003298, -0.04856551, -0.04711195, 
    -0.04648273, -0.04629274, -0.04621351,
  -0.04035198, -0.03907359, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009016, -0.03902347, -0.03970177, -0.0402356, 
    -0.03640241, -0.03826259, -0.03454811, -0.03567765, -0.03289467, 
    -0.03472191, -0.0325357, -0.03294641, -0.03172283, -0.03206963, 
    -0.03054395, -0.03156378, -0.02977613, -0.03078516, -0.03062552, 
    -0.03159786, -0.03788236, -0.03662992, -0.0379576, -0.03777665, 
    -0.03785779, -0.03885455, -0.03936473, -0.04045115, -0.04025215, 
    -0.03945512, -0.03769551, -0.03828567, -0.0368126, -0.03684536, 
    -0.03525804, -0.0359668, -0.03338129, -0.03410057, -0.03205509, 
    -0.03256006, -0.03207865, -0.03222404, -0.03207676, -0.03281991, 
    -0.03249985, -0.03315991, -0.03583318, -0.03503027, -0.03746841, 
    -0.03899861, -0.04004287, -0.0407974, -0.04069003, -0.04048597, 
    -0.0394505, -0.03849666, -0.03778228, -0.03731038, -0.03685007, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351131, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306041, 
    -0.03214354, -0.03366819, -0.03324559, -0.03672529, -0.03812575, 
    -0.03873348, -0.03927216, -0.04060763, -0.0396815, -0.04004452, 
    -0.03918534, -0.03864712, -0.03891259, -0.03729754, -0.03791887, 
    -0.03473647, -0.03607988, -0.03266144, -0.03345493, -0.0324735, 
    -0.03297142, -0.0321219, -0.03288567, -0.03157166, -0.03129108, 
    -0.0314826, -0.03075207, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887662, -0.03867497, -0.0395677, -0.03962287, -0.04045659, 
    -0.0397141, -0.03940124, -0.03861614, -0.03815764, -0.03772589, 
    -0.03679041, -0.03576767, -0.03437591, -0.03340303, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319531, -0.03337771, -0.03139596, 
    -0.03249685, -0.03085631, -0.03094536, -0.03168111, -0.03093531, 
    -0.03884617, -0.03909631, -0.03997475, -0.03928595, -0.04054824, 
    -0.03983764, -0.0394336, -0.03790571, -0.0375766, -0.03727334, 
    -0.03668029, -0.03593025, -0.03464414, -0.03355532, -0.03258535, 
    -0.03265566, -0.03263089, -0.032417, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249703, -0.03095729, -0.03139117, -0.03094725, 
    -0.03122914, -0.03901487, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869577, -0.03738204, -0.03699523, -0.03522776, -0.03594487, 
    -0.03480911, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240871, -0.03381631, -0.03232207, 
    -0.0325895, -0.03214771, -0.03175604, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797697, -0.0374453, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567741, -0.03433011, -0.03483192, 
    -0.03391519, -0.03373347, -0.03512803, -0.03426639, -0.0370929, 
    -0.03662394, -0.03690264, -0.03793476, -0.03471566, -0.03633909, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299791, -0.03070002, 
    -0.02975696, -0.02889069, -0.02790317, -0.03715776, -0.03751612, 
    -0.03687648, -0.03600582, -0.03521299, -0.03418051, -0.03407629, 
    -0.03388602, -0.03339719, -0.03299051, -0.03382596, -0.03288919, 
    -0.0365157, -0.03457757, -0.03765226, -0.03670414, -0.03605671, 
    -0.03633966, -0.03488967, -0.03455472, -0.03321987, -0.03390472, 
    -0.02998751, -0.0316737, -0.02716934, -0.02837385, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629072, -0.03411249, -0.03359264, 
    -0.03317476, -0.0326465, -0.03258992, -0.03228053, -0.03278875, 
    -0.03230051, -0.03417834, -0.03332876, -0.03570153, -0.03511194, 
    -0.03538223, -0.03568055, -0.03476622, -0.03381266, -0.03379264, 
    -0.03349145, -0.03265397, -0.03410389, -0.02977493, -0.03239306, 
    -0.03663808, -0.03573204, -0.03560426, -0.03595205, -0.03364447, 
    -0.03446649, -0.03228806, -0.03286572, -0.03192349, -0.03238898, 
    -0.03245791, -0.03306468, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199434, -0.03426683, -0.03329876, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301851, -0.0353249, -0.03511771, 
    -0.03448297, -0.03323382, -0.03296256, -0.03267466, -0.0328521, 
    -0.03372323, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480884, -0.03372291, -0.03276749, 
    -0.03175048, -0.03150549, -0.03035583, -0.03128898, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.03407919, -0.03340878, -0.03191093, -0.03271292, -0.03177662, 
    -0.03387342, -0.03500367, -0.03530111, -0.03586118, -0.03528839, 
    -0.0353347, -0.03479289, -0.03496628, -0.03368732, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993588, -0.02884545, -0.02776788, 
    -0.02730223, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.0189572, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277074, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459348, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927695, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  296.7043, 297.9638, 297.7187, 298.7369, 298.1718, 298.839, 296.9594, 
    298.0138, 297.3404, 296.8176, 300.7122, 298.7824, 302.7232, 301.4879, 
    304.599, 302.5305, 305.0127, 304.5395, 305.9586, 305.5526, 307.3677, 
    306.1461, 308.3125, 307.0758, 307.2689, 306.1058, 299.1718, 300.4719, 
    299.0945, 299.2805, 299.1971, 298.1834, 297.6734, 296.6083, 296.8015, 
    297.584, 299.3642, 298.7592, 300.2814, 300.2471, 301.9428, 301.1773, 
    304.0388, 303.2234, 305.5696, 304.9851, 305.5421, 305.3731, 305.5443, 
    304.6862, 305.0543, 304.293, 301.3205, 302.1916, 299.5991, 298.0383, 
    297.0055, 296.2741, 296.3775, 296.5744, 297.5886, 298.5448, 299.275, 
    299.7627, 300.2421, 301.6963, 302.4688, 304.2037, 303.8903, 304.4216, 
    304.927, 305.7667, 305.6284, 305.9987, 304.4077, 305.4663, 303.7119, 
    304.1945, 300.3715, 298.9223, 298.3048, 297.7658, 296.4569, 297.3602, 
    297.0038, 297.8525, 298.3925, 298.1254, 299.7759, 299.1344, 302.5147, 
    301.0562, 304.8687, 303.9547, 305.0847, 304.5107, 305.4916, 304.61, 
    306.1367, 306.4692, 306.2419, 307.1161, 304.5604, 305.5419, 298.1179, 
    298.1614, 298.3645, 297.4726, 297.4181, 296.603, 297.3283, 297.6375, 
    298.424, 298.8897, 299.3331, 300.3045, 301.3907, 302.915, 304.0139, 
    304.7522, 304.2995, 304.6992, 304.2523, 304.0431, 306.3445, 305.0576, 
    306.9902, 306.8831, 306.0074, 306.8952, 298.192, 297.9414, 297.0722, 
    297.7523, 296.5143, 297.2066, 297.6052, 299.1476, 299.4875, 299.8009, 
    300.4203, 301.2164, 302.617, 303.8399, 304.9561, 304.8755, 304.9038, 
    305.1498, 304.5368, 305.2499, 305.369, 305.0576, 306.8687, 306.3505, 
    306.8808, 306.5433, 298.0229, 298.4448, 298.2167, 298.6457, 298.3434, 
    299.688, 300.0898, 301.9754, 301.2007, 302.4347, 301.3259, 301.5221, 
    302.4746, 301.3858, 303.7722, 302.1523, 305.1594, 303.543, 305.2595, 
    304.9514, 305.4618, 305.9194, 306.496, 307.562, 307.3149, 308.2081, 
    299.0747, 299.6229, 299.575, 300.1464, 300.5695, 301.4883, 302.9663, 
    302.4099, 303.4322, 303.6376, 302.0849, 303.0374, 299.9883, 300.4791, 
    300.1869, 299.1179, 302.5378, 300.7802, 304.0321, 303.0754, 305.8541, 
    304.4796, 307.1789, 308.3359, 309.4288, 310.7087, 299.9209, 299.5501, 
    300.2145, 301.1352, 301.9919, 303.1336, 303.2507, 303.465, 304.0208, 
    304.4886, 303.5326, 304.6059, 300.5926, 302.6908, 299.4091, 300.3946, 
    301.0809, 300.7799, 302.3464, 302.7165, 304.2238, 303.444, 308.0498, 
    306.0158, 311.6866, 310.0937, 299.4199, 299.9197, 301.6616, 300.8319, 
    303.2101, 303.7976, 304.276, 304.8857, 304.9508, 305.3075, 304.7226, 
    305.2845, 303.136, 304.099, 301.4624, 302.1024, 301.8079, 301.485, 
    302.4824, 303.5475, 303.5706, 303.9128, 304.8756, 303.2197, 308.3125, 
    305.176, 300.4647, 301.4289, 301.5672, 301.1932, 303.7386, 302.8144, 
    305.2989, 304.6331, 305.7232, 305.1822, 305.1027, 304.4029, 303.9637, 
    302.8566, 301.9582, 301.2475, 301.4126, 302.1938, 303.6129, 304.9566, 
    304.6647, 305.6404, 303.0371, 304.1332, 303.7091, 304.8149, 302.3951, 
    304.4547, 301.8702, 302.0962, 302.7961, 304.2075, 304.5209, 304.8534, 
    304.649, 303.649, 303.4856, 302.7791, 302.5841, 302.047, 301.6028, 
    302.0085, 302.4351, 303.6496, 304.747, 305.9258, 306.215, 307.5968, 
    306.4711, 308.33, 306.7484, 309.4906, 304.5749, 306.7026, 302.828, 
    303.2475, 304.007, 305.7372, 304.8098, 305.8948, 303.4792, 302.2206, 
    301.8961, 301.2906, 301.9099, 301.8595, 302.453, 302.2622, 303.69, 
    302.9224, 305.1006, 305.8864, 308.1143, 309.4861, 310.8879, 311.5081, 
    311.6971, 311.7762 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.356892e-08, 6.384848e-08, 6.379413e-08, 6.401962e-08, 6.389453e-08, 
    6.404218e-08, 6.362559e-08, 6.385958e-08, 6.37102e-08, 6.359408e-08, 
    6.445721e-08, 6.402967e-08, 6.490126e-08, 6.462861e-08, 6.531352e-08, 
    6.485884e-08, 6.54052e-08, 6.530039e-08, 6.561581e-08, 6.552545e-08, 
    6.592889e-08, 6.565751e-08, 6.613801e-08, 6.586408e-08, 6.590693e-08, 
    6.564856e-08, 6.41157e-08, 6.440398e-08, 6.409863e-08, 6.413973e-08, 
    6.412129e-08, 6.389712e-08, 6.378416e-08, 6.354755e-08, 6.35905e-08, 
    6.376428e-08, 6.415822e-08, 6.402449e-08, 6.436151e-08, 6.43539e-08, 
    6.472909e-08, 6.455993e-08, 6.519053e-08, 6.50113e-08, 6.552921e-08, 
    6.539896e-08, 6.55231e-08, 6.548546e-08, 6.552359e-08, 6.533256e-08, 
    6.541441e-08, 6.524632e-08, 6.459161e-08, 6.478403e-08, 6.421014e-08, 
    6.386507e-08, 6.363586e-08, 6.347321e-08, 6.34962e-08, 6.354004e-08, 
    6.37653e-08, 6.397708e-08, 6.413847e-08, 6.424643e-08, 6.43528e-08, 
    6.46748e-08, 6.484521e-08, 6.522678e-08, 6.515791e-08, 6.527457e-08, 
    6.538601e-08, 6.557312e-08, 6.554232e-08, 6.562475e-08, 6.527149e-08, 
    6.550627e-08, 6.511868e-08, 6.522469e-08, 6.438174e-08, 6.406056e-08, 
    6.392407e-08, 6.380458e-08, 6.351388e-08, 6.371463e-08, 6.36355e-08, 
    6.382376e-08, 6.394339e-08, 6.388422e-08, 6.424938e-08, 6.410742e-08, 
    6.485531e-08, 6.453317e-08, 6.537302e-08, 6.517205e-08, 6.542118e-08, 
    6.529405e-08, 6.551188e-08, 6.531584e-08, 6.565543e-08, 6.572938e-08, 
    6.567885e-08, 6.587296e-08, 6.530497e-08, 6.55231e-08, 6.388257e-08, 
    6.389222e-08, 6.393717e-08, 6.373956e-08, 6.372747e-08, 6.354637e-08, 
    6.370751e-08, 6.377613e-08, 6.395032e-08, 6.405336e-08, 6.415131e-08, 
    6.436666e-08, 6.460716e-08, 6.494347e-08, 6.518507e-08, 6.534702e-08, 
    6.524771e-08, 6.533539e-08, 6.523738e-08, 6.519144e-08, 6.570168e-08, 
    6.541517e-08, 6.584504e-08, 6.582125e-08, 6.562671e-08, 6.582393e-08, 
    6.389899e-08, 6.384346e-08, 6.365067e-08, 6.380154e-08, 6.352665e-08, 
    6.368052e-08, 6.376901e-08, 6.411039e-08, 6.418539e-08, 6.425494e-08, 
    6.43923e-08, 6.456858e-08, 6.487782e-08, 6.514688e-08, 6.539249e-08, 
    6.537449e-08, 6.538083e-08, 6.54357e-08, 6.529979e-08, 6.545802e-08, 
    6.548457e-08, 6.541514e-08, 6.581807e-08, 6.570296e-08, 6.582075e-08, 
    6.574579e-08, 6.386151e-08, 6.395495e-08, 6.390446e-08, 6.39994e-08, 
    6.393252e-08, 6.422994e-08, 6.431911e-08, 6.473636e-08, 6.456511e-08, 
    6.483764e-08, 6.45928e-08, 6.463618e-08, 6.484655e-08, 6.460603e-08, 
    6.513206e-08, 6.477543e-08, 6.543784e-08, 6.508173e-08, 6.546015e-08, 
    6.539143e-08, 6.55052e-08, 6.560711e-08, 6.573531e-08, 6.597185e-08, 
    6.591708e-08, 6.611489e-08, 6.409424e-08, 6.421543e-08, 6.420476e-08, 
    6.433159e-08, 6.442539e-08, 6.462868e-08, 6.495473e-08, 6.483211e-08, 
    6.505721e-08, 6.51024e-08, 6.476043e-08, 6.497039e-08, 6.429654e-08, 
    6.440542e-08, 6.434059e-08, 6.41038e-08, 6.486038e-08, 6.447211e-08, 
    6.518906e-08, 6.497873e-08, 6.559258e-08, 6.528731e-08, 6.588692e-08, 
    6.614327e-08, 6.638449e-08, 6.666644e-08, 6.428157e-08, 6.419923e-08, 
    6.434667e-08, 6.455067e-08, 6.473994e-08, 6.499156e-08, 6.50173e-08, 
    6.506445e-08, 6.518654e-08, 6.528921e-08, 6.507936e-08, 6.531494e-08, 
    6.443068e-08, 6.489408e-08, 6.41681e-08, 6.438672e-08, 6.453865e-08, 
    6.447199e-08, 6.48181e-08, 6.489968e-08, 6.523117e-08, 6.505981e-08, 
    6.608001e-08, 6.562864e-08, 6.688109e-08, 6.653109e-08, 6.417046e-08, 
    6.428129e-08, 6.466703e-08, 6.448349e-08, 6.500836e-08, 6.513755e-08, 
    6.524257e-08, 6.537682e-08, 6.539132e-08, 6.547086e-08, 6.534052e-08, 
    6.546571e-08, 6.49921e-08, 6.520374e-08, 6.462293e-08, 6.47643e-08, 
    6.469926e-08, 6.462793e-08, 6.484809e-08, 6.508266e-08, 6.508766e-08, 
    6.516288e-08, 6.537484e-08, 6.501048e-08, 6.613828e-08, 6.54418e-08, 
    6.440214e-08, 6.461564e-08, 6.464612e-08, 6.456342e-08, 6.51246e-08, 
    6.492127e-08, 6.546892e-08, 6.532091e-08, 6.556343e-08, 6.544292e-08, 
    6.542518e-08, 6.527041e-08, 6.517404e-08, 6.493059e-08, 6.47325e-08, 
    6.457542e-08, 6.461194e-08, 6.478449e-08, 6.509701e-08, 6.539263e-08, 
    6.532787e-08, 6.5545e-08, 6.49703e-08, 6.521128e-08, 6.511815e-08, 
    6.5361e-08, 6.482886e-08, 6.528204e-08, 6.471303e-08, 6.476292e-08, 
    6.491723e-08, 6.522764e-08, 6.52963e-08, 6.536963e-08, 6.532438e-08, 
    6.510494e-08, 6.506898e-08, 6.491348e-08, 6.487055e-08, 6.475205e-08, 
    6.465395e-08, 6.474359e-08, 6.483771e-08, 6.510503e-08, 6.534592e-08, 
    6.560856e-08, 6.567284e-08, 6.597972e-08, 6.572991e-08, 6.614216e-08, 
    6.579169e-08, 6.639835e-08, 6.530828e-08, 6.578136e-08, 6.492425e-08, 
    6.501659e-08, 6.518361e-08, 6.556667e-08, 6.535986e-08, 6.560172e-08, 
    6.506757e-08, 6.479046e-08, 6.471874e-08, 6.458497e-08, 6.47218e-08, 
    6.471067e-08, 6.484161e-08, 6.479953e-08, 6.51139e-08, 6.494503e-08, 
    6.542474e-08, 6.55998e-08, 6.609416e-08, 6.639722e-08, 6.67057e-08, 
    6.684189e-08, 6.688335e-08, 6.690068e-08 ;

 SOM_C_LEACHED =
  6.799576e-20, 5.784397e-21, 3.186314e-20, 3.781883e-20, 1.091324e-20, 
    1.352854e-20, -7.690232e-21, -2.716396e-20, 3.505336e-20, -2.381964e-20, 
    2.362712e-20, 3.420565e-20, -3.124232e-21, -1.062299e-20, 3.461862e-20, 
    2.621248e-20, 6.352486e-20, 2.816233e-20, -8.239468e-20, 4.558226e-20, 
    -1.036748e-20, -2.228872e-21, 7.602613e-20, 1.834276e-20, 1.831154e-20, 
    -3.353828e-20, -1.264245e-20, 5.340808e-20, 3.135758e-20, -3.589461e-20, 
    -3.177138e-20, 2.63052e-20, 1.005138e-19, -6.687746e-21, -4.955645e-21, 
    -6.218095e-21, 5.259001e-20, -3.429285e-20, 3.268283e-20, -3.905691e-20, 
    2.633893e-20, 4.025091e-20, 8.729365e-21, 1.975519e-20, -1.439565e-20, 
    4.010447e-21, 7.13598e-20, -3.989678e-21, 3.487805e-20, 5.978779e-20, 
    1.929251e-20, -1.964346e-20, -3.946242e-21, 4.120298e-20, 1.816417e-20, 
    1.335093e-20, 6.995167e-21, -2.471493e-21, -5.189719e-20, 6.365055e-21, 
    -7.024981e-20, 3.540338e-20, 2.300081e-22, 5.436196e-20, 1.956477e-20, 
    -9.099482e-21, -5.643635e-20, 3.625111e-20, -4.479015e-20, -7.77256e-20, 
    1.593235e-21, -2.195422e-20, -4.714119e-20, -1.939608e-20, -2.783546e-21, 
    1.600512e-20, -1.214802e-20, 3.19964e-20, -7.950964e-21, 1.287464e-20, 
    -5.226228e-20, 3.526865e-20, 8.712128e-21, -3.357215e-20, -1.611282e-20, 
    -6.596757e-20, -1.666533e-20, -2.213702e-20, -3.826636e-20, 2.620029e-20, 
    -2.070008e-20, -4.134382e-21, -3.725858e-20, 1.257159e-20, -3.566785e-20, 
    6.983666e-21, 3.532867e-21, 1.902074e-20, 4.515321e-20, -2.774799e-20, 
    8.861884e-20, -5.125841e-20, -2.26976e-20, -3.887951e-20, 4.939567e-20, 
    6.898462e-20, -1.131881e-20, -1.027744e-21, 8.024647e-21, -4.908806e-20, 
    -6.990703e-20, 4.090592e-20, 2.088447e-20, -1.680522e-20, -3.662338e-20, 
    2.796942e-20, 2.947277e-20, -2.280889e-20, 3.155092e-21, -6.076785e-20, 
    -7.228953e-20, 7.197974e-20, 1.228787e-20, -4.516528e-20, 2.728294e-21, 
    -6.414388e-20, 1.891423e-20, 1.824324e-20, 2.120318e-20, 8.134926e-20, 
    4.133611e-20, -5.529981e-21, 4.302102e-20, 5.952275e-20, -9.267587e-20, 
    -6.421909e-20, 2.476901e-20, 1.856488e-21, -2.468964e-20, 2.936265e-20, 
    -8.057199e-21, -2.624529e-20, 8.253718e-20, 3.695357e-20, -1.602048e-20, 
    5.053847e-20, -6.271269e-20, 3.020451e-20, -1.103285e-19, -6.802025e-22, 
    5.223765e-20, -9.8812e-20, 5.684968e-20, -7.618499e-20, 2.924768e-21, 
    -2.133959e-20, 3.337591e-20, -6.694773e-21, 3.141091e-21, -9.313816e-20, 
    -7.715976e-20, -3.503665e-20, -1.129557e-20, -2.170056e-20, 
    -3.676581e-20, -4.767825e-20, 5.650884e-20, 1.126752e-21, 6.258447e-20, 
    -1.853261e-20, -1.017641e-19, -2.915833e-20, -3.159542e-20, 1.484597e-20, 
    -4.352514e-20, 5.582953e-22, 4.247375e-21, 1.645368e-20, 2.279192e-21, 
    -4.669785e-20, 3.675786e-20, -3.243836e-20, -8.600927e-21, 1.45277e-20, 
    8.41596e-21, -3.965254e-20, -5.450335e-20, -9.490375e-21, 2.84381e-20, 
    1.176646e-20, 5.429896e-21, -4.306028e-20, -4.744816e-20, -1.192768e-20, 
    -5.002558e-20, 2.651737e-20, 1.183728e-20, -1.266107e-20, 3.845591e-21, 
    5.601912e-20, 2.560926e-20, 1.74259e-20, 3.809755e-20, -3.703054e-20, 
    -3.668875e-20, 7.617168e-20, -4.996352e-20, -5.427616e-20, 6.139945e-20, 
    1.142535e-20, -3.394475e-20, -2.080552e-20, 1.348559e-20, -1.813312e-20, 
    -1.580827e-20, 4.670637e-20, -3.25e-20, -6.747299e-21, -6.909917e-20, 
    6.12812e-21, -1.499891e-20, 5.188069e-21, 6.131123e-20, -1.290714e-20, 
    -9.744207e-21, 3.136244e-20, -1.354973e-20, -7.246205e-20, 6.917312e-20, 
    -1.600377e-21, 6.937805e-20, 3.27791e-20, -6.976646e-20, -4.284513e-21, 
    1.560695e-20, -1.703907e-20, -3.586714e-20, -4.512048e-20, 2.766592e-20, 
    -1.382688e-20, 2.225857e-20, -2.184671e-20, -6.322792e-20, 6.399402e-20, 
    2.489947e-20, -1.2256e-20, 5.022241e-20, 7.805675e-21, 3.604211e-20, 
    1.670381e-20, -3.65866e-20, 3.576515e-20, 1.423109e-21, -6.275372e-20, 
    6.01423e-20, 2.199157e-20, -1.666886e-20, 2.250698e-20, -4.93124e-20, 
    -5.78286e-20, 5.397531e-20, -2.120425e-20, 1.057796e-19, -1.030961e-20, 
    -3.201191e-20, -5.228104e-20, -2.261494e-20, -3.150349e-20, 
    -4.817497e-20, 4.39983e-20, -3.219313e-20, -7.579922e-21, 2.267422e-20, 
    -3.933052e-20, -2.880951e-20, 8.350128e-21, 3.256275e-20, 1.720735e-20, 
    8.123509e-20, 2.090567e-20, -3.019495e-21, -1.323248e-20, 9.544815e-21, 
    1.664707e-20, -5.345702e-21, 7.959429e-21, 4.145767e-20, 9.073537e-21, 
    -6.200361e-21, -2.527503e-20, 3.849913e-20, 4.675566e-20, 5.589579e-21, 
    4.01394e-21, 5.504844e-21, -9.584341e-21, 4.72683e-20, -2.414454e-22, 
    3.552849e-20, -2.021971e-20, -1.248271e-20, -3.249854e-20, -9.656761e-21, 
    -3.888912e-20, -2.146107e-20, -7.872717e-21, 5.177226e-21, -8.563564e-21, 
    3.491871e-20, 1.983495e-20, 3.941384e-20, 5.759656e-21, 2.349276e-20, 
    6.644998e-21, 1.467352e-20, -1.537464e-20, 4.163038e-20, -4.412623e-20, 
    -5.207517e-21, 3.300052e-20, 2.419371e-20, -4.560378e-20, 1.971595e-21, 
    4.840245e-20, 3.095534e-20, -4.106729e-21, -2.902547e-20, -5.048131e-20, 
    -4.815284e-20, -3.651929e-20, -4.511208e-20, -5.828621e-20, 3.376665e-20, 
    4.429075e-20, -4.487058e-22, -3.448296e-20, -4.42431e-20, -6.731025e-20 ;

 SR =
  6.356978e-08, 6.384934e-08, 6.379499e-08, 6.402048e-08, 6.389539e-08, 
    6.404304e-08, 6.362645e-08, 6.386044e-08, 6.371106e-08, 6.359494e-08, 
    6.445807e-08, 6.403054e-08, 6.490213e-08, 6.462948e-08, 6.531439e-08, 
    6.485971e-08, 6.540607e-08, 6.530126e-08, 6.561668e-08, 6.552632e-08, 
    6.592977e-08, 6.565838e-08, 6.61389e-08, 6.586495e-08, 6.590781e-08, 
    6.564943e-08, 6.411657e-08, 6.440485e-08, 6.409949e-08, 6.41406e-08, 
    6.412215e-08, 6.389798e-08, 6.378502e-08, 6.354841e-08, 6.359136e-08, 
    6.376514e-08, 6.415908e-08, 6.402535e-08, 6.436237e-08, 6.435476e-08, 
    6.472996e-08, 6.456079e-08, 6.51914e-08, 6.501217e-08, 6.553009e-08, 
    6.539984e-08, 6.552398e-08, 6.548633e-08, 6.552447e-08, 6.533344e-08, 
    6.541529e-08, 6.524719e-08, 6.459248e-08, 6.478489e-08, 6.421101e-08, 
    6.386593e-08, 6.363672e-08, 6.347406e-08, 6.349706e-08, 6.35409e-08, 
    6.376616e-08, 6.397794e-08, 6.413933e-08, 6.42473e-08, 6.435366e-08, 
    6.467567e-08, 6.484608e-08, 6.522765e-08, 6.515878e-08, 6.527544e-08, 
    6.538689e-08, 6.557399e-08, 6.55432e-08, 6.562563e-08, 6.527236e-08, 
    6.550714e-08, 6.511956e-08, 6.522556e-08, 6.438261e-08, 6.406143e-08, 
    6.392494e-08, 6.380544e-08, 6.351474e-08, 6.371549e-08, 6.363636e-08, 
    6.382462e-08, 6.394425e-08, 6.388508e-08, 6.425024e-08, 6.410828e-08, 
    6.485618e-08, 6.453404e-08, 6.537388e-08, 6.517291e-08, 6.542206e-08, 
    6.529492e-08, 6.551276e-08, 6.53167e-08, 6.565631e-08, 6.573026e-08, 
    6.567973e-08, 6.587384e-08, 6.530584e-08, 6.552398e-08, 6.388343e-08, 
    6.389308e-08, 6.393803e-08, 6.374042e-08, 6.372833e-08, 6.354723e-08, 
    6.370837e-08, 6.377699e-08, 6.395118e-08, 6.405422e-08, 6.415217e-08, 
    6.436752e-08, 6.460803e-08, 6.494434e-08, 6.518594e-08, 6.53479e-08, 
    6.524859e-08, 6.533626e-08, 6.523825e-08, 6.519231e-08, 6.570255e-08, 
    6.541605e-08, 6.584592e-08, 6.582213e-08, 6.562759e-08, 6.582481e-08, 
    6.389985e-08, 6.384432e-08, 6.365153e-08, 6.38024e-08, 6.352751e-08, 
    6.368138e-08, 6.376987e-08, 6.411125e-08, 6.418625e-08, 6.425581e-08, 
    6.439316e-08, 6.456945e-08, 6.487869e-08, 6.514775e-08, 6.539337e-08, 
    6.537537e-08, 6.538171e-08, 6.543657e-08, 6.530066e-08, 6.545889e-08, 
    6.548544e-08, 6.541601e-08, 6.581894e-08, 6.570383e-08, 6.582162e-08, 
    6.574668e-08, 6.386237e-08, 6.395581e-08, 6.390532e-08, 6.400027e-08, 
    6.393338e-08, 6.42308e-08, 6.431998e-08, 6.473723e-08, 6.456598e-08, 
    6.483852e-08, 6.459366e-08, 6.463705e-08, 6.484741e-08, 6.460689e-08, 
    6.513292e-08, 6.47763e-08, 6.543871e-08, 6.50826e-08, 6.546102e-08, 
    6.53923e-08, 6.550608e-08, 6.560798e-08, 6.573618e-08, 6.597273e-08, 
    6.591795e-08, 6.611577e-08, 6.40951e-08, 6.42163e-08, 6.420562e-08, 
    6.433245e-08, 6.442625e-08, 6.462955e-08, 6.49556e-08, 6.483299e-08, 
    6.505808e-08, 6.510327e-08, 6.476129e-08, 6.497127e-08, 6.42974e-08, 
    6.440629e-08, 6.434146e-08, 6.410467e-08, 6.486125e-08, 6.447298e-08, 
    6.518994e-08, 6.49796e-08, 6.559345e-08, 6.528818e-08, 6.58878e-08, 
    6.614415e-08, 6.638538e-08, 6.666732e-08, 6.428244e-08, 6.420009e-08, 
    6.434753e-08, 6.455154e-08, 6.47408e-08, 6.499243e-08, 6.501818e-08, 
    6.506531e-08, 6.518741e-08, 6.529008e-08, 6.508023e-08, 6.531582e-08, 
    6.443155e-08, 6.489495e-08, 6.416896e-08, 6.438758e-08, 6.453951e-08, 
    6.447286e-08, 6.481897e-08, 6.490055e-08, 6.523204e-08, 6.506068e-08, 
    6.608088e-08, 6.562952e-08, 6.688197e-08, 6.653197e-08, 6.417132e-08, 
    6.428215e-08, 6.466789e-08, 6.448436e-08, 6.500922e-08, 6.513842e-08, 
    6.524344e-08, 6.53777e-08, 6.539219e-08, 6.547174e-08, 6.534139e-08, 
    6.546659e-08, 6.499297e-08, 6.520462e-08, 6.46238e-08, 6.476517e-08, 
    6.470013e-08, 6.46288e-08, 6.484896e-08, 6.508353e-08, 6.508854e-08, 
    6.516375e-08, 6.537572e-08, 6.501136e-08, 6.613915e-08, 6.544267e-08, 
    6.440301e-08, 6.461651e-08, 6.464699e-08, 6.456429e-08, 6.512547e-08, 
    6.492213e-08, 6.54698e-08, 6.532179e-08, 6.55643e-08, 6.544379e-08, 
    6.542606e-08, 6.527128e-08, 6.517492e-08, 6.493146e-08, 6.473337e-08, 
    6.457628e-08, 6.461281e-08, 6.478536e-08, 6.509788e-08, 6.539351e-08, 
    6.532875e-08, 6.554587e-08, 6.497117e-08, 6.521216e-08, 6.511902e-08, 
    6.536187e-08, 6.482973e-08, 6.52829e-08, 6.471389e-08, 6.476378e-08, 
    6.49181e-08, 6.522851e-08, 6.529717e-08, 6.53705e-08, 6.532525e-08, 
    6.510581e-08, 6.506986e-08, 6.491435e-08, 6.487141e-08, 6.475292e-08, 
    6.465483e-08, 6.474446e-08, 6.483858e-08, 6.51059e-08, 6.53468e-08, 
    6.560944e-08, 6.567371e-08, 6.59806e-08, 6.573079e-08, 6.614304e-08, 
    6.579257e-08, 6.639924e-08, 6.530915e-08, 6.578225e-08, 6.492512e-08, 
    6.501746e-08, 6.518448e-08, 6.556754e-08, 6.536073e-08, 6.560259e-08, 
    6.506844e-08, 6.479132e-08, 6.471961e-08, 6.458583e-08, 6.472267e-08, 
    6.471154e-08, 6.484247e-08, 6.48004e-08, 6.511478e-08, 6.494591e-08, 
    6.542562e-08, 6.560068e-08, 6.609504e-08, 6.63981e-08, 6.670659e-08, 
    6.684278e-08, 6.688423e-08, 6.690156e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999936, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999936, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999937, 
    0.9999936, 0.9999936, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999936, 
    0.9999937, 0.9999937, 0.9999936, 0.9999937, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999935, 0.9999935, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999937, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999935, 0.9999935, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999937, 0.9999937, 0.9999937, 0.9999937, 0.9999935, 0.9999934, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999936, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999936, 0.9999938, 0.9999937, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999935, 0.9999936, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999937, 0.9999936, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 0.9999937, 
    0.9999936, 0.9999937, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999937, 0.9999937, 0.9999937, 0.9999938, 
    0.9999938, 0.9999938 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.1477056, -0.1477207, -0.1477179, -0.1477299, -0.1477233, -0.1477311, 
    -0.1477088, -0.1477212, -0.1477134, -0.1477071, -0.1477515, -0.1477305, 
    -0.1477674, -0.1477586, -0.1477915, -0.1477659, -0.1477944, -0.1477913, 
    -0.1478011, -0.1477983, -0.1478105, -0.1478024, -0.1478171, -0.1478087, 
    -0.1478099, -0.1478021, -0.147735, -0.1477488, -0.1477341, -0.1477361, 
    -0.1477352, -0.1477234, -0.1477171, -0.1477046, -0.1477069, -0.1477162, 
    -0.147737, -0.1477304, -0.1477475, -0.1477471, -0.1477619, -0.1477562, 
    -0.1477879, -0.147771, -0.1477984, -0.1477944, -0.1477982, -0.1477971, 
    -0.1477982, -0.1477923, -0.1477948, -0.1477896, -0.1477574, -0.1477637, 
    -0.1477397, -0.1477213, -0.1477093, -0.1477006, -0.1477018, -0.1477041, 
    -0.1477162, -0.1477278, -0.1477362, -0.1477416, -0.147747, -0.1477598, 
    -0.1477655, -0.1477889, -0.1477869, -0.1477904, -0.147794, -0.1477997, 
    -0.1477988, -0.1478013, -0.1477904, -0.1477976, -0.1477743, -0.147789, 
    -0.1477476, -0.1477322, -0.1477245, -0.1477184, -0.1477027, -0.1477135, 
    -0.1477092, -0.1477196, -0.147726, -0.1477228, -0.1477418, -0.1477346, 
    -0.1477659, -0.1477551, -0.1477935, -0.1477873, -0.1477951, -0.1477911, 
    -0.1477978, -0.1477918, -0.1478023, -0.1478045, -0.147803, -0.1478091, 
    -0.1477915, -0.1477982, -0.1477227, -0.1477232, -0.1477257, -0.1477148, 
    -0.1477142, -0.1477045, -0.1477132, -0.1477169, -0.1477264, -0.1477318, 
    -0.1477368, -0.1477476, -0.1477578, -0.1477688, -0.1477877, -0.1477928, 
    -0.1477897, -0.1477924, -0.1477894, -0.147788, -0.1478036, -0.1477948, 
    -0.1478082, -0.1478075, -0.1478014, -0.1478075, -0.1477236, -0.1477206, 
    -0.1477101, -0.1477184, -0.1477035, -0.1477117, -0.1477164, -0.1477346, 
    -0.1477385, -0.147742, -0.147749, -0.1477565, -0.1477667, -0.1477865, 
    -0.1477942, -0.1477936, -0.1477938, -0.1477955, -0.1477913, -0.1477962, 
    -0.147797, -0.1477949, -0.1478074, -0.1478038, -0.1478074, -0.1478051, 
    -0.1477216, -0.1477266, -0.1477239, -0.1477289, -0.1477253, -0.1477405, 
    -0.147745, -0.147762, -0.1477564, -0.1477654, -0.1477575, -0.1477588, 
    -0.1477654, -0.1477579, -0.1477745, -0.1477632, -0.1477956, -0.1477728, 
    -0.1477963, -0.1477942, -0.1477977, -0.1478008, -0.1478048, -0.147812, 
    -0.1478104, -0.1478165, -0.1477339, -0.1477399, -0.1477395, -0.1477459, 
    -0.1477506, -0.1477587, -0.1477692, -0.1477653, -0.1477724, -0.1477737, 
    -0.147763, -0.1477696, -0.147744, -0.1477493, -0.1477463, -0.1477343, 
    -0.1477661, -0.1477527, -0.1477878, -0.14777, -0.1478003, -0.1477908, 
    -0.1478094, -0.1478171, -0.1478249, -0.1478334, -0.1477433, -0.1477393, 
    -0.1477467, -0.1477557, -0.1477623, -0.1477703, -0.1477712, -0.1477726, 
    -0.1477878, -0.147791, -0.1477729, -0.1477918, -0.1477502, -0.1477672, 
    -0.1477376, -0.1477484, -0.1477553, -0.1477529, -0.1477649, -0.1477676, 
    -0.1477891, -0.1477724, -0.1478151, -0.1478013, -0.1478402, -0.1478292, 
    -0.1477378, -0.1477434, -0.1477598, -0.1477534, -0.1477709, -0.1477748, 
    -0.1477896, -0.1477936, -0.1477941, -0.1477966, -0.1477926, -0.1477965, 
    -0.1477703, -0.1477883, -0.1477585, -0.1477631, -0.147761, -0.1477587, 
    -0.1477659, -0.147773, -0.1477733, -0.147787, -0.147793, -0.147771, 
    -0.1478166, -0.1477951, -0.1477495, -0.147758, -0.1477592, -0.1477564, 
    -0.1477744, -0.1477682, -0.1477965, -0.147792, -0.1477995, -0.1477957, 
    -0.1477952, -0.1477904, -0.1477874, -0.1477685, -0.147762, -0.1477569, 
    -0.1477581, -0.1477637, -0.1477734, -0.1477941, -0.1477921, -0.1477989, 
    -0.1477697, -0.1477885, -0.1477741, -0.1477932, -0.1477652, -0.1477902, 
    -0.1477615, -0.1477631, -0.1477681, -0.1477889, -0.1477912, -0.1477934, 
    -0.1477921, -0.1477737, -0.1477727, -0.147768, -0.1477665, -0.1477627, 
    -0.1477595, -0.1477624, -0.1477654, -0.1477738, -0.1477927, -0.1478008, 
    -0.1478029, -0.147812, -0.1478043, -0.1478167, -0.1478058, -0.1478248, 
    -0.1477912, -0.1478058, -0.1477684, -0.1477711, -0.1477875, -0.1477994, 
    -0.1477931, -0.1478005, -0.1477726, -0.1477638, -0.1477616, -0.1477572, 
    -0.1477617, -0.1477614, -0.1477657, -0.1477643, -0.1477741, -0.147769, 
    -0.1477951, -0.1478005, -0.1478158, -0.1478251, -0.1478348, -0.147839, 
    -0.1478403, -0.1478408 ;

 TAUY =
  -0.1477056, -0.1477207, -0.1477179, -0.1477299, -0.1477233, -0.1477311, 
    -0.1477088, -0.1477212, -0.1477134, -0.1477071, -0.1477515, -0.1477305, 
    -0.1477674, -0.1477586, -0.1477915, -0.1477659, -0.1477944, -0.1477913, 
    -0.1478011, -0.1477983, -0.1478105, -0.1478024, -0.1478171, -0.1478087, 
    -0.1478099, -0.1478021, -0.147735, -0.1477488, -0.1477341, -0.1477361, 
    -0.1477352, -0.1477234, -0.1477171, -0.1477046, -0.1477069, -0.1477162, 
    -0.147737, -0.1477304, -0.1477475, -0.1477471, -0.1477619, -0.1477562, 
    -0.1477879, -0.147771, -0.1477984, -0.1477944, -0.1477982, -0.1477971, 
    -0.1477982, -0.1477923, -0.1477948, -0.1477896, -0.1477574, -0.1477637, 
    -0.1477397, -0.1477213, -0.1477093, -0.1477006, -0.1477018, -0.1477041, 
    -0.1477162, -0.1477278, -0.1477362, -0.1477416, -0.147747, -0.1477598, 
    -0.1477655, -0.1477889, -0.1477869, -0.1477904, -0.147794, -0.1477997, 
    -0.1477988, -0.1478013, -0.1477904, -0.1477976, -0.1477743, -0.147789, 
    -0.1477476, -0.1477322, -0.1477245, -0.1477184, -0.1477027, -0.1477135, 
    -0.1477092, -0.1477196, -0.147726, -0.1477228, -0.1477418, -0.1477346, 
    -0.1477659, -0.1477551, -0.1477935, -0.1477873, -0.1477951, -0.1477911, 
    -0.1477978, -0.1477918, -0.1478023, -0.1478045, -0.147803, -0.1478091, 
    -0.1477915, -0.1477982, -0.1477227, -0.1477232, -0.1477257, -0.1477148, 
    -0.1477142, -0.1477045, -0.1477132, -0.1477169, -0.1477264, -0.1477318, 
    -0.1477368, -0.1477476, -0.1477578, -0.1477688, -0.1477877, -0.1477928, 
    -0.1477897, -0.1477924, -0.1477894, -0.147788, -0.1478036, -0.1477948, 
    -0.1478082, -0.1478075, -0.1478014, -0.1478075, -0.1477236, -0.1477206, 
    -0.1477101, -0.1477184, -0.1477035, -0.1477117, -0.1477164, -0.1477346, 
    -0.1477385, -0.147742, -0.147749, -0.1477565, -0.1477667, -0.1477865, 
    -0.1477942, -0.1477936, -0.1477938, -0.1477955, -0.1477913, -0.1477962, 
    -0.147797, -0.1477949, -0.1478074, -0.1478038, -0.1478074, -0.1478051, 
    -0.1477216, -0.1477266, -0.1477239, -0.1477289, -0.1477253, -0.1477405, 
    -0.147745, -0.147762, -0.1477564, -0.1477654, -0.1477575, -0.1477588, 
    -0.1477654, -0.1477579, -0.1477745, -0.1477632, -0.1477956, -0.1477728, 
    -0.1477963, -0.1477942, -0.1477977, -0.1478008, -0.1478048, -0.147812, 
    -0.1478104, -0.1478165, -0.1477339, -0.1477399, -0.1477395, -0.1477459, 
    -0.1477506, -0.1477587, -0.1477692, -0.1477653, -0.1477724, -0.1477737, 
    -0.147763, -0.1477696, -0.147744, -0.1477493, -0.1477463, -0.1477343, 
    -0.1477661, -0.1477527, -0.1477878, -0.14777, -0.1478003, -0.1477908, 
    -0.1478094, -0.1478171, -0.1478249, -0.1478334, -0.1477433, -0.1477393, 
    -0.1477467, -0.1477557, -0.1477623, -0.1477703, -0.1477712, -0.1477726, 
    -0.1477878, -0.147791, -0.1477729, -0.1477918, -0.1477502, -0.1477672, 
    -0.1477376, -0.1477484, -0.1477553, -0.1477529, -0.1477649, -0.1477676, 
    -0.1477891, -0.1477724, -0.1478151, -0.1478013, -0.1478402, -0.1478292, 
    -0.1477378, -0.1477434, -0.1477598, -0.1477534, -0.1477709, -0.1477748, 
    -0.1477896, -0.1477936, -0.1477941, -0.1477966, -0.1477926, -0.1477965, 
    -0.1477703, -0.1477883, -0.1477585, -0.1477631, -0.147761, -0.1477587, 
    -0.1477659, -0.147773, -0.1477733, -0.147787, -0.147793, -0.147771, 
    -0.1478166, -0.1477951, -0.1477495, -0.147758, -0.1477592, -0.1477564, 
    -0.1477744, -0.1477682, -0.1477965, -0.147792, -0.1477995, -0.1477957, 
    -0.1477952, -0.1477904, -0.1477874, -0.1477685, -0.147762, -0.1477569, 
    -0.1477581, -0.1477637, -0.1477734, -0.1477941, -0.1477921, -0.1477989, 
    -0.1477697, -0.1477885, -0.1477741, -0.1477932, -0.1477652, -0.1477902, 
    -0.1477615, -0.1477631, -0.1477681, -0.1477889, -0.1477912, -0.1477934, 
    -0.1477921, -0.1477737, -0.1477727, -0.147768, -0.1477665, -0.1477627, 
    -0.1477595, -0.1477624, -0.1477654, -0.1477738, -0.1477927, -0.1478008, 
    -0.1478029, -0.147812, -0.1478043, -0.1478167, -0.1478058, -0.1478248, 
    -0.1477912, -0.1478058, -0.1477684, -0.1477711, -0.1477875, -0.1477994, 
    -0.1477931, -0.1478005, -0.1477726, -0.1477638, -0.1477616, -0.1477572, 
    -0.1477617, -0.1477614, -0.1477657, -0.1477643, -0.1477741, -0.147769, 
    -0.1477951, -0.1478005, -0.1478158, -0.1478251, -0.1478348, -0.147839, 
    -0.1478403, -0.1478408 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.6828, 261.6993, 261.6961, 261.7094, 261.7021, 261.7108, 261.6862, 
    261.7, 261.6912, 261.6843, 261.7353, 261.7101, 261.7617, 261.7456, 
    261.7861, 261.7592, 261.7915, 261.7853, 261.8041, 261.7987, 261.8226, 
    261.8066, 261.8351, 261.8188, 261.8213, 261.806, 261.7152, 261.7321, 
    261.7142, 261.7166, 261.7155, 261.7022, 261.6955, 261.6815, 261.6841, 
    261.6943, 261.7177, 261.7098, 261.7297, 261.7293, 261.7515, 261.7415, 
    261.7788, 261.7683, 261.799, 261.7912, 261.7986, 261.7964, 261.7986, 
    261.7873, 261.7921, 261.7821, 261.7434, 261.7548, 261.7208, 261.7003, 
    261.6868, 261.6772, 261.6785, 261.6811, 261.6944, 261.707, 261.7165, 
    261.7229, 261.7292, 261.7482, 261.7584, 261.7809, 261.7769, 261.7838, 
    261.7904, 261.8015, 261.7997, 261.8046, 261.7836, 261.7975, 261.7747, 
    261.7809, 261.7308, 261.7119, 261.7038, 261.6967, 261.6795, 261.6914, 
    261.6867, 261.6979, 261.705, 261.7015, 261.7231, 261.7147, 261.759, 
    261.7399, 261.7897, 261.7777, 261.7925, 261.785, 261.7979, 261.7863, 
    261.8064, 261.8108, 261.8078, 261.8193, 261.7856, 261.7986, 261.7014, 
    261.7019, 261.7046, 261.6929, 261.6922, 261.6815, 261.691, 261.6951, 
    261.7054, 261.7115, 261.7173, 261.73, 261.7443, 261.7643, 261.7785, 
    261.7881, 261.7822, 261.7874, 261.7816, 261.7789, 261.8091, 261.7921, 
    261.8177, 261.8163, 261.8047, 261.8164, 261.7024, 261.6991, 261.6877, 
    261.6966, 261.6803, 261.6894, 261.6946, 261.7148, 261.7193, 261.7234, 
    261.7316, 261.742, 261.7603, 261.7762, 261.7908, 261.7898, 261.7901, 
    261.7934, 261.7853, 261.7947, 261.7963, 261.7922, 261.8161, 261.8093, 
    261.8163, 261.8118, 261.7001, 261.7057, 261.7027, 261.7083, 261.7043, 
    261.7219, 261.7272, 261.7519, 261.7418, 261.758, 261.7434, 261.746, 
    261.7584, 261.7442, 261.7754, 261.7542, 261.7935, 261.7724, 261.7948, 
    261.7908, 261.7975, 261.8036, 261.8112, 261.8252, 261.822, 261.8337, 
    261.7139, 261.7211, 261.7205, 261.728, 261.7335, 261.7456, 261.765, 
    261.7577, 261.7711, 261.7737, 261.7534, 261.7659, 261.7259, 261.7323, 
    261.7285, 261.7144, 261.7593, 261.7362, 261.7787, 261.7664, 261.8027, 
    261.7845, 261.8202, 261.8353, 261.8497, 261.8663, 261.725, 261.7201, 
    261.7289, 261.7409, 261.7522, 261.7671, 261.7687, 261.7715, 261.7786, 
    261.7847, 261.7723, 261.7862, 261.7337, 261.7613, 261.7183, 261.7312, 
    261.7402, 261.7363, 261.7568, 261.7617, 261.7812, 261.7712, 261.8315, 
    261.8048, 261.8791, 261.8583, 261.7184, 261.725, 261.7478, 261.737, 
    261.7682, 261.7758, 261.7819, 261.7899, 261.7908, 261.7955, 261.7878, 
    261.7952, 261.7672, 261.7796, 261.7453, 261.7536, 261.7498, 261.7455, 
    261.7586, 261.7725, 261.7729, 261.7772, 261.7896, 261.7683, 261.8349, 
    261.7936, 261.7321, 261.7448, 261.7466, 261.7417, 261.775, 261.763, 
    261.7953, 261.7866, 261.801, 261.7938, 261.7928, 261.7836, 261.7779, 
    261.7635, 261.7517, 261.7424, 261.7446, 261.7548, 261.7734, 261.7908, 
    261.787, 261.7999, 261.7659, 261.78, 261.7746, 261.7889, 261.7575, 
    261.7841, 261.7506, 261.7536, 261.7627, 261.781, 261.7851, 261.7895, 
    261.7868, 261.7739, 261.7717, 261.7625, 261.7599, 261.7529, 261.7471, 
    261.7524, 261.758, 261.7739, 261.7881, 261.8036, 261.8075, 261.8256, 
    261.8108, 261.8351, 261.8143, 261.8504, 261.7857, 261.8138, 261.7632, 
    261.7686, 261.7784, 261.8011, 261.7889, 261.8032, 261.7716, 261.7552, 
    261.7509, 261.743, 261.7511, 261.7505, 261.7582, 261.7557, 261.7744, 
    261.7644, 261.7927, 261.8031, 261.8324, 261.8504, 261.8687, 261.8768, 
    261.8793, 261.8803 ;

 TG_R =
  261.6828, 261.6993, 261.6961, 261.7094, 261.7021, 261.7108, 261.6862, 
    261.7, 261.6912, 261.6843, 261.7353, 261.7101, 261.7617, 261.7456, 
    261.7861, 261.7592, 261.7915, 261.7853, 261.8041, 261.7987, 261.8226, 
    261.8066, 261.8351, 261.8188, 261.8213, 261.806, 261.7152, 261.7321, 
    261.7142, 261.7166, 261.7155, 261.7022, 261.6955, 261.6815, 261.6841, 
    261.6943, 261.7177, 261.7098, 261.7297, 261.7293, 261.7515, 261.7415, 
    261.7788, 261.7683, 261.799, 261.7912, 261.7986, 261.7964, 261.7986, 
    261.7873, 261.7921, 261.7821, 261.7434, 261.7548, 261.7208, 261.7003, 
    261.6868, 261.6772, 261.6785, 261.6811, 261.6944, 261.707, 261.7165, 
    261.7229, 261.7292, 261.7482, 261.7584, 261.7809, 261.7769, 261.7838, 
    261.7904, 261.8015, 261.7997, 261.8046, 261.7836, 261.7975, 261.7747, 
    261.7809, 261.7308, 261.7119, 261.7038, 261.6967, 261.6795, 261.6914, 
    261.6867, 261.6979, 261.705, 261.7015, 261.7231, 261.7147, 261.759, 
    261.7399, 261.7897, 261.7777, 261.7925, 261.785, 261.7979, 261.7863, 
    261.8064, 261.8108, 261.8078, 261.8193, 261.7856, 261.7986, 261.7014, 
    261.7019, 261.7046, 261.6929, 261.6922, 261.6815, 261.691, 261.6951, 
    261.7054, 261.7115, 261.7173, 261.73, 261.7443, 261.7643, 261.7785, 
    261.7881, 261.7822, 261.7874, 261.7816, 261.7789, 261.8091, 261.7921, 
    261.8177, 261.8163, 261.8047, 261.8164, 261.7024, 261.6991, 261.6877, 
    261.6966, 261.6803, 261.6894, 261.6946, 261.7148, 261.7193, 261.7234, 
    261.7316, 261.742, 261.7603, 261.7762, 261.7908, 261.7898, 261.7901, 
    261.7934, 261.7853, 261.7947, 261.7963, 261.7922, 261.8161, 261.8093, 
    261.8163, 261.8118, 261.7001, 261.7057, 261.7027, 261.7083, 261.7043, 
    261.7219, 261.7272, 261.7519, 261.7418, 261.758, 261.7434, 261.746, 
    261.7584, 261.7442, 261.7754, 261.7542, 261.7935, 261.7724, 261.7948, 
    261.7908, 261.7975, 261.8036, 261.8112, 261.8252, 261.822, 261.8337, 
    261.7139, 261.7211, 261.7205, 261.728, 261.7335, 261.7456, 261.765, 
    261.7577, 261.7711, 261.7737, 261.7534, 261.7659, 261.7259, 261.7323, 
    261.7285, 261.7144, 261.7593, 261.7362, 261.7787, 261.7664, 261.8027, 
    261.7845, 261.8202, 261.8353, 261.8497, 261.8663, 261.725, 261.7201, 
    261.7289, 261.7409, 261.7522, 261.7671, 261.7687, 261.7715, 261.7786, 
    261.7847, 261.7723, 261.7862, 261.7337, 261.7613, 261.7183, 261.7312, 
    261.7402, 261.7363, 261.7568, 261.7617, 261.7812, 261.7712, 261.8315, 
    261.8048, 261.8791, 261.8583, 261.7184, 261.725, 261.7478, 261.737, 
    261.7682, 261.7758, 261.7819, 261.7899, 261.7908, 261.7955, 261.7878, 
    261.7952, 261.7672, 261.7796, 261.7453, 261.7536, 261.7498, 261.7455, 
    261.7586, 261.7725, 261.7729, 261.7772, 261.7896, 261.7683, 261.8349, 
    261.7936, 261.7321, 261.7448, 261.7466, 261.7417, 261.775, 261.763, 
    261.7953, 261.7866, 261.801, 261.7938, 261.7928, 261.7836, 261.7779, 
    261.7635, 261.7517, 261.7424, 261.7446, 261.7548, 261.7734, 261.7908, 
    261.787, 261.7999, 261.7659, 261.78, 261.7746, 261.7889, 261.7575, 
    261.7841, 261.7506, 261.7536, 261.7627, 261.781, 261.7851, 261.7895, 
    261.7868, 261.7739, 261.7717, 261.7625, 261.7599, 261.7529, 261.7471, 
    261.7524, 261.758, 261.7739, 261.7881, 261.8036, 261.8075, 261.8256, 
    261.8108, 261.8351, 261.8143, 261.8504, 261.7857, 261.8138, 261.7632, 
    261.7686, 261.7784, 261.8011, 261.7889, 261.8032, 261.7716, 261.7552, 
    261.7509, 261.743, 261.7511, 261.7505, 261.7582, 261.7557, 261.7744, 
    261.7644, 261.7927, 261.8031, 261.8324, 261.8504, 261.8687, 261.8768, 
    261.8793, 261.8803 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.015, 254.0168, 254.0165, 254.0179, 254.0172, 254.0181, 254.0154, 
    254.0169, 254.0159, 254.0152, 254.0208, 254.018, 254.0237, 254.022, 
    254.0264, 254.0234, 254.0271, 254.0264, 254.0285, 254.0279, 254.0305, 
    254.0287, 254.0319, 254.0301, 254.0303, 254.0287, 254.0186, 254.0204, 
    254.0185, 254.0187, 254.0186, 254.0172, 254.0164, 254.0149, 254.0152, 
    254.0163, 254.0189, 254.018, 254.0202, 254.0202, 254.0226, 254.0215, 
    254.0257, 254.0245, 254.0279, 254.027, 254.0278, 254.0276, 254.0279, 
    254.0266, 254.0271, 254.026, 254.0217, 254.023, 254.0192, 254.0169, 
    254.0154, 254.0144, 254.0145, 254.0148, 254.0163, 254.0177, 254.0188, 
    254.0195, 254.0202, 254.0222, 254.0234, 254.0259, 254.0255, 254.0262, 
    254.0269, 254.0282, 254.028, 254.0285, 254.0262, 254.0277, 254.0252, 
    254.0259, 254.0202, 254.0182, 254.0173, 254.0165, 254.0146, 254.0159, 
    254.0154, 254.0167, 254.0175, 254.0171, 254.0195, 254.0186, 254.0234, 
    254.0213, 254.0269, 254.0255, 254.0272, 254.0264, 254.0278, 254.0265, 
    254.0287, 254.0292, 254.0289, 254.0302, 254.0264, 254.0278, 254.0171, 
    254.0171, 254.0174, 254.0161, 254.016, 254.0148, 254.0159, 254.0164, 
    254.0175, 254.0182, 254.0188, 254.0202, 254.0218, 254.024, 254.0256, 
    254.0267, 254.026, 254.0266, 254.026, 254.0257, 254.029, 254.0271, 
    254.03, 254.0298, 254.0285, 254.0298, 254.0172, 254.0168, 254.0155, 
    254.0165, 254.0147, 254.0157, 254.0163, 254.0185, 254.0191, 254.0195, 
    254.0204, 254.0216, 254.0236, 254.0254, 254.027, 254.0269, 254.0269, 
    254.0273, 254.0264, 254.0274, 254.0276, 254.0271, 254.0298, 254.029, 
    254.0298, 254.0293, 254.0169, 254.0175, 254.0172, 254.0178, 254.0174, 
    254.0193, 254.0199, 254.0226, 254.0215, 254.0233, 254.0217, 254.022, 
    254.0233, 254.0218, 254.0253, 254.0229, 254.0273, 254.0249, 254.0274, 
    254.027, 254.0277, 254.0284, 254.0293, 254.0308, 254.0304, 254.0317, 
    254.0185, 254.0192, 254.0192, 254.02, 254.0206, 254.022, 254.0241, 
    254.0233, 254.0248, 254.0251, 254.0229, 254.0242, 254.0198, 254.0205, 
    254.0201, 254.0185, 254.0235, 254.0209, 254.0257, 254.0243, 254.0283, 
    254.0263, 254.0302, 254.0319, 254.0335, 254.0353, 254.0197, 254.0192, 
    254.0201, 254.0214, 254.0227, 254.0244, 254.0245, 254.0248, 254.0257, 
    254.0263, 254.0249, 254.0265, 254.0206, 254.0237, 254.0189, 254.0203, 
    254.0214, 254.0209, 254.0232, 254.0238, 254.0259, 254.0248, 254.0314, 
    254.0285, 254.0368, 254.0345, 254.019, 254.0197, 254.0222, 254.021, 
    254.0245, 254.0253, 254.026, 254.0269, 254.027, 254.0275, 254.0267, 
    254.0275, 254.0244, 254.0258, 254.022, 254.0229, 254.0224, 254.022, 
    254.0234, 254.0249, 254.025, 254.0255, 254.0267, 254.0245, 254.0318, 
    254.0272, 254.0205, 254.0219, 254.0221, 254.0216, 254.0252, 254.0239, 
    254.0275, 254.0265, 254.0281, 254.0273, 254.0272, 254.0262, 254.0256, 
    254.024, 254.0227, 254.0216, 254.0219, 254.023, 254.025, 254.027, 
    254.0266, 254.028, 254.0242, 254.0258, 254.0252, 254.0268, 254.0233, 
    254.0262, 254.0225, 254.0229, 254.0239, 254.0259, 254.0264, 254.0268, 
    254.0266, 254.0251, 254.0249, 254.0238, 254.0236, 254.0228, 254.0222, 
    254.0227, 254.0233, 254.0251, 254.0267, 254.0284, 254.0288, 254.0308, 
    254.0292, 254.0318, 254.0295, 254.0335, 254.0264, 254.0295, 254.0239, 
    254.0245, 254.0256, 254.0281, 254.0268, 254.0283, 254.0249, 254.023, 
    254.0226, 254.0217, 254.0226, 254.0225, 254.0234, 254.0231, 254.0252, 
    254.0241, 254.0272, 254.0283, 254.0316, 254.0336, 254.0356, 254.0365, 
    254.0368, 254.0369 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23988, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTCOLCH4 =
  1.357788e-05, 1.337091e-05, 1.341105e-05, 1.324484e-05, 1.333693e-05, 
    1.322826e-05, 1.353582e-05, 1.336272e-05, 1.347312e-05, 1.35592e-05, 
    1.292496e-05, 1.323745e-05, 1.268778e-05, 1.289718e-05, 1.237662e-05, 
    1.272018e-05, 1.230838e-05, 1.238642e-05, 1.215298e-05, 1.221941e-05, 
    1.192567e-05, 1.212244e-05, 1.177643e-05, 1.197235e-05, 1.194146e-05, 
    1.212899e-05, 1.317428e-05, 1.296367e-05, 1.318681e-05, 1.315666e-05, 
    1.317019e-05, 1.333503e-05, 1.341842e-05, 1.359375e-05, 1.356185e-05, 
    1.343311e-05, 1.314312e-05, 1.324125e-05, 1.299458e-05, 1.300013e-05, 
    1.281969e-05, 1.295036e-05, 1.246873e-05, 1.260406e-05, 1.221663e-05, 
    1.2313e-05, 1.222114e-05, 1.224893e-05, 1.222078e-05, 1.236241e-05, 
    1.230154e-05, 1.242687e-05, 1.292581e-05, 1.277748e-05, 1.310511e-05, 
    1.335867e-05, 1.352821e-05, 1.364901e-05, 1.363191e-05, 1.359933e-05, 
    1.343236e-05, 1.327613e-05, 1.315759e-05, 1.307857e-05, 1.300093e-05, 
    1.286152e-05, 1.27306e-05, 1.244152e-05, 1.249326e-05, 1.240572e-05, 
    1.232263e-05, 1.218432e-05, 1.220698e-05, 1.214642e-05, 1.240803e-05, 
    1.223356e-05, 1.252282e-05, 1.244308e-05, 1.297986e-05, 1.321475e-05, 
    1.331516e-05, 1.340333e-05, 1.361876e-05, 1.346985e-05, 1.352848e-05, 
    1.338915e-05, 1.330093e-05, 1.334453e-05, 1.307641e-05, 1.318036e-05, 
    1.272288e-05, 1.297112e-05, 1.233229e-05, 1.248263e-05, 1.229651e-05, 
    1.239116e-05, 1.222942e-05, 1.237489e-05, 1.212396e-05, 1.206999e-05, 
    1.210684e-05, 1.196594e-05, 1.238301e-05, 1.222114e-05, 1.334575e-05, 
    1.333864e-05, 1.330551e-05, 1.34514e-05, 1.346034e-05, 1.359462e-05, 
    1.347512e-05, 1.342435e-05, 1.329582e-05, 1.322004e-05, 1.314818e-05, 
    1.299083e-05, 1.291377e-05, 1.265561e-05, 1.247283e-05, 1.235164e-05, 
    1.242582e-05, 1.236031e-05, 1.243357e-05, 1.246804e-05, 1.209018e-05, 
    1.230097e-05, 1.19861e-05, 1.20033e-05, 1.214498e-05, 1.200136e-05, 
    1.333364e-05, 1.337461e-05, 1.351723e-05, 1.340556e-05, 1.360928e-05, 
    1.34951e-05, 1.342962e-05, 1.317818e-05, 1.312322e-05, 1.307235e-05, 
    1.297216e-05, 1.294364e-05, 1.270567e-05, 1.250157e-05, 1.231781e-05, 
    1.233119e-05, 1.232648e-05, 1.228575e-05, 1.238687e-05, 1.226922e-05, 
    1.224958e-05, 1.2301e-05, 1.200561e-05, 1.208925e-05, 1.200367e-05, 
    1.205805e-05, 1.336129e-05, 1.329241e-05, 1.332961e-05, 1.32597e-05, 
    1.330894e-05, 1.309063e-05, 1.30255e-05, 1.28141e-05, 1.294633e-05, 
    1.273639e-05, 1.292489e-05, 1.289133e-05, 1.272958e-05, 1.291464e-05, 
    1.251275e-05, 1.278408e-05, 1.228417e-05, 1.255073e-05, 1.226764e-05, 
    1.23186e-05, 1.223434e-05, 1.215935e-05, 1.206568e-05, 1.189484e-05, 
    1.193416e-05, 1.179282e-05, 1.319003e-05, 1.310123e-05, 1.310904e-05, 
    1.301639e-05, 1.294808e-05, 1.289713e-05, 1.264704e-05, 1.274062e-05, 
    1.256927e-05, 1.253512e-05, 1.27956e-05, 1.263513e-05, 1.304196e-05, 
    1.296261e-05, 1.300983e-05, 1.318301e-05, 1.2719e-05, 1.291413e-05, 
    1.246983e-05, 1.262879e-05, 1.217002e-05, 1.23962e-05, 1.195587e-05, 
    1.177271e-05, 1.160331e-05, 1.140915e-05, 1.305289e-05, 1.311309e-05, 
    1.30054e-05, 1.295754e-05, 1.281135e-05, 1.261904e-05, 1.259951e-05, 
    1.25638e-05, 1.247172e-05, 1.239478e-05, 1.255253e-05, 1.237556e-05, 
    1.294424e-05, 1.269326e-05, 1.313588e-05, 1.297623e-05, 1.296687e-05, 
    1.291421e-05, 1.275135e-05, 1.268898e-05, 1.243823e-05, 1.256731e-05, 
    1.181761e-05, 1.214357e-05, 1.12642e-05, 1.150183e-05, 1.313415e-05, 
    1.30531e-05, 1.286751e-05, 1.290585e-05, 1.260629e-05, 1.25086e-05, 
    1.242968e-05, 1.232946e-05, 1.231868e-05, 1.225972e-05, 1.235649e-05, 
    1.226352e-05, 1.261864e-05, 1.24588e-05, 1.290157e-05, 1.279262e-05, 
    1.284265e-05, 1.28977e-05, 1.272839e-05, 1.255003e-05, 1.254624e-05, 
    1.248953e-05, 1.233094e-05, 1.260468e-05, 1.177624e-05, 1.228124e-05, 
    1.296499e-05, 1.290721e-05, 1.288365e-05, 1.294764e-05, 1.251836e-05, 
    1.267252e-05, 1.226115e-05, 1.237111e-05, 1.219144e-05, 1.22804e-05, 
    1.229354e-05, 1.240884e-05, 1.248112e-05, 1.266542e-05, 1.281706e-05, 
    1.293835e-05, 1.291007e-05, 1.277712e-05, 1.253919e-05, 1.231771e-05, 
    1.236591e-05, 1.220501e-05, 1.26352e-05, 1.245314e-05, 1.252323e-05, 
    1.234123e-05, 1.274311e-05, 1.240015e-05, 1.283205e-05, 1.279368e-05, 
    1.26756e-05, 1.244088e-05, 1.238948e-05, 1.233481e-05, 1.236852e-05, 
    1.25332e-05, 1.256037e-05, 1.267846e-05, 1.271123e-05, 1.280203e-05, 
    1.28776e-05, 1.280854e-05, 1.273634e-05, 1.253313e-05, 1.235246e-05, 
    1.215829e-05, 1.211124e-05, 1.18892e-05, 1.206961e-05, 1.17735e-05, 
    1.202473e-05, 1.159367e-05, 1.238054e-05, 1.203221e-05, 1.267025e-05, 
    1.260005e-05, 1.247393e-05, 1.218906e-05, 1.234208e-05, 1.216331e-05, 
    1.256143e-05, 1.277255e-05, 1.282765e-05, 1.293095e-05, 1.28253e-05, 
    1.283386e-05, 1.273335e-05, 1.276558e-05, 1.252643e-05, 1.265442e-05, 
    1.229387e-05, 1.216472e-05, 1.180754e-05, 1.159446e-05, 1.138245e-05, 
    1.129048e-05, 1.126269e-05, 1.12511e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23988, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976208e-05, 5.976193e-05, 5.976196e-05, 5.976184e-05, 5.976191e-05, 
    5.976183e-05, 5.976205e-05, 5.976193e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976184e-05, 5.976138e-05, 5.976153e-05, 5.976117e-05, 
    5.976141e-05, 5.976112e-05, 5.976118e-05, 5.976101e-05, 5.976106e-05, 
    5.976085e-05, 5.976099e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976179e-05, 5.976164e-05, 5.97618e-05, 5.976178e-05, 
    5.976179e-05, 5.976191e-05, 5.976197e-05, 5.976209e-05, 5.976207e-05, 
    5.976198e-05, 5.976177e-05, 5.976184e-05, 5.976166e-05, 5.976167e-05, 
    5.976147e-05, 5.976156e-05, 5.976123e-05, 5.976133e-05, 5.976106e-05, 
    5.976113e-05, 5.976106e-05, 5.976108e-05, 5.976106e-05, 5.976116e-05, 
    5.976112e-05, 5.976121e-05, 5.976154e-05, 5.976145e-05, 5.976174e-05, 
    5.976192e-05, 5.976204e-05, 5.976213e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976178e-05, 5.976172e-05, 5.976167e-05, 
    5.97615e-05, 5.976141e-05, 5.976121e-05, 5.976125e-05, 5.976119e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.976101e-05, 5.976119e-05, 
    5.976107e-05, 5.976127e-05, 5.976122e-05, 5.976165e-05, 5.976182e-05, 
    5.976189e-05, 5.976195e-05, 5.976211e-05, 5.9762e-05, 5.976204e-05, 
    5.976194e-05, 5.976188e-05, 5.976191e-05, 5.976172e-05, 5.976179e-05, 
    5.976141e-05, 5.976157e-05, 5.976114e-05, 5.976124e-05, 5.976111e-05, 
    5.976118e-05, 5.976107e-05, 5.976117e-05, 5.976099e-05, 5.976095e-05, 
    5.976098e-05, 5.976088e-05, 5.976117e-05, 5.976106e-05, 5.976191e-05, 
    5.976191e-05, 5.976189e-05, 5.976199e-05, 5.976199e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976188e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976154e-05, 5.976136e-05, 5.976123e-05, 5.976115e-05, 
    5.97612e-05, 5.976116e-05, 5.976121e-05, 5.976123e-05, 5.976097e-05, 
    5.976111e-05, 5.976089e-05, 5.976091e-05, 5.976101e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.97621e-05, 
    5.976202e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976172e-05, 
    5.976165e-05, 5.976155e-05, 5.976139e-05, 5.976126e-05, 5.976113e-05, 
    5.976114e-05, 5.976113e-05, 5.97611e-05, 5.976118e-05, 5.976109e-05, 
    5.976108e-05, 5.976111e-05, 5.976091e-05, 5.976097e-05, 5.976091e-05, 
    5.976094e-05, 5.976193e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976189e-05, 5.976173e-05, 5.976169e-05, 5.976147e-05, 5.976156e-05, 
    5.976142e-05, 5.976154e-05, 5.976152e-05, 5.976141e-05, 5.976154e-05, 
    5.976126e-05, 5.976145e-05, 5.97611e-05, 5.976129e-05, 5.976109e-05, 
    5.976113e-05, 5.976107e-05, 5.976102e-05, 5.976095e-05, 5.976083e-05, 
    5.976086e-05, 5.976075e-05, 5.97618e-05, 5.976174e-05, 5.976174e-05, 
    5.976168e-05, 5.976163e-05, 5.976153e-05, 5.976135e-05, 5.976142e-05, 
    5.97613e-05, 5.976128e-05, 5.976146e-05, 5.976135e-05, 5.97617e-05, 
    5.976164e-05, 5.976167e-05, 5.97618e-05, 5.976141e-05, 5.976161e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976074e-05, 5.976061e-05, 5.976047e-05, 5.97617e-05, 5.976175e-05, 
    5.976167e-05, 5.976157e-05, 5.976147e-05, 5.976134e-05, 5.976132e-05, 
    5.97613e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976117e-05, 
    5.976163e-05, 5.976139e-05, 5.976177e-05, 5.976165e-05, 5.976157e-05, 
    5.976161e-05, 5.976143e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976077e-05, 5.976101e-05, 5.976036e-05, 5.976054e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.97616e-05, 5.976133e-05, 5.976126e-05, 
    5.976121e-05, 5.976114e-05, 5.976113e-05, 5.976109e-05, 5.976115e-05, 
    5.976109e-05, 5.976134e-05, 5.976123e-05, 5.976153e-05, 5.976145e-05, 
    5.976149e-05, 5.976153e-05, 5.976141e-05, 5.976129e-05, 5.976129e-05, 
    5.976125e-05, 5.976114e-05, 5.976133e-05, 5.976074e-05, 5.97611e-05, 
    5.976164e-05, 5.976153e-05, 5.976151e-05, 5.976156e-05, 5.976127e-05, 
    5.976137e-05, 5.976109e-05, 5.976117e-05, 5.976104e-05, 5.97611e-05, 
    5.976111e-05, 5.976119e-05, 5.976124e-05, 5.976137e-05, 5.976147e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976128e-05, 5.976113e-05, 
    5.976116e-05, 5.976105e-05, 5.976135e-05, 5.976122e-05, 5.976127e-05, 
    5.976114e-05, 5.976142e-05, 5.976118e-05, 5.976148e-05, 5.976146e-05, 
    5.976137e-05, 5.976121e-05, 5.976118e-05, 5.976114e-05, 5.976116e-05, 
    5.976128e-05, 5.97613e-05, 5.976138e-05, 5.97614e-05, 5.976146e-05, 
    5.976151e-05, 5.976146e-05, 5.976142e-05, 5.976128e-05, 5.976115e-05, 
    5.976102e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976074e-05, 
    5.976092e-05, 5.976061e-05, 5.976117e-05, 5.976093e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976104e-05, 5.976114e-05, 5.976102e-05, 
    5.97613e-05, 5.976144e-05, 5.976148e-05, 5.976155e-05, 5.976147e-05, 
    5.976148e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976136e-05, 
    5.976111e-05, 5.976102e-05, 5.976076e-05, 5.976061e-05, 5.976045e-05, 
    5.976038e-05, 5.976036e-05, 5.976035e-05 ;

 TOTLITC_1m =
  5.976208e-05, 5.976193e-05, 5.976196e-05, 5.976184e-05, 5.976191e-05, 
    5.976183e-05, 5.976205e-05, 5.976193e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976184e-05, 5.976138e-05, 5.976153e-05, 5.976117e-05, 
    5.976141e-05, 5.976112e-05, 5.976118e-05, 5.976101e-05, 5.976106e-05, 
    5.976085e-05, 5.976099e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976179e-05, 5.976164e-05, 5.97618e-05, 5.976178e-05, 
    5.976179e-05, 5.976191e-05, 5.976197e-05, 5.976209e-05, 5.976207e-05, 
    5.976198e-05, 5.976177e-05, 5.976184e-05, 5.976166e-05, 5.976167e-05, 
    5.976147e-05, 5.976156e-05, 5.976123e-05, 5.976133e-05, 5.976106e-05, 
    5.976113e-05, 5.976106e-05, 5.976108e-05, 5.976106e-05, 5.976116e-05, 
    5.976112e-05, 5.976121e-05, 5.976154e-05, 5.976145e-05, 5.976174e-05, 
    5.976192e-05, 5.976204e-05, 5.976213e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976178e-05, 5.976172e-05, 5.976167e-05, 
    5.97615e-05, 5.976141e-05, 5.976121e-05, 5.976125e-05, 5.976119e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.976101e-05, 5.976119e-05, 
    5.976107e-05, 5.976127e-05, 5.976122e-05, 5.976165e-05, 5.976182e-05, 
    5.976189e-05, 5.976195e-05, 5.976211e-05, 5.9762e-05, 5.976204e-05, 
    5.976194e-05, 5.976188e-05, 5.976191e-05, 5.976172e-05, 5.976179e-05, 
    5.976141e-05, 5.976157e-05, 5.976114e-05, 5.976124e-05, 5.976111e-05, 
    5.976118e-05, 5.976107e-05, 5.976117e-05, 5.976099e-05, 5.976095e-05, 
    5.976098e-05, 5.976088e-05, 5.976117e-05, 5.976106e-05, 5.976191e-05, 
    5.976191e-05, 5.976189e-05, 5.976199e-05, 5.976199e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976188e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976154e-05, 5.976136e-05, 5.976123e-05, 5.976115e-05, 
    5.97612e-05, 5.976116e-05, 5.976121e-05, 5.976123e-05, 5.976097e-05, 
    5.976111e-05, 5.976089e-05, 5.976091e-05, 5.976101e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.97621e-05, 
    5.976202e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976172e-05, 
    5.976165e-05, 5.976155e-05, 5.976139e-05, 5.976126e-05, 5.976113e-05, 
    5.976114e-05, 5.976113e-05, 5.97611e-05, 5.976118e-05, 5.976109e-05, 
    5.976108e-05, 5.976111e-05, 5.976091e-05, 5.976097e-05, 5.976091e-05, 
    5.976094e-05, 5.976193e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976189e-05, 5.976173e-05, 5.976169e-05, 5.976147e-05, 5.976156e-05, 
    5.976142e-05, 5.976154e-05, 5.976152e-05, 5.976141e-05, 5.976154e-05, 
    5.976126e-05, 5.976145e-05, 5.97611e-05, 5.976129e-05, 5.976109e-05, 
    5.976113e-05, 5.976107e-05, 5.976102e-05, 5.976095e-05, 5.976083e-05, 
    5.976086e-05, 5.976075e-05, 5.97618e-05, 5.976174e-05, 5.976174e-05, 
    5.976168e-05, 5.976163e-05, 5.976153e-05, 5.976135e-05, 5.976142e-05, 
    5.97613e-05, 5.976128e-05, 5.976146e-05, 5.976135e-05, 5.97617e-05, 
    5.976164e-05, 5.976167e-05, 5.97618e-05, 5.976141e-05, 5.976161e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976074e-05, 5.976061e-05, 5.976047e-05, 5.97617e-05, 5.976175e-05, 
    5.976167e-05, 5.976157e-05, 5.976147e-05, 5.976134e-05, 5.976132e-05, 
    5.97613e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976117e-05, 
    5.976163e-05, 5.976139e-05, 5.976177e-05, 5.976165e-05, 5.976157e-05, 
    5.976161e-05, 5.976143e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976077e-05, 5.976101e-05, 5.976036e-05, 5.976054e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.97616e-05, 5.976133e-05, 5.976126e-05, 
    5.976121e-05, 5.976114e-05, 5.976113e-05, 5.976109e-05, 5.976115e-05, 
    5.976109e-05, 5.976134e-05, 5.976123e-05, 5.976153e-05, 5.976145e-05, 
    5.976149e-05, 5.976153e-05, 5.976141e-05, 5.976129e-05, 5.976129e-05, 
    5.976125e-05, 5.976114e-05, 5.976133e-05, 5.976074e-05, 5.97611e-05, 
    5.976164e-05, 5.976153e-05, 5.976151e-05, 5.976156e-05, 5.976127e-05, 
    5.976137e-05, 5.976109e-05, 5.976117e-05, 5.976104e-05, 5.97611e-05, 
    5.976111e-05, 5.976119e-05, 5.976124e-05, 5.976137e-05, 5.976147e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976128e-05, 5.976113e-05, 
    5.976116e-05, 5.976105e-05, 5.976135e-05, 5.976122e-05, 5.976127e-05, 
    5.976114e-05, 5.976142e-05, 5.976118e-05, 5.976148e-05, 5.976146e-05, 
    5.976137e-05, 5.976121e-05, 5.976118e-05, 5.976114e-05, 5.976116e-05, 
    5.976128e-05, 5.97613e-05, 5.976138e-05, 5.97614e-05, 5.976146e-05, 
    5.976151e-05, 5.976146e-05, 5.976142e-05, 5.976128e-05, 5.976115e-05, 
    5.976102e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976074e-05, 
    5.976092e-05, 5.976061e-05, 5.976117e-05, 5.976093e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976104e-05, 5.976114e-05, 5.976102e-05, 
    5.97613e-05, 5.976144e-05, 5.976148e-05, 5.976155e-05, 5.976147e-05, 
    5.976148e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976136e-05, 
    5.976111e-05, 5.976102e-05, 5.976076e-05, 5.976061e-05, 5.976045e-05, 
    5.976038e-05, 5.976036e-05, 5.976035e-05 ;

 TOTLITN =
  1.37593e-06, 1.375926e-06, 1.375927e-06, 1.375924e-06, 1.375926e-06, 
    1.375923e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 1.37593e-06, 
    1.375917e-06, 1.375924e-06, 1.375911e-06, 1.375915e-06, 1.375905e-06, 
    1.375911e-06, 1.375903e-06, 1.375905e-06, 1.3759e-06, 1.375902e-06, 
    1.375896e-06, 1.3759e-06, 1.375893e-06, 1.375897e-06, 1.375896e-06, 
    1.3759e-06, 1.375922e-06, 1.375918e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375931e-06, 1.37593e-06, 
    1.375927e-06, 1.375922e-06, 1.375924e-06, 1.375919e-06, 1.375919e-06, 
    1.375913e-06, 1.375916e-06, 1.375907e-06, 1.375909e-06, 1.375902e-06, 
    1.375903e-06, 1.375902e-06, 1.375902e-06, 1.375902e-06, 1.375905e-06, 
    1.375903e-06, 1.375906e-06, 1.375915e-06, 1.375912e-06, 1.375921e-06, 
    1.375926e-06, 1.375929e-06, 1.375932e-06, 1.375931e-06, 1.375931e-06, 
    1.375927e-06, 1.375924e-06, 1.375922e-06, 1.37592e-06, 1.375919e-06, 
    1.375914e-06, 1.375912e-06, 1.375906e-06, 1.375907e-06, 1.375905e-06, 
    1.375904e-06, 1.375901e-06, 1.375901e-06, 1.3759e-06, 1.375905e-06, 
    1.375902e-06, 1.375908e-06, 1.375906e-06, 1.375918e-06, 1.375923e-06, 
    1.375925e-06, 1.375927e-06, 1.375931e-06, 1.375928e-06, 1.375929e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.37592e-06, 1.375922e-06, 
    1.375911e-06, 1.375916e-06, 1.375904e-06, 1.375907e-06, 1.375903e-06, 
    1.375905e-06, 1.375902e-06, 1.375905e-06, 1.3759e-06, 1.375899e-06, 
    1.375899e-06, 1.375897e-06, 1.375905e-06, 1.375902e-06, 1.375926e-06, 
    1.375926e-06, 1.375925e-06, 1.375928e-06, 1.375928e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.375922e-06, 
    1.375919e-06, 1.375915e-06, 1.37591e-06, 1.375907e-06, 1.375904e-06, 
    1.375906e-06, 1.375905e-06, 1.375906e-06, 1.375907e-06, 1.375899e-06, 
    1.375903e-06, 1.375897e-06, 1.375897e-06, 1.3759e-06, 1.375897e-06, 
    1.375926e-06, 1.375926e-06, 1.375929e-06, 1.375927e-06, 1.375931e-06, 
    1.375929e-06, 1.375927e-06, 1.375922e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375916e-06, 1.375911e-06, 1.375907e-06, 1.375904e-06, 
    1.375904e-06, 1.375904e-06, 1.375903e-06, 1.375905e-06, 1.375903e-06, 
    1.375902e-06, 1.375903e-06, 1.375897e-06, 1.375899e-06, 1.375897e-06, 
    1.375898e-06, 1.375926e-06, 1.375925e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.375921e-06, 1.375919e-06, 1.375913e-06, 1.375916e-06, 
    1.375912e-06, 1.375915e-06, 1.375915e-06, 1.375912e-06, 1.375915e-06, 
    1.375907e-06, 1.375913e-06, 1.375903e-06, 1.375908e-06, 1.375903e-06, 
    1.375904e-06, 1.375902e-06, 1.375901e-06, 1.375899e-06, 1.375895e-06, 
    1.375896e-06, 1.375893e-06, 1.375923e-06, 1.375921e-06, 1.375921e-06, 
    1.375919e-06, 1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375912e-06, 
    1.375908e-06, 1.375908e-06, 1.375913e-06, 1.37591e-06, 1.37592e-06, 
    1.375918e-06, 1.375919e-06, 1.375922e-06, 1.375911e-06, 1.375917e-06, 
    1.375907e-06, 1.37591e-06, 1.375901e-06, 1.375905e-06, 1.375896e-06, 
    1.375893e-06, 1.375889e-06, 1.375885e-06, 1.37592e-06, 1.375921e-06, 
    1.375919e-06, 1.375916e-06, 1.375913e-06, 1.37591e-06, 1.375909e-06, 
    1.375908e-06, 1.375907e-06, 1.375905e-06, 1.375908e-06, 1.375905e-06, 
    1.375918e-06, 1.375911e-06, 1.375922e-06, 1.375918e-06, 1.375916e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375894e-06, 1.3759e-06, 1.375882e-06, 1.375887e-06, 1.375922e-06, 
    1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 1.375907e-06, 
    1.375906e-06, 1.375904e-06, 1.375904e-06, 1.375902e-06, 1.375904e-06, 
    1.375903e-06, 1.37591e-06, 1.375906e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375908e-06, 
    1.375907e-06, 1.375904e-06, 1.375909e-06, 1.375893e-06, 1.375903e-06, 
    1.375918e-06, 1.375915e-06, 1.375915e-06, 1.375916e-06, 1.375908e-06, 
    1.375911e-06, 1.375902e-06, 1.375905e-06, 1.375901e-06, 1.375903e-06, 
    1.375903e-06, 1.375905e-06, 1.375907e-06, 1.37591e-06, 1.375913e-06, 
    1.375916e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.375905e-06, 1.375901e-06, 1.37591e-06, 1.375906e-06, 1.375908e-06, 
    1.375904e-06, 1.375912e-06, 1.375905e-06, 1.375914e-06, 1.375913e-06, 
    1.375911e-06, 1.375906e-06, 1.375905e-06, 1.375904e-06, 1.375905e-06, 
    1.375908e-06, 1.375908e-06, 1.375911e-06, 1.375911e-06, 1.375913e-06, 
    1.375914e-06, 1.375913e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.3759e-06, 1.3759e-06, 1.375895e-06, 1.375899e-06, 1.375893e-06, 
    1.375898e-06, 1.375889e-06, 1.375905e-06, 1.375898e-06, 1.37591e-06, 
    1.375909e-06, 1.375907e-06, 1.375901e-06, 1.375904e-06, 1.375901e-06, 
    1.375908e-06, 1.375912e-06, 1.375913e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375912e-06, 1.375912e-06, 1.375908e-06, 1.37591e-06, 
    1.375903e-06, 1.375901e-06, 1.375893e-06, 1.375889e-06, 1.375884e-06, 
    1.375883e-06, 1.375882e-06, 1.375882e-06 ;

 TOTLITN_1m =
  1.37593e-06, 1.375926e-06, 1.375927e-06, 1.375924e-06, 1.375926e-06, 
    1.375923e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 1.37593e-06, 
    1.375917e-06, 1.375924e-06, 1.375911e-06, 1.375915e-06, 1.375905e-06, 
    1.375911e-06, 1.375903e-06, 1.375905e-06, 1.3759e-06, 1.375902e-06, 
    1.375896e-06, 1.3759e-06, 1.375893e-06, 1.375897e-06, 1.375896e-06, 
    1.3759e-06, 1.375922e-06, 1.375918e-06, 1.375923e-06, 1.375922e-06, 
    1.375922e-06, 1.375926e-06, 1.375927e-06, 1.375931e-06, 1.37593e-06, 
    1.375927e-06, 1.375922e-06, 1.375924e-06, 1.375919e-06, 1.375919e-06, 
    1.375913e-06, 1.375916e-06, 1.375907e-06, 1.375909e-06, 1.375902e-06, 
    1.375903e-06, 1.375902e-06, 1.375902e-06, 1.375902e-06, 1.375905e-06, 
    1.375903e-06, 1.375906e-06, 1.375915e-06, 1.375912e-06, 1.375921e-06, 
    1.375926e-06, 1.375929e-06, 1.375932e-06, 1.375931e-06, 1.375931e-06, 
    1.375927e-06, 1.375924e-06, 1.375922e-06, 1.37592e-06, 1.375919e-06, 
    1.375914e-06, 1.375912e-06, 1.375906e-06, 1.375907e-06, 1.375905e-06, 
    1.375904e-06, 1.375901e-06, 1.375901e-06, 1.3759e-06, 1.375905e-06, 
    1.375902e-06, 1.375908e-06, 1.375906e-06, 1.375918e-06, 1.375923e-06, 
    1.375925e-06, 1.375927e-06, 1.375931e-06, 1.375928e-06, 1.375929e-06, 
    1.375927e-06, 1.375925e-06, 1.375926e-06, 1.37592e-06, 1.375922e-06, 
    1.375911e-06, 1.375916e-06, 1.375904e-06, 1.375907e-06, 1.375903e-06, 
    1.375905e-06, 1.375902e-06, 1.375905e-06, 1.3759e-06, 1.375899e-06, 
    1.375899e-06, 1.375897e-06, 1.375905e-06, 1.375902e-06, 1.375926e-06, 
    1.375926e-06, 1.375925e-06, 1.375928e-06, 1.375928e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.375922e-06, 
    1.375919e-06, 1.375915e-06, 1.37591e-06, 1.375907e-06, 1.375904e-06, 
    1.375906e-06, 1.375905e-06, 1.375906e-06, 1.375907e-06, 1.375899e-06, 
    1.375903e-06, 1.375897e-06, 1.375897e-06, 1.3759e-06, 1.375897e-06, 
    1.375926e-06, 1.375926e-06, 1.375929e-06, 1.375927e-06, 1.375931e-06, 
    1.375929e-06, 1.375927e-06, 1.375922e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375916e-06, 1.375911e-06, 1.375907e-06, 1.375904e-06, 
    1.375904e-06, 1.375904e-06, 1.375903e-06, 1.375905e-06, 1.375903e-06, 
    1.375902e-06, 1.375903e-06, 1.375897e-06, 1.375899e-06, 1.375897e-06, 
    1.375898e-06, 1.375926e-06, 1.375925e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.375921e-06, 1.375919e-06, 1.375913e-06, 1.375916e-06, 
    1.375912e-06, 1.375915e-06, 1.375915e-06, 1.375912e-06, 1.375915e-06, 
    1.375907e-06, 1.375913e-06, 1.375903e-06, 1.375908e-06, 1.375903e-06, 
    1.375904e-06, 1.375902e-06, 1.375901e-06, 1.375899e-06, 1.375895e-06, 
    1.375896e-06, 1.375893e-06, 1.375923e-06, 1.375921e-06, 1.375921e-06, 
    1.375919e-06, 1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375912e-06, 
    1.375908e-06, 1.375908e-06, 1.375913e-06, 1.37591e-06, 1.37592e-06, 
    1.375918e-06, 1.375919e-06, 1.375922e-06, 1.375911e-06, 1.375917e-06, 
    1.375907e-06, 1.37591e-06, 1.375901e-06, 1.375905e-06, 1.375896e-06, 
    1.375893e-06, 1.375889e-06, 1.375885e-06, 1.37592e-06, 1.375921e-06, 
    1.375919e-06, 1.375916e-06, 1.375913e-06, 1.37591e-06, 1.375909e-06, 
    1.375908e-06, 1.375907e-06, 1.375905e-06, 1.375908e-06, 1.375905e-06, 
    1.375918e-06, 1.375911e-06, 1.375922e-06, 1.375918e-06, 1.375916e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375894e-06, 1.3759e-06, 1.375882e-06, 1.375887e-06, 1.375922e-06, 
    1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 1.375907e-06, 
    1.375906e-06, 1.375904e-06, 1.375904e-06, 1.375902e-06, 1.375904e-06, 
    1.375903e-06, 1.37591e-06, 1.375906e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375908e-06, 
    1.375907e-06, 1.375904e-06, 1.375909e-06, 1.375893e-06, 1.375903e-06, 
    1.375918e-06, 1.375915e-06, 1.375915e-06, 1.375916e-06, 1.375908e-06, 
    1.375911e-06, 1.375902e-06, 1.375905e-06, 1.375901e-06, 1.375903e-06, 
    1.375903e-06, 1.375905e-06, 1.375907e-06, 1.37591e-06, 1.375913e-06, 
    1.375916e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.375905e-06, 1.375901e-06, 1.37591e-06, 1.375906e-06, 1.375908e-06, 
    1.375904e-06, 1.375912e-06, 1.375905e-06, 1.375914e-06, 1.375913e-06, 
    1.375911e-06, 1.375906e-06, 1.375905e-06, 1.375904e-06, 1.375905e-06, 
    1.375908e-06, 1.375908e-06, 1.375911e-06, 1.375911e-06, 1.375913e-06, 
    1.375914e-06, 1.375913e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.3759e-06, 1.3759e-06, 1.375895e-06, 1.375899e-06, 1.375893e-06, 
    1.375898e-06, 1.375889e-06, 1.375905e-06, 1.375898e-06, 1.37591e-06, 
    1.375909e-06, 1.375907e-06, 1.375901e-06, 1.375904e-06, 1.375901e-06, 
    1.375908e-06, 1.375912e-06, 1.375913e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375912e-06, 1.375912e-06, 1.375908e-06, 1.37591e-06, 
    1.375903e-06, 1.375901e-06, 1.375893e-06, 1.375889e-06, 1.375884e-06, 
    1.375883e-06, 1.375882e-06, 1.375882e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773745, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773748, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773737, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.773751, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773745, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773748, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773737, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.773751, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  243.0869, 243.0901, 243.0895, 243.0921, 243.0907, 243.0923, 243.0875, 
    243.0902, 243.0885, 243.0872, 243.097, 243.0922, 243.1021, 243.0991, 
    243.1068, 243.1016, 243.1079, 243.1067, 243.1103, 243.1093, 243.1137, 
    243.1108, 243.1161, 243.1131, 243.1135, 243.1107, 243.0932, 243.0963, 
    243.093, 243.0934, 243.0933, 243.0907, 243.0893, 243.0866, 243.0871, 
    243.0891, 243.0937, 243.0921, 243.096, 243.0959, 243.1002, 243.0983, 
    243.1055, 243.1035, 243.1093, 243.1078, 243.1092, 243.1088, 243.1093, 
    243.1071, 243.108, 243.1061, 243.0986, 243.1008, 243.0943, 243.0902, 
    243.0876, 243.0858, 243.086, 243.0865, 243.0891, 243.0916, 243.0935, 
    243.0947, 243.0959, 243.0995, 243.1015, 243.1059, 243.1051, 243.1064, 
    243.1077, 243.1098, 243.1095, 243.1104, 243.1064, 243.109, 243.1047, 
    243.1059, 243.0961, 243.0926, 243.0909, 243.0896, 243.0862, 243.0885, 
    243.0876, 243.0898, 243.0912, 243.0905, 243.0947, 243.0931, 243.1016, 
    243.098, 243.1075, 243.1053, 243.1081, 243.1067, 243.1091, 243.1069, 
    243.1107, 243.1115, 243.111, 243.1132, 243.1068, 243.1092, 243.0905, 
    243.0906, 243.0912, 243.0888, 243.0887, 243.0866, 243.0885, 243.0893, 
    243.0913, 243.0925, 243.0936, 243.0961, 243.0988, 243.1026, 243.1054, 
    243.1073, 243.1061, 243.1071, 243.106, 243.1055, 243.1112, 243.108, 
    243.1129, 243.1126, 243.1104, 243.1126, 243.0907, 243.0901, 243.0878, 
    243.0896, 243.0864, 243.0882, 243.0892, 243.0931, 243.094, 243.0948, 
    243.0964, 243.0984, 243.1019, 243.105, 243.1078, 243.1076, 243.1076, 
    243.1082, 243.1067, 243.1085, 243.1088, 243.108, 243.1126, 243.1113, 
    243.1126, 243.1118, 243.0903, 243.0914, 243.0908, 243.0918, 243.0911, 
    243.0945, 243.0955, 243.1003, 243.0983, 243.1014, 243.0987, 243.0992, 
    243.1015, 243.0988, 243.1048, 243.1007, 243.1083, 243.1041, 243.1085, 
    243.1078, 243.1091, 243.1102, 243.1116, 243.1143, 243.1137, 243.1159, 
    243.093, 243.0943, 243.0942, 243.0957, 243.0967, 243.0991, 243.1028, 
    243.1014, 243.104, 243.1045, 243.1006, 243.103, 243.0953, 243.0965, 
    243.0958, 243.093, 243.1017, 243.0972, 243.1055, 243.1031, 243.11, 
    243.1065, 243.1133, 243.1161, 243.1189, 243.122, 243.0951, 243.0942, 
    243.0959, 243.0981, 243.1003, 243.1032, 243.1035, 243.104, 243.1054, 
    243.1066, 243.1042, 243.1069, 243.0967, 243.1021, 243.0938, 243.0963, 
    243.098, 243.0973, 243.1013, 243.1022, 243.1059, 243.104, 243.1154, 
    243.1104, 243.1244, 243.1205, 243.0938, 243.0951, 243.0995, 243.0974, 
    243.1034, 243.1049, 243.1061, 243.1076, 243.1078, 243.1086, 243.1072, 
    243.1086, 243.1032, 243.1056, 243.099, 243.1006, 243.0999, 243.0991, 
    243.1016, 243.1042, 243.1043, 243.1051, 243.1074, 243.1034, 243.116, 
    243.1082, 243.0965, 243.0989, 243.0993, 243.0983, 243.1047, 243.1024, 
    243.1086, 243.107, 243.1097, 243.1083, 243.1081, 243.1064, 243.1053, 
    243.1025, 243.1003, 243.0985, 243.0989, 243.1008, 243.1044, 243.1077, 
    243.107, 243.1095, 243.103, 243.1057, 243.1046, 243.1074, 243.1014, 
    243.1063, 243.1001, 243.1006, 243.1024, 243.1058, 243.1067, 243.1075, 
    243.107, 243.1045, 243.1041, 243.1023, 243.1018, 243.1005, 243.0994, 
    243.1004, 243.1014, 243.1045, 243.1072, 243.1102, 243.1109, 243.1143, 
    243.1115, 243.116, 243.112, 243.1189, 243.1067, 243.112, 243.1025, 
    243.1035, 243.1053, 243.1097, 243.1074, 243.1101, 243.1041, 243.1009, 
    243.1001, 243.0986, 243.1002, 243.1, 243.1015, 243.101, 243.1046, 
    243.1027, 243.1081, 243.1101, 243.1156, 243.119, 243.1225, 243.124, 
    243.1245, 243.1246 ;

 TREFMNAV_R =
  243.0869, 243.0901, 243.0895, 243.0921, 243.0907, 243.0923, 243.0875, 
    243.0902, 243.0885, 243.0872, 243.097, 243.0922, 243.1021, 243.0991, 
    243.1068, 243.1016, 243.1079, 243.1067, 243.1103, 243.1093, 243.1137, 
    243.1108, 243.1161, 243.1131, 243.1135, 243.1107, 243.0932, 243.0963, 
    243.093, 243.0934, 243.0933, 243.0907, 243.0893, 243.0866, 243.0871, 
    243.0891, 243.0937, 243.0921, 243.096, 243.0959, 243.1002, 243.0983, 
    243.1055, 243.1035, 243.1093, 243.1078, 243.1092, 243.1088, 243.1093, 
    243.1071, 243.108, 243.1061, 243.0986, 243.1008, 243.0943, 243.0902, 
    243.0876, 243.0858, 243.086, 243.0865, 243.0891, 243.0916, 243.0935, 
    243.0947, 243.0959, 243.0995, 243.1015, 243.1059, 243.1051, 243.1064, 
    243.1077, 243.1098, 243.1095, 243.1104, 243.1064, 243.109, 243.1047, 
    243.1059, 243.0961, 243.0926, 243.0909, 243.0896, 243.0862, 243.0885, 
    243.0876, 243.0898, 243.0912, 243.0905, 243.0947, 243.0931, 243.1016, 
    243.098, 243.1075, 243.1053, 243.1081, 243.1067, 243.1091, 243.1069, 
    243.1107, 243.1115, 243.111, 243.1132, 243.1068, 243.1092, 243.0905, 
    243.0906, 243.0912, 243.0888, 243.0887, 243.0866, 243.0885, 243.0893, 
    243.0913, 243.0925, 243.0936, 243.0961, 243.0988, 243.1026, 243.1054, 
    243.1073, 243.1061, 243.1071, 243.106, 243.1055, 243.1112, 243.108, 
    243.1129, 243.1126, 243.1104, 243.1126, 243.0907, 243.0901, 243.0878, 
    243.0896, 243.0864, 243.0882, 243.0892, 243.0931, 243.094, 243.0948, 
    243.0964, 243.0984, 243.1019, 243.105, 243.1078, 243.1076, 243.1076, 
    243.1082, 243.1067, 243.1085, 243.1088, 243.108, 243.1126, 243.1113, 
    243.1126, 243.1118, 243.0903, 243.0914, 243.0908, 243.0918, 243.0911, 
    243.0945, 243.0955, 243.1003, 243.0983, 243.1014, 243.0987, 243.0992, 
    243.1015, 243.0988, 243.1048, 243.1007, 243.1083, 243.1041, 243.1085, 
    243.1078, 243.1091, 243.1102, 243.1116, 243.1143, 243.1137, 243.1159, 
    243.093, 243.0943, 243.0942, 243.0957, 243.0967, 243.0991, 243.1028, 
    243.1014, 243.104, 243.1045, 243.1006, 243.103, 243.0953, 243.0965, 
    243.0958, 243.093, 243.1017, 243.0972, 243.1055, 243.1031, 243.11, 
    243.1065, 243.1133, 243.1161, 243.1189, 243.122, 243.0951, 243.0942, 
    243.0959, 243.0981, 243.1003, 243.1032, 243.1035, 243.104, 243.1054, 
    243.1066, 243.1042, 243.1069, 243.0967, 243.1021, 243.0938, 243.0963, 
    243.098, 243.0973, 243.1013, 243.1022, 243.1059, 243.104, 243.1154, 
    243.1104, 243.1244, 243.1205, 243.0938, 243.0951, 243.0995, 243.0974, 
    243.1034, 243.1049, 243.1061, 243.1076, 243.1078, 243.1086, 243.1072, 
    243.1086, 243.1032, 243.1056, 243.099, 243.1006, 243.0999, 243.0991, 
    243.1016, 243.1042, 243.1043, 243.1051, 243.1074, 243.1034, 243.116, 
    243.1082, 243.0965, 243.0989, 243.0993, 243.0983, 243.1047, 243.1024, 
    243.1086, 243.107, 243.1097, 243.1083, 243.1081, 243.1064, 243.1053, 
    243.1025, 243.1003, 243.0985, 243.0989, 243.1008, 243.1044, 243.1077, 
    243.107, 243.1095, 243.103, 243.1057, 243.1046, 243.1074, 243.1014, 
    243.1063, 243.1001, 243.1006, 243.1024, 243.1058, 243.1067, 243.1075, 
    243.107, 243.1045, 243.1041, 243.1023, 243.1018, 243.1005, 243.0994, 
    243.1004, 243.1014, 243.1045, 243.1072, 243.1102, 243.1109, 243.1143, 
    243.1115, 243.116, 243.112, 243.1189, 243.1067, 243.112, 243.1025, 
    243.1035, 243.1053, 243.1097, 243.1074, 243.1101, 243.1041, 243.1009, 
    243.1001, 243.0986, 243.1002, 243.1, 243.1015, 243.101, 243.1046, 
    243.1027, 243.1081, 243.1101, 243.1156, 243.119, 243.1225, 243.124, 
    243.1245, 243.1246 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7644, 270.7623, 270.7627, 270.761, 270.7619, 270.7608, 270.7639, 
    270.7622, 270.7633, 270.7642, 270.7578, 270.7609, 270.7544, 270.7564, 
    270.7513, 270.7547, 270.7506, 270.7513, 270.749, 270.7496, 270.7467, 
    270.7486, 270.7451, 270.7471, 270.7468, 270.7487, 270.7603, 270.7582, 
    270.7604, 270.7601, 270.7602, 270.7619, 270.7628, 270.7645, 270.7642, 
    270.7629, 270.7599, 270.7609, 270.7584, 270.7585, 270.7556, 270.7569, 
    270.7522, 270.7535, 270.7496, 270.7506, 270.7497, 270.7499, 270.7497, 
    270.7511, 270.7505, 270.7517, 270.7567, 270.7552, 270.7596, 270.7622, 
    270.7639, 270.7651, 270.7649, 270.7646, 270.7629, 270.7613, 270.7601, 
    270.7593, 270.7585, 270.7561, 270.7548, 270.7519, 270.7524, 270.7516, 
    270.7507, 270.7493, 270.7495, 270.7489, 270.7516, 270.7498, 270.7527, 
    270.7519, 270.7584, 270.7607, 270.7617, 270.7626, 270.7648, 270.7633, 
    270.7639, 270.7625, 270.7616, 270.762, 270.7592, 270.7603, 270.7547, 
    270.7571, 270.7508, 270.7523, 270.7504, 270.7514, 270.7498, 270.7512, 
    270.7487, 270.7481, 270.7485, 270.747, 270.7513, 270.7497, 270.762, 
    270.7619, 270.7616, 270.7631, 270.7632, 270.7646, 270.7633, 270.7628, 
    270.7615, 270.7607, 270.76, 270.7584, 270.7566, 270.7541, 270.7522, 
    270.751, 270.7517, 270.7511, 270.7518, 270.7521, 270.7484, 270.7505, 
    270.7473, 270.7474, 270.7489, 270.7474, 270.7619, 270.7623, 270.7638, 
    270.7626, 270.7647, 270.7635, 270.7629, 270.7603, 270.7597, 270.7592, 
    270.7582, 270.7568, 270.7545, 270.7525, 270.7506, 270.7508, 270.7507, 
    270.7503, 270.7513, 270.7502, 270.75, 270.7505, 270.7474, 270.7483, 
    270.7474, 270.748, 270.7621, 270.7615, 270.7618, 270.7611, 270.7617, 
    270.7594, 270.7588, 270.7556, 270.7569, 270.7549, 270.7567, 270.7563, 
    270.7549, 270.7566, 270.7527, 270.7553, 270.7503, 270.7531, 270.7501, 
    270.7506, 270.7498, 270.749, 270.748, 270.7463, 270.7467, 270.7452, 
    270.7604, 270.7595, 270.7596, 270.7586, 270.7579, 270.7564, 270.7539, 
    270.7549, 270.7531, 270.7528, 270.7554, 270.7538, 270.7589, 270.7581, 
    270.7586, 270.7603, 270.7547, 270.7576, 270.7522, 270.7538, 270.7491, 
    270.7515, 270.7469, 270.7451, 270.7432, 270.7411, 270.759, 270.7596, 
    270.7585, 270.757, 270.7556, 270.7537, 270.7534, 270.7531, 270.7522, 
    270.7514, 270.753, 270.7512, 270.758, 270.7544, 270.7599, 270.7583, 
    270.7571, 270.7576, 270.7549, 270.7543, 270.7519, 270.7531, 270.7455, 
    270.7489, 270.7395, 270.7421, 270.7598, 270.759, 270.7561, 270.7575, 
    270.7535, 270.7526, 270.7518, 270.7508, 270.7506, 270.7501, 270.751, 
    270.7501, 270.7537, 270.7521, 270.7564, 270.7554, 270.7559, 270.7564, 
    270.7547, 270.753, 270.7529, 270.7524, 270.7509, 270.7535, 270.7452, 
    270.7504, 270.7581, 270.7565, 270.7563, 270.7569, 270.7527, 270.7542, 
    270.7501, 270.7512, 270.7494, 270.7503, 270.7504, 270.7516, 270.7523, 
    270.7541, 270.7556, 270.7568, 270.7565, 270.7552, 270.7529, 270.7506, 
    270.7512, 270.7495, 270.7538, 270.752, 270.7527, 270.7509, 270.7549, 
    270.7516, 270.7557, 270.7554, 270.7542, 270.7519, 270.7514, 270.7508, 
    270.7512, 270.7528, 270.7531, 270.7542, 270.7546, 270.7555, 270.7562, 
    270.7555, 270.7548, 270.7528, 270.751, 270.749, 270.7485, 270.7463, 
    270.7482, 270.7452, 270.7478, 270.7432, 270.7513, 270.7478, 270.7542, 
    270.7534, 270.7523, 270.7494, 270.7509, 270.7491, 270.7531, 270.7552, 
    270.7557, 270.7567, 270.7557, 270.7558, 270.7548, 270.7551, 270.7527, 
    270.754, 270.7504, 270.7491, 270.7454, 270.7431, 270.7408, 270.7397, 
    270.7394, 270.7393 ;

 TREFMXAV_R =
  270.7644, 270.7623, 270.7627, 270.761, 270.7619, 270.7608, 270.7639, 
    270.7622, 270.7633, 270.7642, 270.7578, 270.7609, 270.7544, 270.7564, 
    270.7513, 270.7547, 270.7506, 270.7513, 270.749, 270.7496, 270.7467, 
    270.7486, 270.7451, 270.7471, 270.7468, 270.7487, 270.7603, 270.7582, 
    270.7604, 270.7601, 270.7602, 270.7619, 270.7628, 270.7645, 270.7642, 
    270.7629, 270.7599, 270.7609, 270.7584, 270.7585, 270.7556, 270.7569, 
    270.7522, 270.7535, 270.7496, 270.7506, 270.7497, 270.7499, 270.7497, 
    270.7511, 270.7505, 270.7517, 270.7567, 270.7552, 270.7596, 270.7622, 
    270.7639, 270.7651, 270.7649, 270.7646, 270.7629, 270.7613, 270.7601, 
    270.7593, 270.7585, 270.7561, 270.7548, 270.7519, 270.7524, 270.7516, 
    270.7507, 270.7493, 270.7495, 270.7489, 270.7516, 270.7498, 270.7527, 
    270.7519, 270.7584, 270.7607, 270.7617, 270.7626, 270.7648, 270.7633, 
    270.7639, 270.7625, 270.7616, 270.762, 270.7592, 270.7603, 270.7547, 
    270.7571, 270.7508, 270.7523, 270.7504, 270.7514, 270.7498, 270.7512, 
    270.7487, 270.7481, 270.7485, 270.747, 270.7513, 270.7497, 270.762, 
    270.7619, 270.7616, 270.7631, 270.7632, 270.7646, 270.7633, 270.7628, 
    270.7615, 270.7607, 270.76, 270.7584, 270.7566, 270.7541, 270.7522, 
    270.751, 270.7517, 270.7511, 270.7518, 270.7521, 270.7484, 270.7505, 
    270.7473, 270.7474, 270.7489, 270.7474, 270.7619, 270.7623, 270.7638, 
    270.7626, 270.7647, 270.7635, 270.7629, 270.7603, 270.7597, 270.7592, 
    270.7582, 270.7568, 270.7545, 270.7525, 270.7506, 270.7508, 270.7507, 
    270.7503, 270.7513, 270.7502, 270.75, 270.7505, 270.7474, 270.7483, 
    270.7474, 270.748, 270.7621, 270.7615, 270.7618, 270.7611, 270.7617, 
    270.7594, 270.7588, 270.7556, 270.7569, 270.7549, 270.7567, 270.7563, 
    270.7549, 270.7566, 270.7527, 270.7553, 270.7503, 270.7531, 270.7501, 
    270.7506, 270.7498, 270.749, 270.748, 270.7463, 270.7467, 270.7452, 
    270.7604, 270.7595, 270.7596, 270.7586, 270.7579, 270.7564, 270.7539, 
    270.7549, 270.7531, 270.7528, 270.7554, 270.7538, 270.7589, 270.7581, 
    270.7586, 270.7603, 270.7547, 270.7576, 270.7522, 270.7538, 270.7491, 
    270.7515, 270.7469, 270.7451, 270.7432, 270.7411, 270.759, 270.7596, 
    270.7585, 270.757, 270.7556, 270.7537, 270.7534, 270.7531, 270.7522, 
    270.7514, 270.753, 270.7512, 270.758, 270.7544, 270.7599, 270.7583, 
    270.7571, 270.7576, 270.7549, 270.7543, 270.7519, 270.7531, 270.7455, 
    270.7489, 270.7395, 270.7421, 270.7598, 270.759, 270.7561, 270.7575, 
    270.7535, 270.7526, 270.7518, 270.7508, 270.7506, 270.7501, 270.751, 
    270.7501, 270.7537, 270.7521, 270.7564, 270.7554, 270.7559, 270.7564, 
    270.7547, 270.753, 270.7529, 270.7524, 270.7509, 270.7535, 270.7452, 
    270.7504, 270.7581, 270.7565, 270.7563, 270.7569, 270.7527, 270.7542, 
    270.7501, 270.7512, 270.7494, 270.7503, 270.7504, 270.7516, 270.7523, 
    270.7541, 270.7556, 270.7568, 270.7565, 270.7552, 270.7529, 270.7506, 
    270.7512, 270.7495, 270.7538, 270.752, 270.7527, 270.7509, 270.7549, 
    270.7516, 270.7557, 270.7554, 270.7542, 270.7519, 270.7514, 270.7508, 
    270.7512, 270.7528, 270.7531, 270.7542, 270.7546, 270.7555, 270.7562, 
    270.7555, 270.7548, 270.7528, 270.751, 270.749, 270.7485, 270.7463, 
    270.7482, 270.7452, 270.7478, 270.7432, 270.7513, 270.7478, 270.7542, 
    270.7534, 270.7523, 270.7494, 270.7509, 270.7491, 270.7531, 270.7552, 
    270.7557, 270.7567, 270.7557, 270.7558, 270.7548, 270.7551, 270.7527, 
    270.754, 270.7504, 270.7491, 270.7454, 270.7431, 270.7408, 270.7397, 
    270.7394, 270.7393 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.2031, 255.203, 255.203, 255.2029, 255.203, 255.2029, 255.2031, 255.203, 
    255.2031, 255.2031, 255.2027, 255.2029, 255.2024, 255.2026, 255.2022, 
    255.2024, 255.2021, 255.2022, 255.202, 255.2021, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2018, 255.202, 255.2029, 255.2027, 255.2029, 
    255.2028, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.203, 
    255.2028, 255.2029, 255.2027, 255.2027, 255.2025, 255.2026, 255.2023, 
    255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2021, 255.2022, 255.2026, 255.2025, 255.2028, 255.203, 255.2031, 
    255.2032, 255.2032, 255.2032, 255.203, 255.2029, 255.2028, 255.2028, 
    255.2027, 255.2025, 255.2025, 255.2022, 255.2023, 255.2022, 255.2021, 
    255.202, 255.2021, 255.202, 255.2022, 255.2021, 255.2023, 255.2022, 
    255.2027, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.2031, 
    255.203, 255.2029, 255.203, 255.2028, 255.2029, 255.2024, 255.2026, 
    255.2021, 255.2023, 255.2021, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.203, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2022, 255.2022, 255.2022, 255.2023, 255.202, 255.2021, 255.2019, 
    255.2019, 255.202, 255.2019, 255.203, 255.203, 255.2031, 255.203, 
    255.2032, 255.2031, 255.203, 255.2029, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 
    255.2022, 255.2021, 255.2021, 255.2021, 255.2019, 255.202, 255.2019, 
    255.2019, 255.203, 255.2029, 255.203, 255.2029, 255.2029, 255.2028, 
    255.2027, 255.2025, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 
    255.2026, 255.2023, 255.2025, 255.2021, 255.2023, 255.2021, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2018, 255.2018, 255.2017, 255.2029, 
    255.2028, 255.2028, 255.2027, 255.2027, 255.2026, 255.2024, 255.2025, 
    255.2023, 255.2023, 255.2025, 255.2024, 255.2027, 255.2027, 255.2027, 
    255.2029, 255.2024, 255.2027, 255.2023, 255.2024, 255.202, 255.2022, 
    255.2019, 255.2017, 255.2016, 255.2014, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2025, 255.2024, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2027, 255.2024, 255.2028, 255.2027, 255.2026, 
    255.2027, 255.2025, 255.2024, 255.2022, 255.2023, 255.2018, 255.202, 
    255.2013, 255.2015, 255.2028, 255.2028, 255.2025, 255.2027, 255.2023, 
    255.2023, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 255.2021, 
    255.2024, 255.2022, 255.2026, 255.2025, 255.2025, 255.2026, 255.2024, 
    255.2023, 255.2023, 255.2023, 255.2022, 255.2023, 255.2017, 255.2021, 
    255.2027, 255.2026, 255.2026, 255.2026, 255.2023, 255.2024, 255.2021, 
    255.2022, 255.202, 255.2021, 255.2021, 255.2022, 255.2023, 255.2024, 
    255.2025, 255.2026, 255.2026, 255.2025, 255.2023, 255.2021, 255.2022, 
    255.2021, 255.2024, 255.2022, 255.2023, 255.2021, 255.2025, 255.2022, 
    255.2025, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 255.2022, 
    255.2023, 255.2023, 255.2024, 255.2024, 255.2025, 255.2025, 255.2025, 
    255.2025, 255.2023, 255.2022, 255.202, 255.202, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2016, 255.2022, 255.2019, 255.2024, 255.2023, 
    255.2023, 255.202, 255.2021, 255.202, 255.2023, 255.2025, 255.2025, 
    255.2026, 255.2025, 255.2025, 255.2025, 255.2025, 255.2023, 255.2024, 
    255.2021, 255.202, 255.2017, 255.2016, 255.2014, 255.2013, 255.2013, 
    255.2013 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  255.2031, 255.203, 255.203, 255.2029, 255.203, 255.2029, 255.2031, 255.203, 
    255.2031, 255.2031, 255.2027, 255.2029, 255.2024, 255.2026, 255.2022, 
    255.2024, 255.2021, 255.2022, 255.202, 255.2021, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2018, 255.202, 255.2029, 255.2027, 255.2029, 
    255.2028, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.203, 
    255.2028, 255.2029, 255.2027, 255.2027, 255.2025, 255.2026, 255.2023, 
    255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2021, 255.2022, 255.2026, 255.2025, 255.2028, 255.203, 255.2031, 
    255.2032, 255.2032, 255.2032, 255.203, 255.2029, 255.2028, 255.2028, 
    255.2027, 255.2025, 255.2025, 255.2022, 255.2023, 255.2022, 255.2021, 
    255.202, 255.2021, 255.202, 255.2022, 255.2021, 255.2023, 255.2022, 
    255.2027, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.2031, 
    255.203, 255.2029, 255.203, 255.2028, 255.2029, 255.2024, 255.2026, 
    255.2021, 255.2023, 255.2021, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.203, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2022, 255.2022, 255.2022, 255.2023, 255.202, 255.2021, 255.2019, 
    255.2019, 255.202, 255.2019, 255.203, 255.203, 255.2031, 255.203, 
    255.2032, 255.2031, 255.203, 255.2029, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 
    255.2022, 255.2021, 255.2021, 255.2021, 255.2019, 255.202, 255.2019, 
    255.2019, 255.203, 255.2029, 255.203, 255.2029, 255.2029, 255.2028, 
    255.2027, 255.2025, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 
    255.2026, 255.2023, 255.2025, 255.2021, 255.2023, 255.2021, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2018, 255.2018, 255.2017, 255.2029, 
    255.2028, 255.2028, 255.2027, 255.2027, 255.2026, 255.2024, 255.2025, 
    255.2023, 255.2023, 255.2025, 255.2024, 255.2027, 255.2027, 255.2027, 
    255.2029, 255.2024, 255.2027, 255.2023, 255.2024, 255.202, 255.2022, 
    255.2019, 255.2017, 255.2016, 255.2014, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2025, 255.2024, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2027, 255.2024, 255.2028, 255.2027, 255.2026, 
    255.2027, 255.2025, 255.2024, 255.2022, 255.2023, 255.2018, 255.202, 
    255.2013, 255.2015, 255.2028, 255.2028, 255.2025, 255.2027, 255.2023, 
    255.2023, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 255.2021, 
    255.2024, 255.2022, 255.2026, 255.2025, 255.2025, 255.2026, 255.2024, 
    255.2023, 255.2023, 255.2023, 255.2022, 255.2023, 255.2017, 255.2021, 
    255.2027, 255.2026, 255.2026, 255.2026, 255.2023, 255.2024, 255.2021, 
    255.2022, 255.202, 255.2021, 255.2021, 255.2022, 255.2023, 255.2024, 
    255.2025, 255.2026, 255.2026, 255.2025, 255.2023, 255.2021, 255.2022, 
    255.2021, 255.2024, 255.2022, 255.2023, 255.2021, 255.2025, 255.2022, 
    255.2025, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 255.2022, 
    255.2023, 255.2023, 255.2024, 255.2024, 255.2025, 255.2025, 255.2025, 
    255.2025, 255.2023, 255.2022, 255.202, 255.202, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2016, 255.2022, 255.2019, 255.2024, 255.2023, 
    255.2023, 255.202, 255.2021, 255.202, 255.2023, 255.2025, 255.2025, 
    255.2026, 255.2025, 255.2025, 255.2025, 255.2025, 255.2023, 255.2024, 
    255.2021, 255.202, 255.2017, 255.2016, 255.2014, 255.2013, 255.2013, 
    255.2013 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6895, 253.6914, 253.691, 253.6926, 253.6917, 253.6927, 253.6899, 
    253.6915, 253.6905, 253.6897, 253.6955, 253.6926, 253.6985, 253.6967, 
    253.7013, 253.6982, 253.702, 253.7013, 253.7034, 253.7028, 253.7055, 
    253.7037, 253.707, 253.7051, 253.7054, 253.7037, 253.6932, 253.6951, 
    253.6931, 253.6934, 253.6933, 253.6917, 253.6909, 253.6894, 253.6897, 
    253.6908, 253.6935, 253.6926, 253.6949, 253.6949, 253.6974, 253.6963, 
    253.7005, 253.6993, 253.7029, 253.702, 253.7028, 253.7025, 253.7028, 
    253.7015, 253.7021, 253.7009, 253.6965, 253.6978, 253.6939, 253.6915, 
    253.69, 253.6889, 253.689, 253.6893, 253.6908, 253.6923, 253.6934, 
    253.6941, 253.6949, 253.697, 253.6982, 253.7008, 253.7003, 253.7011, 
    253.7019, 253.7031, 253.7029, 253.7035, 253.7011, 253.7027, 253.7001, 
    253.7008, 253.6949, 253.6929, 253.6919, 253.6911, 253.6891, 253.6905, 
    253.69, 253.6913, 253.6921, 253.6917, 253.6942, 253.6932, 253.6982, 
    253.6961, 253.7018, 253.7004, 253.7021, 253.7012, 253.7027, 253.7014, 
    253.7037, 253.7042, 253.7038, 253.7052, 253.7013, 253.7028, 253.6917, 
    253.6917, 253.692, 253.6907, 253.6906, 253.6894, 253.6905, 253.6909, 
    253.6921, 253.6928, 253.6935, 253.6949, 253.6965, 253.6988, 253.7005, 
    253.7016, 253.7009, 253.7015, 253.7009, 253.7005, 253.704, 253.7021, 
    253.705, 253.7048, 253.7035, 253.7048, 253.6918, 253.6914, 253.6901, 
    253.6911, 253.6892, 253.6903, 253.6909, 253.6932, 253.6937, 253.6942, 
    253.6951, 253.6963, 253.6984, 253.7002, 253.7019, 253.7018, 253.7018, 
    253.7022, 253.7013, 253.7024, 253.7025, 253.7021, 253.7048, 253.704, 
    253.7048, 253.7043, 253.6915, 253.6922, 253.6918, 253.6924, 253.692, 
    253.694, 253.6946, 253.6974, 253.6963, 253.6981, 253.6965, 253.6968, 
    253.6981, 253.6966, 253.7001, 253.6977, 253.7022, 253.6997, 253.7024, 
    253.7019, 253.7027, 253.7034, 253.7042, 253.7058, 253.7055, 253.7068, 
    253.6931, 253.6939, 253.6938, 253.6947, 253.6953, 253.6967, 253.6989, 
    253.6981, 253.6996, 253.7, 253.6976, 253.699, 253.6945, 253.6952, 
    253.6948, 253.6931, 253.6983, 253.6956, 253.7005, 253.6991, 253.7033, 
    253.7012, 253.7053, 253.707, 253.7087, 253.7105, 253.6944, 253.6938, 
    253.6948, 253.6962, 253.6975, 253.6992, 253.6994, 253.6997, 253.7005, 
    253.7012, 253.6998, 253.7014, 253.6953, 253.6985, 253.6936, 253.695, 
    253.6961, 253.6957, 253.698, 253.6986, 253.7008, 253.6997, 253.7065, 
    253.7035, 253.712, 253.7096, 253.6936, 253.6944, 253.697, 253.6957, 
    253.6993, 253.7002, 253.7009, 253.7018, 253.7019, 253.7024, 253.7016, 
    253.7024, 253.6992, 253.7006, 253.6967, 253.6976, 253.6972, 253.6967, 
    253.6982, 253.6998, 253.6998, 253.7003, 253.7017, 253.6993, 253.7068, 
    253.7021, 253.6952, 253.6966, 253.6968, 253.6963, 253.7001, 253.6987, 
    253.7024, 253.7014, 253.7031, 253.7023, 253.7021, 253.7011, 253.7004, 
    253.6988, 253.6974, 253.6964, 253.6966, 253.6978, 253.6999, 253.7019, 
    253.7014, 253.703, 253.6991, 253.7007, 253.7, 253.7017, 253.6981, 
    253.701, 253.6973, 253.6976, 253.6987, 253.7007, 253.7013, 253.7017, 
    253.7015, 253.7, 253.6997, 253.6987, 253.6984, 253.6976, 253.6969, 
    253.6975, 253.6981, 253.7, 253.7016, 253.7034, 253.7038, 253.7058, 
    253.7041, 253.7069, 253.7045, 253.7086, 253.7013, 253.7045, 253.6987, 
    253.6994, 253.7005, 253.703, 253.7017, 253.7033, 253.6997, 253.6978, 
    253.6973, 253.6964, 253.6974, 253.6973, 253.6982, 253.6979, 253.7, 
    253.6989, 253.7021, 253.7033, 253.7067, 253.7087, 253.7108, 253.7118, 
    253.7121, 253.7122,
  255.2212, 255.223, 255.2226, 255.224, 255.2233, 255.2242, 255.2216, 
    255.223, 255.2221, 255.2214, 255.2267, 255.2241, 255.2296, 255.2279, 
    255.2322, 255.2293, 255.2328, 255.2322, 255.2342, 255.2336, 255.2361, 
    255.2345, 255.2375, 255.2357, 255.236, 255.2344, 255.2247, 255.2264, 
    255.2246, 255.2248, 255.2247, 255.2233, 255.2225, 255.2211, 255.2214, 
    255.2224, 255.2249, 255.2241, 255.2262, 255.2262, 255.2285, 255.2275, 
    255.2315, 255.2303, 255.2336, 255.2328, 255.2336, 255.2334, 255.2336, 
    255.2324, 255.2329, 255.2318, 255.2277, 255.2289, 255.2253, 255.223, 
    255.2216, 255.2206, 255.2208, 255.221, 255.2224, 255.2238, 255.2248, 
    255.2255, 255.2262, 255.2281, 255.2292, 255.2317, 255.2313, 255.232, 
    255.2327, 255.2339, 255.2337, 255.2342, 255.232, 255.2335, 255.231, 
    255.2317, 255.2263, 255.2243, 255.2234, 255.2227, 255.2209, 255.2221, 
    255.2216, 255.2228, 255.2236, 255.2232, 255.2255, 255.2246, 255.2293, 
    255.2273, 255.2326, 255.2314, 255.2329, 255.2321, 255.2335, 255.2323, 
    255.2344, 255.2349, 255.2346, 255.2358, 255.2322, 255.2336, 255.2232, 
    255.2233, 255.2235, 255.2223, 255.2222, 255.2211, 255.2221, 255.2225, 
    255.2236, 255.2243, 255.2249, 255.2263, 255.2278, 255.2299, 255.2314, 
    255.2325, 255.2318, 255.2324, 255.2318, 255.2315, 255.2347, 255.2329, 
    255.2356, 255.2355, 255.2342, 255.2355, 255.2233, 255.223, 255.2217, 
    255.2227, 255.221, 255.2219, 255.2225, 255.2246, 255.2251, 255.2255, 
    255.2264, 255.2275, 255.2295, 255.2312, 255.2328, 255.2327, 255.2327, 
    255.233, 255.2322, 255.2332, 255.2333, 255.2329, 255.2355, 255.2347, 
    255.2355, 255.235, 255.2231, 255.2237, 255.2233, 255.2239, 255.2235, 
    255.2254, 255.2259, 255.2286, 255.2275, 255.2292, 255.2277, 255.228, 
    255.2292, 255.2278, 255.2311, 255.2288, 255.233, 255.2307, 255.2332, 
    255.2328, 255.2335, 255.2341, 255.2349, 255.2364, 255.2361, 255.2374, 
    255.2245, 255.2253, 255.2252, 255.226, 255.2266, 255.2279, 255.23, 
    255.2292, 255.2306, 255.2309, 255.2288, 255.2301, 255.2258, 255.2265, 
    255.2261, 255.2246, 255.2294, 255.2269, 255.2315, 255.2301, 255.234, 
    255.2321, 255.2359, 255.2375, 255.2391, 255.2409, 255.2257, 255.2252, 
    255.2261, 255.2274, 255.2286, 255.2302, 255.2304, 255.2307, 255.2314, 
    255.2321, 255.2307, 255.2323, 255.2266, 255.2296, 255.225, 255.2263, 
    255.2273, 255.2269, 255.2291, 255.2296, 255.2317, 255.2307, 255.2371, 
    255.2342, 255.2423, 255.24, 255.225, 255.2257, 255.2281, 255.227, 
    255.2303, 255.2311, 255.2318, 255.2327, 255.2328, 255.2332, 255.2324, 
    255.2332, 255.2302, 255.2316, 255.2279, 255.2288, 255.2284, 255.2279, 
    255.2293, 255.2308, 255.2308, 255.2313, 255.2325, 255.2303, 255.2374, 
    255.233, 255.2265, 255.2278, 255.228, 255.2275, 255.231, 255.2298, 
    255.2332, 255.2323, 255.2338, 255.2331, 255.233, 255.232, 255.2314, 
    255.2298, 255.2286, 255.2276, 255.2278, 255.2289, 255.2309, 255.2327, 
    255.2323, 255.2337, 255.2301, 255.2316, 255.231, 255.2326, 255.2292, 
    255.2319, 255.2285, 255.2288, 255.2297, 255.2317, 255.2321, 255.2326, 
    255.2323, 255.2309, 255.2307, 255.2297, 255.2294, 255.2287, 255.2281, 
    255.2286, 255.2292, 255.2309, 255.2325, 255.2341, 255.2345, 255.2364, 
    255.2348, 255.2374, 255.2352, 255.2391, 255.2322, 255.2352, 255.2298, 
    255.2304, 255.2314, 255.2338, 255.2325, 255.2341, 255.2307, 255.2289, 
    255.2285, 255.2276, 255.2285, 255.2284, 255.2293, 255.229, 255.231, 
    255.2299, 255.233, 255.2341, 255.2372, 255.2391, 255.2412, 255.242, 
    255.2423, 255.2424,
  257.2871, 257.2885, 257.2883, 257.2894, 257.2888, 257.2895, 257.2874, 
    257.2886, 257.2879, 257.2873, 257.2916, 257.2895, 257.2939, 257.2925, 
    257.2961, 257.2937, 257.2965, 257.296, 257.2976, 257.2972, 257.2993, 
    257.2979, 257.3004, 257.2989, 257.2991, 257.2978, 257.2899, 257.2913, 
    257.2898, 257.29, 257.2899, 257.2888, 257.2882, 257.287, 257.2873, 
    257.2881, 257.2901, 257.2895, 257.2912, 257.2911, 257.2931, 257.2922, 
    257.2954, 257.2945, 257.2972, 257.2965, 257.2971, 257.297, 257.2972, 
    257.2962, 257.2966, 257.2957, 257.2924, 257.2933, 257.2904, 257.2886, 
    257.2875, 257.2867, 257.2868, 257.287, 257.2881, 257.2892, 257.29, 
    257.2906, 257.2911, 257.2927, 257.2936, 257.2956, 257.2953, 257.2959, 
    257.2964, 257.2974, 257.2973, 257.2977, 257.2959, 257.2971, 257.2951, 
    257.2956, 257.2912, 257.2896, 257.2889, 257.2883, 257.2869, 257.2879, 
    257.2875, 257.2885, 257.289, 257.2888, 257.2906, 257.2899, 257.2937, 
    257.2921, 257.2964, 257.2953, 257.2966, 257.296, 257.2971, 257.2961, 
    257.2979, 257.2982, 257.298, 257.299, 257.296, 257.2971, 257.2887, 
    257.2888, 257.289, 257.288, 257.2879, 257.287, 257.2878, 257.2882, 
    257.2891, 257.2896, 257.2901, 257.2912, 257.2924, 257.2942, 257.2954, 
    257.2963, 257.2957, 257.2962, 257.2957, 257.2954, 257.2981, 257.2966, 
    257.2989, 257.2987, 257.2977, 257.2987, 257.2888, 257.2885, 257.2876, 
    257.2883, 257.2869, 257.2877, 257.2881, 257.2899, 257.2903, 257.2906, 
    257.2914, 257.2922, 257.2938, 257.2952, 257.2965, 257.2964, 257.2964, 
    257.2967, 257.296, 257.2968, 257.297, 257.2966, 257.2987, 257.2981, 
    257.2987, 257.2983, 257.2886, 257.2891, 257.2888, 257.2893, 257.289, 
    257.2905, 257.2909, 257.2931, 257.2922, 257.2936, 257.2924, 257.2926, 
    257.2936, 257.2924, 257.2951, 257.2933, 257.2967, 257.2948, 257.2968, 
    257.2965, 257.2971, 257.2976, 257.2983, 257.2995, 257.2992, 257.3003, 
    257.2898, 257.2904, 257.2904, 257.291, 257.2915, 257.2925, 257.2942, 
    257.2936, 257.2947, 257.295, 257.2932, 257.2943, 257.2908, 257.2914, 
    257.2911, 257.2899, 257.2937, 257.2917, 257.2954, 257.2943, 257.2975, 
    257.2959, 257.2991, 257.3004, 257.3017, 257.3032, 257.2908, 257.2903, 
    257.2911, 257.2921, 257.2931, 257.2944, 257.2946, 257.2948, 257.2954, 
    257.296, 257.2948, 257.2961, 257.2915, 257.2939, 257.2902, 257.2913, 
    257.2921, 257.2917, 257.2935, 257.2939, 257.2956, 257.2948, 257.3, 
    257.2977, 257.3043, 257.3024, 257.2902, 257.2908, 257.2927, 257.2918, 
    257.2945, 257.2952, 257.2957, 257.2964, 257.2965, 257.2969, 257.2962, 
    257.2969, 257.2944, 257.2955, 257.2925, 257.2932, 257.2929, 257.2925, 
    257.2937, 257.2949, 257.2949, 257.2953, 257.2963, 257.2945, 257.3003, 
    257.2967, 257.2914, 257.2924, 257.2926, 257.2922, 257.2951, 257.294, 
    257.2969, 257.2961, 257.2974, 257.2968, 257.2967, 257.2959, 257.2953, 
    257.2941, 257.2931, 257.2923, 257.2924, 257.2933, 257.295, 257.2965, 
    257.2961, 257.2973, 257.2943, 257.2955, 257.295, 257.2963, 257.2936, 
    257.2958, 257.293, 257.2932, 257.294, 257.2956, 257.296, 257.2964, 
    257.2961, 257.295, 257.2948, 257.294, 257.2938, 257.2932, 257.2927, 
    257.2931, 257.2936, 257.295, 257.2962, 257.2976, 257.2979, 257.2995, 
    257.2982, 257.3003, 257.2985, 257.3017, 257.296, 257.2985, 257.2941, 
    257.2946, 257.2954, 257.2974, 257.2963, 257.2975, 257.2948, 257.2934, 
    257.293, 257.2923, 257.293, 257.293, 257.2936, 257.2934, 257.295, 
    257.2942, 257.2966, 257.2975, 257.3001, 257.3017, 257.3034, 257.3041, 
    257.3044, 257.3044,
  259.794, 259.7949, 259.7947, 259.7954, 259.795, 259.7954, 259.7942, 
    259.7949, 259.7945, 259.7941, 259.7967, 259.7954, 259.798, 259.7972, 
    259.7993, 259.7979, 259.7996, 259.7993, 259.8003, 259.8, 259.8012, 
    259.8004, 259.8019, 259.8011, 259.8012, 259.8004, 259.7957, 259.7965, 
    259.7956, 259.7957, 259.7957, 259.795, 259.7947, 259.794, 259.7941, 
    259.7946, 259.7958, 259.7954, 259.7964, 259.7964, 259.7975, 259.797, 
    259.799, 259.7984, 259.8, 259.7996, 259.8, 259.7999, 259.8, 259.7994, 
    259.7997, 259.7991, 259.7971, 259.7977, 259.796, 259.7949, 259.7943, 
    259.7938, 259.7939, 259.794, 259.7946, 259.7953, 259.7957, 259.7961, 
    259.7964, 259.7973, 259.7979, 259.799, 259.7989, 259.7992, 259.7996, 
    259.8001, 259.8, 259.8003, 259.7992, 259.7999, 259.7987, 259.799, 
    259.7964, 259.7955, 259.7951, 259.7947, 259.7939, 259.7945, 259.7943, 
    259.7948, 259.7952, 259.795, 259.7961, 259.7957, 259.7979, 259.7969, 
    259.7995, 259.7989, 259.7997, 259.7993, 259.8, 259.7993, 259.8004, 
    259.8006, 259.8005, 259.8011, 259.7993, 259.8, 259.795, 259.795, 
    259.7951, 259.7946, 259.7945, 259.794, 259.7945, 259.7947, 259.7952, 
    259.7955, 259.7958, 259.7964, 259.7971, 259.7982, 259.7989, 259.7994, 
    259.7991, 259.7994, 259.7991, 259.799, 259.8005, 259.7997, 259.801, 
    259.8009, 259.8003, 259.8009, 259.795, 259.7949, 259.7943, 259.7947, 
    259.7939, 259.7944, 259.7946, 259.7957, 259.7959, 259.7961, 259.7965, 
    259.797, 259.798, 259.7988, 259.7996, 259.7995, 259.7995, 259.7997, 
    259.7993, 259.7998, 259.7999, 259.7997, 259.8009, 259.8006, 259.8009, 
    259.8007, 259.7949, 259.7952, 259.795, 259.7953, 259.7951, 259.796, 
    259.7963, 259.7975, 259.797, 259.7979, 259.7971, 259.7972, 259.7979, 
    259.7971, 259.7987, 259.7976, 259.7997, 259.7986, 259.7998, 259.7996, 
    259.7999, 259.8003, 259.8007, 259.8014, 259.8012, 259.8018, 259.7956, 
    259.796, 259.796, 259.7963, 259.7966, 259.7972, 259.7982, 259.7979, 
    259.7985, 259.7987, 259.7976, 259.7982, 259.7962, 259.7965, 259.7964, 
    259.7956, 259.7979, 259.7967, 259.799, 259.7983, 259.8002, 259.7992, 
    259.8011, 259.8019, 259.8027, 259.8036, 259.7962, 259.7959, 259.7964, 
    259.797, 259.7975, 259.7983, 259.7984, 259.7986, 259.799, 259.7993, 
    259.7986, 259.7993, 259.7966, 259.798, 259.7958, 259.7965, 259.7969, 
    259.7968, 259.7978, 259.7981, 259.7991, 259.7986, 259.8017, 259.8003, 
    259.8044, 259.8032, 259.7958, 259.7962, 259.7973, 259.7968, 259.7984, 
    259.7988, 259.7991, 259.7995, 259.7996, 259.7998, 259.7994, 259.7998, 
    259.7983, 259.799, 259.7972, 259.7976, 259.7975, 259.7972, 259.7979, 
    259.7986, 259.7986, 259.7989, 259.7995, 259.7984, 259.8019, 259.7997, 
    259.7965, 259.7972, 259.7973, 259.797, 259.7987, 259.7981, 259.7998, 
    259.7993, 259.8001, 259.7997, 259.7997, 259.7992, 259.7989, 259.7981, 
    259.7975, 259.7971, 259.7972, 259.7977, 259.7986, 259.7996, 259.7994, 
    259.8, 259.7983, 259.799, 259.7987, 259.7995, 259.7978, 259.7992, 
    259.7975, 259.7976, 259.7981, 259.799, 259.7993, 259.7995, 259.7994, 
    259.7987, 259.7986, 259.7981, 259.7979, 259.7976, 259.7973, 259.7976, 
    259.7979, 259.7987, 259.7994, 259.8003, 259.8004, 259.8014, 259.8006, 
    259.8019, 259.8008, 259.8027, 259.7993, 259.8008, 259.7981, 259.7984, 
    259.7989, 259.8001, 259.7995, 259.8002, 259.7986, 259.7977, 259.7975, 
    259.7971, 259.7975, 259.7975, 259.7979, 259.7978, 259.7987, 259.7982, 
    259.7997, 259.8002, 259.8018, 259.8028, 259.8038, 259.8042, 259.8044, 
    259.8044,
  262.0097, 262.0099, 262.0099, 262.0101, 262.01, 262.0101, 262.0098, 
    262.0099, 262.0099, 262.0098, 262.0104, 262.0101, 262.0108, 262.0106, 
    262.0111, 262.0107, 262.0112, 262.0111, 262.0114, 262.0114, 262.0117, 
    262.0115, 262.0119, 262.0117, 262.0117, 262.0114, 262.0102, 262.0104, 
    262.0101, 262.0102, 262.0102, 262.01, 262.0099, 262.0097, 262.0098, 
    262.0099, 262.0102, 262.0101, 262.0103, 262.0103, 262.0107, 262.0105, 
    262.011, 262.0109, 262.0114, 262.0112, 262.0114, 262.0113, 262.0114, 
    262.0112, 262.0112, 262.0111, 262.0105, 262.0107, 262.0102, 262.0099, 
    262.0098, 262.0097, 262.0097, 262.0097, 262.0099, 262.01, 262.0102, 
    262.0103, 262.0103, 262.0106, 262.0107, 262.0111, 262.011, 262.0111, 
    262.0112, 262.0114, 262.0114, 262.0114, 262.0111, 262.0113, 262.011, 
    262.0111, 262.0103, 262.0101, 262.01, 262.0099, 262.0097, 262.0099, 
    262.0098, 262.0099, 262.01, 262.01, 262.0103, 262.0102, 262.0107, 
    262.0105, 262.0112, 262.011, 262.0113, 262.0111, 262.0113, 262.0112, 
    262.0114, 262.0115, 262.0115, 262.0117, 262.0111, 262.0113, 262.01, 
    262.01, 262.01, 262.0099, 262.0099, 262.0097, 262.0099, 262.0099, 262.01, 
    262.0101, 262.0102, 262.0103, 262.0106, 262.0108, 262.011, 262.0112, 
    262.0111, 262.0112, 262.0111, 262.011, 262.0115, 262.0112, 262.0116, 
    262.0116, 262.0114, 262.0116, 262.01, 262.0099, 262.0098, 262.0099, 
    262.0097, 262.0098, 262.0099, 262.0102, 262.0102, 262.0103, 262.0104, 
    262.0105, 262.0108, 262.011, 262.0112, 262.0112, 262.0112, 262.0113, 
    262.0111, 262.0113, 262.0113, 262.0112, 262.0116, 262.0115, 262.0116, 
    262.0115, 262.0099, 262.01, 262.01, 262.0101, 262.01, 262.0103, 262.0103, 
    262.0107, 262.0105, 262.0107, 262.0105, 262.0106, 262.0107, 262.0106, 
    262.011, 262.0107, 262.0113, 262.011, 262.0113, 262.0112, 262.0113, 
    262.0114, 262.0115, 262.0117, 262.0117, 262.0119, 262.0101, 262.0102, 
    262.0102, 262.0103, 262.0104, 262.0106, 262.0108, 262.0107, 262.0109, 
    262.011, 262.0107, 262.0109, 262.0103, 262.0104, 262.0103, 262.0102, 
    262.0108, 262.0104, 262.011, 262.0109, 262.0114, 262.0111, 262.0117, 
    262.0119, 262.0121, 262.0124, 262.0103, 262.0102, 262.0103, 262.0105, 
    262.0107, 262.0109, 262.0109, 262.0109, 262.011, 262.0111, 262.011, 
    262.0112, 262.0104, 262.0108, 262.0102, 262.0104, 262.0105, 262.0104, 
    262.0107, 262.0108, 262.0111, 262.0109, 262.0118, 262.0114, 262.0126, 
    262.0123, 262.0102, 262.0103, 262.0106, 262.0104, 262.0109, 262.011, 
    262.0111, 262.0112, 262.0112, 262.0113, 262.0112, 262.0113, 262.0109, 
    262.011, 262.0106, 262.0107, 262.0106, 262.0106, 262.0107, 262.011, 
    262.011, 262.011, 262.0112, 262.0109, 262.0119, 262.0113, 262.0104, 
    262.0106, 262.0106, 262.0105, 262.011, 262.0108, 262.0113, 262.0112, 
    262.0114, 262.0113, 262.0113, 262.0111, 262.011, 262.0108, 262.0107, 
    262.0105, 262.0106, 262.0107, 262.011, 262.0112, 262.0112, 262.0114, 
    262.0109, 262.011, 262.011, 262.0112, 262.0107, 262.0111, 262.0107, 
    262.0107, 262.0108, 262.0111, 262.0111, 262.0112, 262.0112, 262.011, 
    262.0109, 262.0108, 262.0108, 262.0107, 262.0106, 262.0107, 262.0107, 
    262.011, 262.0112, 262.0114, 262.0115, 262.0117, 262.0115, 262.0119, 
    262.0116, 262.0121, 262.0111, 262.0116, 262.0108, 262.0109, 262.011, 
    262.0114, 262.0112, 262.0114, 262.0109, 262.0107, 262.0107, 262.0105, 
    262.0107, 262.0107, 262.0107, 262.0107, 262.011, 262.0108, 262.0113, 
    262.0114, 262.0119, 262.0121, 262.0125, 262.0126, 262.0126, 262.0127,
  262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985,
  263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1113, 263.1236, 263.1212, 263.1312, 263.1257, 263.1322, 263.1138, 
    263.1241, 263.1176, 263.1124, 263.1503, 263.1316, 263.1697, 263.1578, 
    263.1877, 263.1678, 263.1916, 263.1871, 263.2007, 263.1968, 263.214, 
    263.2025, 263.223, 263.2113, 263.2131, 263.2021, 263.1354, 263.1479, 
    263.1347, 263.1365, 263.1357, 263.1258, 263.1208, 263.1104, 263.1123, 
    263.1199, 263.1373, 263.1314, 263.1462, 263.1459, 263.1622, 263.1548, 
    263.1823, 263.1746, 263.197, 263.1914, 263.1967, 263.1951, 263.1967, 
    263.1885, 263.192, 263.1848, 263.1562, 263.1646, 263.1396, 263.1243, 
    263.1143, 263.1071, 263.1081, 263.11, 263.12, 263.1293, 263.1364, 
    263.1412, 263.1458, 263.1598, 263.1673, 263.1839, 263.1809, 263.186, 
    263.1908, 263.1988, 263.1975, 263.201, 263.1859, 263.196, 263.1792, 
    263.1838, 263.147, 263.133, 263.1269, 263.1217, 263.1089, 263.1177, 
    263.1143, 263.1226, 263.1278, 263.1252, 263.1413, 263.135, 263.1677, 
    263.1537, 263.1902, 263.1815, 263.1923, 263.1868, 263.1962, 263.1878, 
    263.2024, 263.2055, 263.2034, 263.2117, 263.1873, 263.1967, 263.1252, 
    263.1256, 263.1276, 263.1188, 263.1183, 263.1103, 263.1174, 263.1205, 
    263.1281, 263.1327, 263.137, 263.1464, 263.1569, 263.1716, 263.1821, 
    263.1891, 263.1848, 263.1886, 263.1844, 263.1824, 263.2043, 263.192, 
    263.2105, 263.2095, 263.2011, 263.2096, 263.1259, 263.1234, 263.1149, 
    263.1216, 263.1095, 263.1162, 263.1201, 263.1352, 263.1385, 263.1415, 
    263.1475, 263.1552, 263.1687, 263.1804, 263.1911, 263.1903, 263.1906, 
    263.1929, 263.1871, 263.1939, 263.195, 263.1921, 263.2093, 263.2044, 
    263.2094, 263.2062, 263.1242, 263.1284, 263.1261, 263.1303, 263.1273, 
    263.1404, 263.1443, 263.1625, 263.1551, 263.167, 263.1563, 263.1582, 
    263.1673, 263.1569, 263.1798, 263.1642, 263.193, 263.1776, 263.194, 
    263.191, 263.1959, 263.2003, 263.2058, 263.2159, 263.2136, 263.222, 
    263.1345, 263.1398, 263.1393, 263.1449, 263.149, 263.1579, 263.1721, 
    263.1667, 263.1765, 263.1785, 263.1636, 263.1728, 263.1433, 263.1481, 
    263.1453, 263.1349, 263.1679, 263.151, 263.1823, 263.1731, 263.1997, 
    263.1865, 263.2122, 263.2232, 263.2335, 263.2455, 263.1427, 263.1391, 
    263.1455, 263.1544, 263.1627, 263.1737, 263.1748, 263.1768, 263.1822, 
    263.1866, 263.1775, 263.1877, 263.1491, 263.1694, 263.1377, 263.1472, 
    263.1539, 263.151, 263.1661, 263.1697, 263.1841, 263.1767, 263.2205, 
    263.2012, 263.2547, 263.2397, 263.1378, 263.1427, 263.1595, 263.1515, 
    263.1744, 263.1801, 263.1846, 263.1904, 263.191, 263.1945, 263.1889, 
    263.1942, 263.1737, 263.1829, 263.1576, 263.1638, 263.1609, 263.1578, 
    263.1674, 263.1776, 263.1779, 263.1811, 263.1902, 263.1745, 263.2229, 
    263.1931, 263.148, 263.1573, 263.1586, 263.155, 263.1795, 263.1706, 
    263.1944, 263.188, 263.1984, 263.1933, 263.1925, 263.1858, 263.1816, 
    263.171, 263.1624, 263.1555, 263.1571, 263.1646, 263.1783, 263.1911, 
    263.1883, 263.1976, 263.1728, 263.1832, 263.1792, 263.1897, 263.1666, 
    263.1862, 263.1616, 263.1637, 263.1704, 263.1839, 263.187, 263.1901, 
    263.1882, 263.1786, 263.1771, 263.1703, 263.1684, 263.1632, 263.159, 
    263.1629, 263.167, 263.1786, 263.1891, 263.2003, 263.2031, 263.2162, 
    263.2055, 263.2231, 263.2081, 263.234, 263.1874, 263.2077, 263.1708, 
    263.1748, 263.182, 263.1985, 263.1897, 263.2, 263.177, 263.1649, 
    263.1618, 263.1559, 263.1619, 263.1614, 263.1672, 263.1653, 263.179, 
    263.1717, 263.1925, 263.2, 263.2211, 263.234, 263.2472, 263.253, 
    263.2548, 263.2555 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9096, 253.9104, 253.9103, 253.911, 253.9106, 253.911, 253.9098, 
    253.9105, 253.91, 253.9097, 253.9123, 253.911, 253.9136, 253.9128, 
    253.9149, 253.9135, 253.9152, 253.9149, 253.9158, 253.9155, 253.9167, 
    253.9159, 253.9174, 253.9165, 253.9167, 253.9159, 253.9113, 253.9121, 
    253.9112, 253.9113, 253.9113, 253.9106, 253.9102, 253.9095, 253.9097, 
    253.9102, 253.9114, 253.911, 253.912, 253.912, 253.9131, 253.9126, 
    253.9145, 253.914, 253.9155, 253.9151, 253.9155, 253.9154, 253.9155, 
    253.9149, 253.9152, 253.9147, 253.9127, 253.9133, 253.9115, 253.9105, 
    253.9098, 253.9093, 253.9094, 253.9095, 253.9102, 253.9108, 253.9113, 
    253.9117, 253.912, 253.9129, 253.9135, 253.9146, 253.9144, 253.9148, 
    253.9151, 253.9157, 253.9156, 253.9158, 253.9148, 253.9155, 253.9143, 
    253.9146, 253.912, 253.9111, 253.9107, 253.9103, 253.9094, 253.91, 
    253.9098, 253.9104, 253.9107, 253.9106, 253.9117, 253.9112, 253.9135, 
    253.9125, 253.9151, 253.9145, 253.9152, 253.9148, 253.9155, 253.9149, 
    253.9159, 253.9161, 253.916, 253.9166, 253.9149, 253.9155, 253.9106, 
    253.9106, 253.9107, 253.9101, 253.9101, 253.9095, 253.91, 253.9102, 
    253.9108, 253.9111, 253.9114, 253.912, 253.9128, 253.9138, 253.9145, 
    253.915, 253.9147, 253.915, 253.9147, 253.9145, 253.9161, 253.9152, 
    253.9165, 253.9164, 253.9158, 253.9164, 253.9106, 253.9104, 253.9098, 
    253.9103, 253.9095, 253.9099, 253.9102, 253.9112, 253.9115, 253.9117, 
    253.9121, 253.9126, 253.9136, 253.9144, 253.9151, 253.9151, 253.9151, 
    253.9153, 253.9149, 253.9153, 253.9154, 253.9152, 253.9164, 253.9161, 
    253.9164, 253.9162, 253.9105, 253.9108, 253.9106, 253.9109, 253.9107, 
    253.9116, 253.9119, 253.9131, 253.9126, 253.9135, 253.9127, 253.9128, 
    253.9135, 253.9128, 253.9143, 253.9133, 253.9153, 253.9142, 253.9153, 
    253.9151, 253.9155, 253.9158, 253.9162, 253.9169, 253.9167, 253.9173, 
    253.9112, 253.9116, 253.9115, 253.9119, 253.9122, 253.9128, 253.9138, 
    253.9135, 253.9141, 253.9143, 253.9132, 253.9138, 253.9118, 253.9121, 
    253.912, 253.9112, 253.9135, 253.9123, 253.9145, 253.9139, 253.9157, 
    253.9148, 253.9166, 253.9174, 253.9181, 253.919, 253.9118, 253.9115, 
    253.912, 253.9126, 253.9132, 253.9139, 253.914, 253.9141, 253.9145, 
    253.9148, 253.9142, 253.9149, 253.9122, 253.9136, 253.9114, 253.9121, 
    253.9126, 253.9124, 253.9134, 253.9137, 253.9146, 253.9141, 253.9172, 
    253.9158, 253.9196, 253.9185, 253.9114, 253.9118, 253.9129, 253.9124, 
    253.914, 253.9144, 253.9147, 253.9151, 253.9151, 253.9154, 253.915, 
    253.9154, 253.9139, 253.9146, 253.9128, 253.9132, 253.913, 253.9128, 
    253.9135, 253.9142, 253.9142, 253.9144, 253.915, 253.914, 253.9173, 
    253.9152, 253.9121, 253.9128, 253.9129, 253.9126, 253.9143, 253.9137, 
    253.9154, 253.9149, 253.9156, 253.9153, 253.9152, 253.9148, 253.9145, 
    253.9137, 253.9131, 253.9127, 253.9128, 253.9133, 253.9142, 253.9151, 
    253.9149, 253.9156, 253.9139, 253.9146, 253.9143, 253.915, 253.9134, 
    253.9147, 253.9131, 253.9132, 253.9137, 253.9146, 253.9148, 253.9151, 
    253.9149, 253.9143, 253.9142, 253.9137, 253.9136, 253.9132, 253.9129, 
    253.9132, 253.9135, 253.9143, 253.915, 253.9158, 253.916, 253.9169, 
    253.9161, 253.9173, 253.9163, 253.9181, 253.9149, 253.9163, 253.9137, 
    253.914, 253.9145, 253.9156, 253.915, 253.9158, 253.9142, 253.9133, 
    253.9131, 253.9127, 253.9131, 253.9131, 253.9135, 253.9133, 253.9143, 
    253.9138, 253.9152, 253.9157, 253.9172, 253.9182, 253.9191, 253.9195, 
    253.9196, 253.9197 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1456413, 0.1456405, 0.1456406, 0.1456399, 0.1456403, 0.1456399, 
    0.1456411, 0.1456404, 0.1456409, 0.1456413, 0.1456387, 0.1456399, 
    0.1456375, 0.1456382, 0.1456364, 0.1456376, 0.1456362, 0.1456365, 
    0.1456357, 0.1456359, 0.1456351, 0.1456356, 0.1456347, 0.1456352, 
    0.1456351, 0.1456356, 0.1456397, 0.1456388, 0.1456397, 0.1456396, 
    0.1456396, 0.1456403, 0.1456407, 0.1456414, 0.1456413, 0.1456407, 
    0.1456395, 0.1456399, 0.145639, 0.145639, 0.1456379, 0.1456384, 
    0.1456367, 0.1456372, 0.1456359, 0.1456362, 0.1456359, 0.145636, 
    0.1456359, 0.1456364, 0.1456362, 0.1456366, 0.1456383, 0.1456378, 
    0.1456394, 0.1456404, 0.1456411, 0.1456416, 0.1456416, 0.1456414, 
    0.1456407, 0.1456401, 0.1456396, 0.1456393, 0.145639, 0.1456381, 
    0.1456376, 0.1456366, 0.1456368, 0.1456365, 0.1456362, 0.1456358, 
    0.1456359, 0.1456357, 0.1456365, 0.145636, 0.1456369, 0.1456366, 
    0.1456389, 0.1456398, 0.1456402, 0.1456406, 0.1456415, 0.1456409, 
    0.1456411, 0.1456405, 0.1456402, 0.1456403, 0.1456393, 0.1456397, 
    0.1456376, 0.1456385, 0.1456363, 0.1456368, 0.1456362, 0.1456365, 
    0.145636, 0.1456364, 0.1456356, 0.1456355, 0.1456356, 0.1456352, 
    0.1456364, 0.1456359, 0.1456404, 0.1456403, 0.1456402, 0.1456408, 
    0.1456408, 0.1456414, 0.1456409, 0.1456407, 0.1456401, 0.1456398, 
    0.1456396, 0.1456389, 0.1456383, 0.1456374, 0.1456367, 0.1456363, 
    0.1456366, 0.1456364, 0.1456366, 0.1456367, 0.1456355, 0.1456362, 
    0.1456352, 0.1456353, 0.1456357, 0.1456353, 0.1456403, 0.1456405, 
    0.1456411, 0.1456406, 0.1456415, 0.145641, 0.1456407, 0.1456397, 
    0.1456394, 0.1456393, 0.1456389, 0.1456384, 0.1456375, 0.1456368, 
    0.1456362, 0.1456363, 0.1456363, 0.1456361, 0.1456365, 0.1456361, 
    0.145636, 0.1456362, 0.1456353, 0.1456355, 0.1456353, 0.1456354, 
    0.1456404, 0.1456401, 0.1456403, 0.14564, 0.1456402, 0.1456393, 
    0.1456391, 0.1456379, 0.1456384, 0.1456376, 0.1456383, 0.1456382, 
    0.1456376, 0.1456383, 0.1456369, 0.1456378, 0.1456361, 0.145637, 
    0.1456361, 0.1456362, 0.145636, 0.1456357, 0.1456355, 0.145635, 
    0.1456351, 0.1456347, 0.1456397, 0.1456394, 0.1456394, 0.145639, 
    0.1456388, 0.1456382, 0.1456373, 0.1456377, 0.1456371, 0.145637, 
    0.1456379, 0.1456373, 0.1456391, 0.1456388, 0.145639, 0.1456397, 
    0.1456376, 0.1456386, 0.1456367, 0.1456373, 0.1456358, 0.1456365, 
    0.1456351, 0.1456346, 0.1456342, 0.1456337, 0.1456392, 0.1456394, 
    0.145639, 0.1456384, 0.1456379, 0.1456372, 0.1456372, 0.1456371, 
    0.1456367, 0.1456365, 0.145637, 0.1456364, 0.1456388, 0.1456375, 
    0.1456395, 0.1456389, 0.1456385, 0.1456386, 0.1456377, 0.1456375, 
    0.1456366, 0.1456371, 0.1456348, 0.1456357, 0.1456334, 0.1456339, 
    0.1456395, 0.1456392, 0.1456381, 0.1456386, 0.1456372, 0.1456369, 
    0.1456366, 0.1456363, 0.1456362, 0.1456361, 0.1456363, 0.1456361, 
    0.1456372, 0.1456367, 0.1456382, 0.1456378, 0.145638, 0.1456382, 
    0.1456376, 0.145637, 0.145637, 0.1456368, 0.1456363, 0.1456372, 
    0.1456347, 0.1456361, 0.1456388, 0.1456382, 0.1456382, 0.1456384, 
    0.1456369, 0.1456374, 0.1456361, 0.1456364, 0.1456358, 0.1456361, 
    0.1456362, 0.1456365, 0.1456368, 0.1456374, 0.1456379, 0.1456383, 
    0.1456383, 0.1456378, 0.145637, 0.1456362, 0.1456364, 0.1456359, 
    0.1456373, 0.1456367, 0.1456369, 0.1456363, 0.1456377, 0.1456365, 
    0.145638, 0.1456378, 0.1456374, 0.1456366, 0.1456365, 0.1456363, 
    0.1456364, 0.145637, 0.1456371, 0.1456375, 0.1456376, 0.1456379, 
    0.1456381, 0.1456379, 0.1456376, 0.145637, 0.1456363, 0.1456357, 
    0.1456356, 0.145635, 0.1456355, 0.1456346, 0.1456353, 0.1456342, 
    0.1456364, 0.1456354, 0.1456374, 0.1456372, 0.1456367, 0.1456358, 
    0.1456363, 0.1456358, 0.1456371, 0.1456378, 0.145638, 0.1456383, 
    0.145638, 0.145638, 0.1456376, 0.1456378, 0.1456369, 0.1456374, 
    0.1456362, 0.1456358, 0.1456347, 0.1456342, 0.1456337, 0.1456334, 
    0.1456334, 0.1456334,
  0.1512737, 0.1512784, 0.1512775, 0.1512813, 0.1512792, 0.1512817, 
    0.1512747, 0.1512786, 0.1512761, 0.1512742, 0.1512886, 0.1512815, 
    0.1512963, 0.1512917, 0.1513034, 0.1512955, 0.151305, 0.1513032, 
    0.1513087, 0.1513071, 0.151314, 0.1513094, 0.1513178, 0.151313, 
    0.1513137, 0.1513093, 0.151283, 0.1512877, 0.1512827, 0.1512834, 
    0.1512831, 0.1512793, 0.1512773, 0.1512734, 0.1512741, 0.151277, 
    0.1512837, 0.1512814, 0.1512872, 0.1512871, 0.1512934, 0.1512906, 
    0.1513013, 0.1512983, 0.1513072, 0.1513049, 0.1513071, 0.1513065, 
    0.1513071, 0.1513038, 0.1513052, 0.1513023, 0.1512911, 0.1512944, 
    0.1512846, 0.1512786, 0.1512749, 0.1512721, 0.1512725, 0.1512732, 
    0.151277, 0.1512807, 0.1512834, 0.1512852, 0.151287, 0.1512924, 
    0.1512953, 0.1513019, 0.1513008, 0.1513027, 0.1513047, 0.151308, 
    0.1513074, 0.1513088, 0.1513027, 0.1513068, 0.1513001, 0.1513019, 
    0.1512873, 0.1512821, 0.1512796, 0.1512777, 0.1512728, 0.1512762, 
    0.1512748, 0.1512781, 0.1512801, 0.1512791, 0.1512853, 0.1512829, 
    0.1512955, 0.1512901, 0.1513045, 0.151301, 0.1513053, 0.1513031, 
    0.1513069, 0.1513035, 0.1513094, 0.1513106, 0.1513098, 0.1513132, 
    0.1513033, 0.1513071, 0.151279, 0.1512792, 0.15128, 0.1512766, 0.1512764, 
    0.1512734, 0.1512761, 0.1512772, 0.1512802, 0.1512819, 0.1512836, 
    0.1512873, 0.1512913, 0.1512971, 0.1513012, 0.1513041, 0.1513023, 
    0.1513039, 0.1513022, 0.1513014, 0.1513101, 0.1513052, 0.1513127, 
    0.1513123, 0.1513089, 0.1513123, 0.1512793, 0.1512784, 0.1512751, 
    0.1512777, 0.151273, 0.1512756, 0.1512771, 0.1512828, 0.1512842, 
    0.1512854, 0.1512877, 0.1512907, 0.1512959, 0.1513005, 0.1513048, 
    0.1513045, 0.1513046, 0.1513056, 0.1513032, 0.151306, 0.1513064, 
    0.1513052, 0.1513122, 0.1513102, 0.1513123, 0.151311, 0.1512787, 
    0.1512803, 0.1512794, 0.151281, 0.1512799, 0.1512849, 0.1512864, 
    0.1512935, 0.1512906, 0.1512952, 0.1512911, 0.1512918, 0.1512953, 
    0.1512914, 0.1513003, 0.1512941, 0.1513056, 0.1512993, 0.151306, 
    0.1513048, 0.1513068, 0.1513085, 0.1513108, 0.1513149, 0.1513139, 
    0.1513174, 0.1512826, 0.1512846, 0.1512845, 0.1512867, 0.1512883, 
    0.1512917, 0.1512973, 0.1512952, 0.1512991, 0.1512998, 0.151294, 
    0.1512975, 0.151286, 0.1512878, 0.1512868, 0.1512828, 0.1512956, 
    0.151289, 0.1513013, 0.1512977, 0.1513083, 0.1513029, 0.1513134, 
    0.1513178, 0.1513222, 0.151327, 0.1512858, 0.1512844, 0.1512869, 
    0.1512903, 0.1512936, 0.1512979, 0.1512984, 0.1512992, 0.1513013, 
    0.1513031, 0.1512994, 0.1513035, 0.1512882, 0.1512962, 0.1512839, 
    0.1512875, 0.1512901, 0.151289, 0.151295, 0.1512964, 0.151302, 0.1512991, 
    0.1513166, 0.1513088, 0.1513309, 0.1513247, 0.1512839, 0.1512858, 
    0.1512923, 0.1512893, 0.1512982, 0.1513004, 0.1513023, 0.1513045, 
    0.1513048, 0.1513062, 0.1513039, 0.1513061, 0.1512979, 0.1513016, 
    0.1512917, 0.151294, 0.1512929, 0.1512917, 0.1512955, 0.1512994, 
    0.1512996, 0.1513008, 0.1513042, 0.1512983, 0.1513175, 0.1513054, 
    0.1512879, 0.1512914, 0.151292, 0.1512906, 0.1513002, 0.1512967, 
    0.1513062, 0.1513036, 0.1513078, 0.1513057, 0.1513054, 0.1513027, 
    0.1513011, 0.1512969, 0.1512935, 0.1512908, 0.1512915, 0.1512944, 
    0.1512997, 0.1513048, 0.1513037, 0.1513075, 0.1512976, 0.1513017, 
    0.1513001, 0.1513043, 0.1512951, 0.1513027, 0.1512932, 0.151294, 
    0.1512967, 0.1513019, 0.1513032, 0.1513044, 0.1513037, 0.1512998, 
    0.1512993, 0.1512966, 0.1512958, 0.1512939, 0.1512922, 0.1512937, 
    0.1512953, 0.1512999, 0.151304, 0.1513086, 0.1513097, 0.1513149, 
    0.1513105, 0.1513176, 0.1513114, 0.1513222, 0.1513032, 0.1513114, 
    0.1512968, 0.1512984, 0.1513011, 0.1513077, 0.1513043, 0.1513084, 
    0.1512992, 0.1512944, 0.1512933, 0.151291, 0.1512933, 0.1512931, 
    0.1512954, 0.1512947, 0.1513, 0.1512972, 0.1513054, 0.1513084, 0.151317, 
    0.1513223, 0.1513278, 0.1513303, 0.151331, 0.1513313,
  0.1611244, 0.1611304, 0.1611293, 0.1611341, 0.1611315, 0.1611346, 
    0.1611257, 0.1611306, 0.1611275, 0.161125, 0.1611434, 0.1611343, 
    0.1611533, 0.1611474, 0.1611624, 0.1611523, 0.1611645, 0.1611622, 
    0.1611693, 0.1611672, 0.1611761, 0.1611702, 0.1611809, 0.1611748, 
    0.1611757, 0.16117, 0.1611363, 0.1611422, 0.1611359, 0.1611367, 
    0.1611364, 0.1611315, 0.161129, 0.161124, 0.1611249, 0.1611286, 
    0.1611371, 0.1611343, 0.1611416, 0.1611415, 0.1611496, 0.1611459, 
    0.1611598, 0.1611558, 0.1611673, 0.1611644, 0.1611672, 0.1611664, 
    0.1611672, 0.1611629, 0.1611647, 0.161161, 0.1611466, 0.1611508, 
    0.1611383, 0.1611307, 0.1611259, 0.1611224, 0.1611229, 0.1611238, 
    0.1611286, 0.1611333, 0.1611368, 0.1611391, 0.1611414, 0.1611482, 
    0.1611521, 0.1611605, 0.1611591, 0.1611616, 0.1611641, 0.1611683, 
    0.1611676, 0.1611694, 0.1611616, 0.1611668, 0.1611582, 0.1611605, 
    0.1611417, 0.1611351, 0.161132, 0.1611295, 0.1611233, 0.1611276, 
    0.1611259, 0.16113, 0.1611325, 0.1611313, 0.1611392, 0.1611361, 
    0.1611523, 0.1611453, 0.1611638, 0.1611594, 0.1611649, 0.1611621, 
    0.1611669, 0.1611626, 0.1611701, 0.1611717, 0.1611706, 0.161175, 
    0.1611623, 0.1611671, 0.1611312, 0.1611314, 0.1611324, 0.1611281, 
    0.1611278, 0.161124, 0.1611274, 0.1611289, 0.1611327, 0.1611349, 
    0.161137, 0.1611417, 0.1611469, 0.1611543, 0.1611597, 0.1611633, 
    0.1611611, 0.161163, 0.1611608, 0.1611598, 0.1611711, 0.1611647, 
    0.1611744, 0.1611739, 0.1611695, 0.1611739, 0.1611316, 0.1611304, 
    0.1611262, 0.1611295, 0.1611236, 0.1611268, 0.1611287, 0.1611361, 
    0.1611378, 0.1611393, 0.1611423, 0.1611461, 0.1611528, 0.1611588, 
    0.1611643, 0.1611639, 0.161164, 0.1611652, 0.1611622, 0.1611657, 
    0.1611663, 0.1611648, 0.1611738, 0.1611712, 0.1611739, 0.1611722, 
    0.1611308, 0.1611328, 0.1611317, 0.1611337, 0.1611323, 0.1611387, 
    0.1611406, 0.1611497, 0.161146, 0.1611519, 0.1611467, 0.1611476, 
    0.161152, 0.161147, 0.1611584, 0.1611505, 0.1611653, 0.1611572, 
    0.1611658, 0.1611643, 0.1611668, 0.161169, 0.1611719, 0.1611772, 
    0.161176, 0.1611805, 0.1611358, 0.1611384, 0.1611382, 0.161141, 0.161143, 
    0.1611474, 0.1611546, 0.1611519, 0.1611569, 0.1611578, 0.1611503, 
    0.1611549, 0.1611402, 0.1611425, 0.1611411, 0.161136, 0.1611524, 
    0.1611439, 0.1611597, 0.1611551, 0.1611687, 0.1611619, 0.1611753, 
    0.1611809, 0.1611866, 0.1611929, 0.1611399, 0.1611381, 0.1611413, 
    0.1611456, 0.1611499, 0.1611554, 0.161156, 0.161157, 0.1611597, 0.161162, 
    0.1611573, 0.1611626, 0.1611429, 0.1611532, 0.1611374, 0.161142, 
    0.1611454, 0.161144, 0.1611516, 0.1611534, 0.1611606, 0.1611569, 
    0.1611795, 0.1611694, 0.1611979, 0.1611898, 0.1611375, 0.1611399, 
    0.1611482, 0.1611443, 0.1611558, 0.1611586, 0.161161, 0.1611639, 
    0.1611643, 0.161166, 0.1611631, 0.1611659, 0.1611554, 0.1611601, 
    0.1611473, 0.1611504, 0.161149, 0.1611474, 0.1611523, 0.1611573, 
    0.1611575, 0.1611591, 0.1611635, 0.1611558, 0.1611806, 0.161165, 
    0.1611425, 0.161147, 0.1611478, 0.161146, 0.1611583, 0.1611538, 0.161166, 
    0.1611627, 0.1611681, 0.1611654, 0.161165, 0.1611616, 0.1611594, 
    0.161154, 0.1611497, 0.1611463, 0.1611471, 0.1611508, 0.1611577, 
    0.1611642, 0.1611628, 0.1611677, 0.1611549, 0.1611602, 0.1611581, 
    0.1611636, 0.1611518, 0.1611615, 0.1611493, 0.1611504, 0.1611537, 
    0.1611605, 0.1611621, 0.1611637, 0.1611628, 0.1611578, 0.1611571, 
    0.1611537, 0.1611527, 0.1611502, 0.161148, 0.1611499, 0.161152, 
    0.1611579, 0.1611632, 0.1611691, 0.1611705, 0.1611772, 0.1611716, 
    0.1611807, 0.1611728, 0.1611866, 0.1611622, 0.1611727, 0.1611539, 
    0.161156, 0.1611595, 0.161168, 0.1611635, 0.1611688, 0.1611571, 
    0.1611509, 0.1611494, 0.1611465, 0.1611495, 0.1611492, 0.1611521, 
    0.1611512, 0.1611581, 0.1611544, 0.161165, 0.1611688, 0.1611799, 
    0.1611868, 0.1611939, 0.1611971, 0.161198, 0.1611984,
  0.1753341, 0.1753387, 0.1753378, 0.1753414, 0.1753394, 0.1753418, 
    0.1753351, 0.1753388, 0.1753365, 0.1753346, 0.1753484, 0.1753416, 
    0.175356, 0.1753515, 0.175363, 0.1753552, 0.1753646, 0.1753629, 
    0.1753683, 0.1753668, 0.1753737, 0.1753691, 0.1753774, 0.1753726, 
    0.1753733, 0.1753689, 0.175343, 0.1753476, 0.1753427, 0.1753434, 
    0.1753431, 0.1753394, 0.1753376, 0.1753339, 0.1753345, 0.1753373, 
    0.1753437, 0.1753415, 0.1753471, 0.175347, 0.1753532, 0.1753504, 
    0.175361, 0.175358, 0.1753668, 0.1753646, 0.1753667, 0.1753661, 
    0.1753667, 0.1753634, 0.1753648, 0.1753619, 0.1753509, 0.1753541, 
    0.1753446, 0.1753388, 0.1753352, 0.1753327, 0.175333, 0.1753337, 
    0.1753373, 0.1753408, 0.1753434, 0.1753452, 0.175347, 0.1753521, 
    0.175355, 0.1753615, 0.1753604, 0.1753624, 0.1753643, 0.1753676, 
    0.175367, 0.1753684, 0.1753624, 0.1753664, 0.1753598, 0.1753616, 
    0.1753472, 0.1753421, 0.1753398, 0.1753379, 0.1753333, 0.1753365, 
    0.1753352, 0.1753383, 0.1753402, 0.1753393, 0.1753452, 0.1753429, 
    0.1753552, 0.1753499, 0.1753641, 0.1753607, 0.1753649, 0.1753628, 
    0.1753665, 0.1753631, 0.175369, 0.1753702, 0.1753694, 0.1753728, 
    0.1753629, 0.1753667, 0.1753392, 0.1753394, 0.1753401, 0.1753369, 
    0.1753367, 0.1753338, 0.1753364, 0.1753375, 0.1753404, 0.175342, 
    0.1753436, 0.1753471, 0.1753511, 0.1753567, 0.1753609, 0.1753637, 
    0.175362, 0.1753635, 0.1753618, 0.175361, 0.1753698, 0.1753648, 
    0.1753723, 0.1753719, 0.1753685, 0.1753719, 0.1753395, 0.1753386, 
    0.1753355, 0.1753379, 0.1753335, 0.1753359, 0.1753373, 0.1753429, 
    0.1753442, 0.1753453, 0.1753476, 0.1753505, 0.1753556, 0.1753602, 
    0.1753645, 0.1753642, 0.1753643, 0.1753652, 0.1753629, 0.1753656, 
    0.175366, 0.1753648, 0.1753718, 0.1753698, 0.1753719, 0.1753706, 
    0.1753389, 0.1753404, 0.1753396, 0.1753411, 0.17534, 0.1753448, 
    0.1753463, 0.1753532, 0.1753504, 0.175355, 0.1753509, 0.1753516, 
    0.175355, 0.1753511, 0.1753599, 0.1753539, 0.1753652, 0.175359, 
    0.1753656, 0.1753644, 0.1753664, 0.1753681, 0.1753704, 0.1753745, 
    0.1753736, 0.1753771, 0.1753427, 0.1753446, 0.1753445, 0.1753466, 
    0.1753481, 0.1753515, 0.175357, 0.1753549, 0.1753587, 0.1753595, 
    0.1753537, 0.1753572, 0.175346, 0.1753477, 0.1753467, 0.1753428, 
    0.1753553, 0.1753488, 0.1753609, 0.1753574, 0.1753679, 0.1753626, 
    0.175373, 0.1753774, 0.1753819, 0.1753869, 0.1753457, 0.1753444, 
    0.1753469, 0.1753501, 0.1753534, 0.1753576, 0.1753581, 0.1753588, 
    0.1753609, 0.1753627, 0.175359, 0.1753631, 0.175348, 0.1753559, 
    0.1753439, 0.1753474, 0.17535, 0.1753489, 0.1753547, 0.1753561, 
    0.1753616, 0.1753588, 0.1753763, 0.1753684, 0.1753909, 0.1753844, 
    0.1753439, 0.1753458, 0.1753521, 0.1753491, 0.1753579, 0.1753601, 
    0.1753619, 0.1753642, 0.1753644, 0.1753658, 0.1753636, 0.1753657, 
    0.1753576, 0.1753612, 0.1753514, 0.1753538, 0.1753527, 0.1753515, 
    0.1753552, 0.1753591, 0.1753592, 0.1753605, 0.1753639, 0.1753579, 
    0.1753772, 0.175365, 0.1753478, 0.1753512, 0.1753518, 0.1753504, 
    0.1753599, 0.1753564, 0.1753658, 0.1753632, 0.1753674, 0.1753653, 
    0.175365, 0.1753624, 0.1753607, 0.1753566, 0.1753532, 0.1753507, 
    0.1753512, 0.1753541, 0.1753593, 0.1753644, 0.1753633, 0.1753671, 
    0.1753573, 0.1753613, 0.1753597, 0.1753639, 0.1753549, 0.1753623, 
    0.1753529, 0.1753538, 0.1753563, 0.1753615, 0.1753628, 0.175364, 
    0.1753633, 0.1753595, 0.1753589, 0.1753563, 0.1753555, 0.1753536, 
    0.1753519, 0.1753534, 0.175355, 0.1753595, 0.1753636, 0.1753682, 
    0.1753693, 0.1753745, 0.1753702, 0.1753772, 0.1753711, 0.1753819, 
    0.1753629, 0.175371, 0.1753565, 0.175358, 0.1753608, 0.1753674, 
    0.1753639, 0.175368, 0.1753589, 0.1753542, 0.175353, 0.1753508, 
    0.1753531, 0.1753529, 0.1753551, 0.1753544, 0.1753597, 0.1753568, 
    0.175365, 0.175368, 0.1753767, 0.175382, 0.1753877, 0.1753902, 0.1753909, 
    0.1753913,
  0.1899464, 0.1899478, 0.1899475, 0.1899487, 0.189948, 0.1899488, 0.1899467, 
    0.1899478, 0.1899471, 0.1899466, 0.1899509, 0.1899487, 0.1899534, 
    0.1899519, 0.1899557, 0.1899531, 0.1899563, 0.1899557, 0.1899576, 
    0.189957, 0.1899594, 0.1899578, 0.1899608, 0.189959, 0.1899593, 
    0.1899578, 0.1899492, 0.1899506, 0.1899491, 0.1899493, 0.1899492, 
    0.189948, 0.1899475, 0.1899463, 0.1899465, 0.1899474, 0.1899494, 
    0.1899487, 0.1899505, 0.1899504, 0.1899524, 0.1899515, 0.189955, 
    0.189954, 0.189957, 0.1899562, 0.189957, 0.1899568, 0.189957, 0.1899559, 
    0.1899563, 0.1899554, 0.1899517, 0.1899527, 0.1899496, 0.1899478, 
    0.1899468, 0.189946, 0.1899461, 0.1899463, 0.1899474, 0.1899485, 
    0.1899493, 0.1899499, 0.1899504, 0.1899521, 0.189953, 0.1899552, 
    0.1899548, 0.1899555, 0.1899562, 0.1899573, 0.1899571, 0.1899576, 
    0.1899555, 0.1899569, 0.1899546, 0.1899552, 0.1899505, 0.1899489, 
    0.1899481, 0.1899476, 0.1899462, 0.1899471, 0.1899467, 0.1899477, 
    0.1899483, 0.189948, 0.1899499, 0.1899491, 0.1899531, 0.1899514, 
    0.1899561, 0.1899549, 0.1899564, 0.1899556, 0.1899569, 0.1899558, 
    0.1899578, 0.1899582, 0.1899579, 0.1899591, 0.1899557, 0.189957, 
    0.189948, 0.189948, 0.1899483, 0.1899472, 0.1899472, 0.1899463, 
    0.1899471, 0.1899474, 0.1899483, 0.1899488, 0.1899493, 0.1899505, 
    0.1899517, 0.1899536, 0.189955, 0.1899559, 0.1899554, 0.1899559, 
    0.1899553, 0.1899551, 0.1899581, 0.1899563, 0.1899589, 0.1899588, 
    0.1899576, 0.1899588, 0.1899481, 0.1899478, 0.1899468, 0.1899476, 
    0.1899462, 0.189947, 0.1899474, 0.1899491, 0.1899495, 0.1899499, 
    0.1899506, 0.1899516, 0.1899532, 0.1899548, 0.1899562, 0.1899561, 
    0.1899562, 0.1899565, 0.1899557, 0.1899566, 0.1899568, 0.1899564, 
    0.1899588, 0.1899581, 0.1899588, 0.1899583, 0.1899479, 0.1899484, 
    0.1899481, 0.1899486, 0.1899482, 0.1899497, 0.1899502, 0.1899524, 
    0.1899515, 0.189953, 0.1899517, 0.1899519, 0.189953, 0.1899518, 
    0.1899547, 0.1899526, 0.1899565, 0.1899544, 0.1899566, 0.1899562, 
    0.1899569, 0.1899575, 0.1899583, 0.1899597, 0.1899594, 0.1899606, 
    0.1899491, 0.1899497, 0.1899496, 0.1899503, 0.1899508, 0.1899519, 
    0.1899537, 0.189953, 0.1899543, 0.1899545, 0.1899526, 0.1899538, 
    0.1899501, 0.1899507, 0.1899503, 0.1899491, 0.1899531, 0.189951, 
    0.189955, 0.1899538, 0.1899574, 0.1899556, 0.1899592, 0.1899608, 
    0.1899624, 0.1899642, 0.18995, 0.1899496, 0.1899504, 0.1899514, 
    0.1899525, 0.1899539, 0.189954, 0.1899543, 0.189955, 0.1899556, 
    0.1899544, 0.1899558, 0.1899507, 0.1899533, 0.1899494, 0.1899506, 
    0.1899514, 0.189951, 0.1899529, 0.1899534, 0.1899552, 0.1899543, 
    0.1899604, 0.1899576, 0.1899657, 0.1899633, 0.1899495, 0.18995, 
    0.1899521, 0.1899511, 0.189954, 0.1899547, 0.1899553, 0.1899561, 
    0.1899562, 0.1899567, 0.1899559, 0.1899567, 0.1899539, 0.1899551, 
    0.1899519, 0.1899526, 0.1899523, 0.1899519, 0.1899531, 0.1899544, 
    0.1899544, 0.1899549, 0.189956, 0.189954, 0.1899607, 0.1899564, 
    0.1899507, 0.1899518, 0.189952, 0.1899515, 0.1899547, 0.1899535, 
    0.1899567, 0.1899558, 0.1899572, 0.1899565, 0.1899564, 0.1899555, 
    0.1899549, 0.1899536, 0.1899524, 0.1899516, 0.1899518, 0.1899527, 
    0.1899545, 0.1899562, 0.1899558, 0.1899571, 0.1899538, 0.1899551, 
    0.1899546, 0.189956, 0.189953, 0.1899555, 0.1899524, 0.1899526, 
    0.1899535, 0.1899552, 0.1899557, 0.1899561, 0.1899558, 0.1899545, 
    0.1899543, 0.1899535, 0.1899532, 0.1899526, 0.189952, 0.1899525, 
    0.189953, 0.1899545, 0.1899559, 0.1899575, 0.1899579, 0.1899597, 
    0.1899582, 0.1899607, 0.1899585, 0.1899624, 0.1899557, 0.1899585, 
    0.1899535, 0.189954, 0.189955, 0.1899572, 0.189956, 0.1899574, 0.1899543, 
    0.1899527, 0.1899524, 0.1899517, 0.1899524, 0.1899523, 0.1899531, 
    0.1899528, 0.1899546, 0.1899536, 0.1899564, 0.1899574, 0.1899605, 
    0.1899624, 0.1899645, 0.1899654, 0.1899657, 0.1899658,
  0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.1973189, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.1973191, 0.197319, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.197319, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.197319, 0.197319, 0.197319, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.197319, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 0.197319, 0.197319, 
    0.1973189, 0.197319, 0.1973189, 0.1973189, 0.197319, 0.1973189, 0.197319, 
    0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.197319, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973191, 0.1973191, 0.1973192, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 0.1973193, 
    0.1973192, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.197319, 0.197319, 0.197319, 0.1973191, 
    0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.197319, 0.1973191, 0.1973192, 0.1973193, 
    0.1973193, 0.1973193,
  0.1984799, 0.1984798, 0.1984799, 0.1984798, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 
    0.1984799, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984799, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984798, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984796, 
    0.1984796, 0.1984796,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.611717, 5.61177, 5.61176, 5.611802, 5.611779, 5.611805, 5.611728, 
    5.611771, 5.611744, 5.611722, 5.61188, 5.611804, 5.611965, 5.611915, 
    5.612043, 5.611956, 5.612062, 5.612042, 5.612103, 5.612086, 5.612161, 
    5.612111, 5.612201, 5.612149, 5.612157, 5.612109, 5.61182, 5.61187, 
    5.611817, 5.611824, 5.611821, 5.611779, 5.611757, 5.611714, 5.611722, 
    5.611754, 5.611827, 5.611803, 5.611866, 5.611865, 5.611934, 5.611903, 
    5.61202, 5.611987, 5.612086, 5.612061, 5.612085, 5.612078, 5.612085, 
    5.612048, 5.612064, 5.612031, 5.611908, 5.611944, 5.611837, 5.611771, 
    5.61173, 5.6117, 5.611704, 5.611712, 5.611754, 5.611794, 5.611825, 
    5.611845, 5.611865, 5.611922, 5.611954, 5.612027, 5.612014, 5.612036, 
    5.612059, 5.612094, 5.612089, 5.612104, 5.612036, 5.612081, 5.612007, 
    5.612027, 5.611866, 5.61181, 5.611783, 5.611762, 5.611707, 5.611744, 
    5.61173, 5.611766, 5.611788, 5.611777, 5.611845, 5.611819, 5.611956, 
    5.611897, 5.612056, 5.612017, 5.612065, 5.612041, 5.612082, 5.612045, 
    5.61211, 5.612124, 5.612114, 5.612152, 5.612043, 5.612084, 5.611777, 
    5.611778, 5.611787, 5.611749, 5.611747, 5.611713, 5.611743, 5.611756, 
    5.61179, 5.611808, 5.611827, 5.611867, 5.611911, 5.611973, 5.612019, 
    5.612051, 5.612032, 5.612049, 5.61203, 5.612021, 5.612119, 5.612064, 
    5.612146, 5.612142, 5.612104, 5.612143, 5.61178, 5.61177, 5.611733, 
    5.611762, 5.61171, 5.611738, 5.611754, 5.611818, 5.611834, 5.611846, 
    5.611872, 5.611905, 5.611961, 5.612011, 5.61206, 5.612057, 5.612058, 
    5.612068, 5.612042, 5.612072, 5.612077, 5.612064, 5.612142, 5.61212, 
    5.612142, 5.612128, 5.611773, 5.61179, 5.611781, 5.611798, 5.611785, 
    5.61184, 5.611857, 5.611934, 5.611904, 5.611953, 5.611909, 5.611917, 
    5.611953, 5.611912, 5.612007, 5.611941, 5.612069, 5.611997, 5.612073, 
    5.61206, 5.612082, 5.612101, 5.612125, 5.61217, 5.61216, 5.612197, 
    5.611816, 5.611838, 5.611837, 5.611861, 5.611878, 5.611916, 5.611976, 
    5.611953, 5.611995, 5.612003, 5.61194, 5.611978, 5.611854, 5.611873, 
    5.611862, 5.611817, 5.611958, 5.611886, 5.61202, 5.61198, 5.612098, 
    5.612039, 5.612154, 5.612201, 5.612248, 5.612299, 5.611851, 5.611836, 
    5.611864, 5.6119, 5.611936, 5.611982, 5.611988, 5.611996, 5.61202, 
    5.61204, 5.611998, 5.612045, 5.611876, 5.611964, 5.61183, 5.611869, 
    5.611898, 5.611887, 5.611951, 5.611966, 5.612028, 5.611996, 5.612189, 
    5.612104, 5.612341, 5.612275, 5.611831, 5.611851, 5.611922, 5.611888, 
    5.611986, 5.61201, 5.612031, 5.612056, 5.61206, 5.612075, 5.61205, 
    5.612074, 5.611982, 5.612023, 5.611915, 5.61194, 5.611929, 5.611916, 
    5.611957, 5.611999, 5.612, 5.612014, 5.612052, 5.611986, 5.612197, 
    5.612065, 5.611874, 5.611912, 5.611919, 5.611904, 5.612007, 5.611969, 
    5.612074, 5.612046, 5.612093, 5.61207, 5.612066, 5.612036, 5.612017, 
    5.611971, 5.611935, 5.611906, 5.611913, 5.611944, 5.612001, 5.61206, 
    5.612047, 5.61209, 5.611979, 5.612024, 5.612005, 5.612054, 5.611952, 
    5.612034, 5.611931, 5.611941, 5.611969, 5.612026, 5.612041, 5.612055, 
    5.612047, 5.612003, 5.611997, 5.611969, 5.61196, 5.611939, 5.611921, 
    5.611937, 5.611954, 5.612003, 5.612051, 5.612101, 5.612114, 5.612169, 
    5.612123, 5.612198, 5.612131, 5.612247, 5.612041, 5.612132, 5.61197, 
    5.611988, 5.612018, 5.612092, 5.612053, 5.612099, 5.611997, 5.611945, 
    5.611932, 5.611907, 5.611933, 5.611931, 5.611955, 5.611948, 5.612005, 
    5.611974, 5.612066, 5.612099, 5.612193, 5.612249, 5.612309, 5.612334, 
    5.612342, 5.612345 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  5.913043e-15, 5.911911e-15, 5.912125e-15, 5.911225e-15, 5.911717e-15, 
    5.911133e-15, 5.912804e-15, 5.911874e-15, 5.912462e-15, 5.912928e-15, 
    5.90951e-15, 5.911182e-15, 5.907686e-15, 5.908765e-15, 5.906031e-15, 
    5.907866e-15, 5.905658e-15, 5.906063e-15, 5.904795e-15, 5.905156e-15, 
    5.903582e-15, 5.904627e-15, 5.902733e-15, 5.90382e-15, 5.903658e-15, 
    5.904665e-15, 5.910825e-15, 5.909724e-15, 5.910895e-15, 5.910737e-15, 
    5.910803e-15, 5.911714e-15, 5.912187e-15, 5.913115e-15, 5.912942e-15, 
    5.912253e-15, 5.910665e-15, 5.91119e-15, 5.909828e-15, 5.909858e-15, 
    5.908359e-15, 5.909035e-15, 5.906503e-15, 5.907218e-15, 5.905141e-15, 
    5.905665e-15, 5.905169e-15, 5.905316e-15, 5.905167e-15, 5.905935e-15, 
    5.905607e-15, 5.906276e-15, 5.908912e-15, 5.908144e-15, 5.91045e-15, 
    5.911872e-15, 5.912767e-15, 5.913418e-15, 5.913326e-15, 5.913155e-15, 
    5.912249e-15, 5.911382e-15, 5.910727e-15, 5.910293e-15, 5.909862e-15, 
    5.908616e-15, 5.907911e-15, 5.90637e-15, 5.906629e-15, 5.906175e-15, 
    5.905716e-15, 5.904971e-15, 5.905091e-15, 5.904767e-15, 5.906174e-15, 
    5.905245e-15, 5.906783e-15, 5.906363e-15, 5.909817e-15, 5.911045e-15, 
    5.911629e-15, 5.912087e-15, 5.913256e-15, 5.912453e-15, 5.912771e-15, 
    5.911999e-15, 5.911518e-15, 5.911753e-15, 5.910281e-15, 5.910855e-15, 
    5.90787e-15, 5.909153e-15, 5.90577e-15, 5.906575e-15, 5.905575e-15, 
    5.906081e-15, 5.905219e-15, 5.905994e-15, 5.904641e-15, 5.904355e-15, 
    5.904551e-15, 5.903771e-15, 5.906039e-15, 5.905176e-15, 5.911762e-15, 
    5.911725e-15, 5.91154e-15, 5.912353e-15, 5.912399e-15, 5.913123e-15, 
    5.912472e-15, 5.912201e-15, 5.911484e-15, 5.911075e-15, 5.910681e-15, 
    5.909814e-15, 5.908859e-15, 5.907506e-15, 5.906523e-15, 5.905869e-15, 
    5.906265e-15, 5.905916e-15, 5.906309e-15, 5.90649e-15, 5.904467e-15, 
    5.905608e-15, 5.903883e-15, 5.903976e-15, 5.904762e-15, 5.903966e-15, 
    5.911697e-15, 5.911917e-15, 5.912704e-15, 5.912088e-15, 5.913201e-15, 
    5.912587e-15, 5.912239e-15, 5.910859e-15, 5.910539e-15, 5.910265e-15, 
    5.909707e-15, 5.909001e-15, 5.907767e-15, 5.906683e-15, 5.905687e-15, 
    5.905759e-15, 5.905734e-15, 5.905519e-15, 5.906061e-15, 5.905429e-15, 
    5.90533e-15, 5.9056e-15, 5.903989e-15, 5.904448e-15, 5.903978e-15, 
    5.904275e-15, 5.911844e-15, 5.91147e-15, 5.911673e-15, 5.911296e-15, 
    5.911567e-15, 5.910382e-15, 5.910026e-15, 5.908348e-15, 5.909018e-15, 
    5.907932e-15, 5.908902e-15, 5.908735e-15, 5.907926e-15, 5.908845e-15, 
    5.906758e-15, 5.908199e-15, 5.90551e-15, 5.906976e-15, 5.90542e-15, 
    5.905691e-15, 5.905235e-15, 5.904836e-15, 5.90432e-15, 5.90339e-15, 
    5.903602e-15, 5.902814e-15, 5.910908e-15, 5.910431e-15, 5.91046e-15, 
    5.909951e-15, 5.909579e-15, 5.908756e-15, 5.907452e-15, 5.907937e-15, 
    5.907032e-15, 5.906855e-15, 5.908223e-15, 5.907395e-15, 5.910102e-15, 
    5.909678e-15, 5.90992e-15, 5.910878e-15, 5.907844e-15, 5.909408e-15, 
    5.906509e-15, 5.907352e-15, 5.904895e-15, 5.906129e-15, 5.903722e-15, 
    5.902732e-15, 5.901738e-15, 5.900653e-15, 5.910156e-15, 5.910481e-15, 
    5.909887e-15, 5.909091e-15, 5.908314e-15, 5.907304e-15, 5.907193e-15, 
    5.907008e-15, 5.906511e-15, 5.906102e-15, 5.906962e-15, 5.905998e-15, 
    5.909607e-15, 5.907703e-15, 5.910617e-15, 5.909756e-15, 5.909131e-15, 
    5.909392e-15, 5.90799e-15, 5.907664e-15, 5.906348e-15, 5.907021e-15, 
    5.902988e-15, 5.90477e-15, 5.899784e-15, 5.901181e-15, 5.910598e-15, 
    5.910151e-15, 5.908616e-15, 5.909344e-15, 5.907229e-15, 5.906716e-15, 
    5.906286e-15, 5.905761e-15, 5.905694e-15, 5.905381e-15, 5.905895e-15, 
    5.905396e-15, 5.907301e-15, 5.906447e-15, 5.908775e-15, 5.908215e-15, 
    5.908468e-15, 5.908755e-15, 5.907871e-15, 5.906952e-15, 5.906911e-15, 
    5.90662e-15, 5.90584e-15, 5.90722e-15, 5.902798e-15, 5.905561e-15, 
    5.909665e-15, 5.908834e-15, 5.908689e-15, 5.909015e-15, 5.906768e-15, 
    5.907584e-15, 5.905385e-15, 5.905974e-15, 5.905005e-15, 5.905488e-15, 
    5.90556e-15, 5.906177e-15, 5.906567e-15, 5.907551e-15, 5.908345e-15, 
    5.908965e-15, 5.908819e-15, 5.908138e-15, 5.906891e-15, 5.905698e-15, 
    5.905961e-15, 5.905078e-15, 5.907383e-15, 5.906426e-15, 5.906803e-15, 
    5.905817e-15, 5.907955e-15, 5.9062e-15, 5.908412e-15, 5.908214e-15, 
    5.9076e-15, 5.906376e-15, 5.906073e-15, 5.905789e-15, 5.90596e-15, 
    5.906855e-15, 5.906993e-15, 5.90761e-15, 5.907791e-15, 5.908255e-15, 
    5.90865e-15, 5.908295e-15, 5.907926e-15, 5.906846e-15, 5.905885e-15, 
    5.904834e-15, 5.904568e-15, 5.903395e-15, 5.904379e-15, 5.902787e-15, 
    5.904184e-15, 5.901744e-15, 5.906066e-15, 5.904183e-15, 5.907565e-15, 
    5.907194e-15, 5.906547e-15, 5.905021e-15, 5.905822e-15, 5.904875e-15, 
    5.906996e-15, 5.908126e-15, 5.908391e-15, 5.908931e-15, 5.908379e-15, 
    5.908423e-15, 5.907896e-15, 5.908064e-15, 5.90681e-15, 5.907482e-15, 
    5.905567e-15, 5.904877e-15, 5.902904e-15, 5.901712e-15, 5.900467e-15, 
    5.899929e-15, 5.899764e-15, 5.899696e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  7.058777, 7.085488, 7.080293, 7.101874, 7.089901, 7.104038, 7.064192, 
    7.086545, 7.072272, 7.061187, 7.143488, 7.10284, 7.185709, 7.159791, 
    7.225058, 7.181663, 7.233835, 7.223818, 7.254036, 7.24537, 7.284096, 
    7.258039, 7.304257, 7.277875, 7.281991, 7.257178, 7.111099, 7.138443, 
    7.109459, 7.113399, 7.111634, 7.090144, 7.079324, 7.056748, 7.060845, 
    7.077434, 7.115171, 7.102352, 7.13447, 7.133749, 7.169341, 7.153276, 
    7.213317, 7.196216, 7.245732, 7.233252, 7.245143, 7.241538, 7.24519, 
    7.226894, 7.234728, 7.21865, 7.15628, 7.174561, 7.120138, 7.087057, 
    7.065169, 7.049659, 7.05185, 7.056026, 7.07753, 7.097808, 7.113287, 
    7.123577, 7.133646, 7.164152, 7.180373, 7.216771, 7.210205, 7.221342, 
    7.232012, 7.249937, 7.246986, 7.254889, 7.221057, 7.243524, 7.206463, 
    7.216583, 7.136334, 7.105811, 7.092708, 7.081289, 7.053534, 7.07269, 
    7.065132, 7.083131, 7.094581, 7.088918, 7.123857, 7.110306, 7.181334, 
    7.150729, 7.230767, 7.211553, 7.23538, 7.223217, 7.244063, 7.2253, 
    7.257836, 7.26493, 7.26008, 7.278739, 7.224259, 7.245138, 7.088758, 
    7.08968, 7.093987, 7.075071, 7.073917, 7.056633, 7.072015, 7.07857, 
    7.095248, 7.105119, 7.114516, 7.134952, 7.157749, 7.189738, 7.212797, 
    7.228283, 7.218788, 7.22717, 7.217798, 7.213411, 7.262268, 7.234798, 
    7.276053, 7.273767, 7.255075, 7.274025, 7.090329, 7.085017, 7.066585, 
    7.081007, 7.054754, 7.069434, 7.077882, 7.11058, 7.117792, 7.124378, 
    7.137384, 7.154097, 7.183487, 7.209144, 7.232635, 7.230913, 7.231519, 
    7.236769, 7.223763, 7.238906, 7.241446, 7.234801, 7.273461, 7.2624, 
    7.273718, 7.266517, 7.086745, 7.095688, 7.090854, 7.099945, 7.093535, 
    7.122001, 7.130435, 7.170018, 7.153765, 7.17966, 7.156396, 7.160511, 
    7.180485, 7.157655, 7.207718, 7.173728, 7.236973, 7.202903, 7.239111, 
    7.232533, 7.243432, 7.253197, 7.265507, 7.288247, 7.282979, 7.302035, 
    7.109042, 7.120636, 7.119637, 7.131634, 7.140515, 7.159805, 7.190817, 
    7.179146, 7.200595, 7.204903, 7.172328, 7.192306, 7.128311, 7.138609, 
    7.132483, 7.109954, 7.181821, 7.144931, 7.213177, 7.193108, 7.251803, 
    7.222557, 7.280077, 7.304749, 7.328072, 7.355347, 7.126898, 7.119115, 
    7.133065, 7.152384, 7.170373, 7.194328, 7.196788, 7.201282, 7.212942, 
    7.222753, 7.202693, 7.225214, 7.140981, 7.185034, 7.116126, 7.136835, 
    7.151248, 7.144932, 7.177815, 7.185579, 7.217194, 7.200843, 7.298645, 
    7.255248, 7.376198, 7.342238, 7.116358, 7.126876, 7.163437, 7.146025, 
    7.195935, 7.208258, 7.218296, 7.231128, 7.232522, 7.240135, 7.227661, 
    7.239645, 7.19438, 7.214582, 7.159262, 7.17269, 7.166513, 7.159736, 
    7.180668, 7.203006, 7.2035, 7.210671, 7.230885, 7.196138, 7.304233, 
    7.237303, 7.138319, 7.158547, 7.161458, 7.153612, 7.207021, 7.187631, 
    7.239951, 7.225785, 7.249012, 7.237462, 7.235763, 7.220955, 7.211744, 
    7.188516, 7.169664, 7.154751, 7.158218, 7.174608, 7.204378, 7.232641, 
    7.22644, 7.247244, 7.192307, 7.215295, 7.206398, 7.229618, 7.178833, 
    7.222015, 7.167822, 7.172564, 7.187247, 7.216846, 7.223431, 7.230439, 
    7.226117, 7.205138, 7.201712, 7.186893, 7.182798, 7.171533, 7.162209, 
    7.170723, 7.179671, 7.205153, 7.22817, 7.253334, 7.259509, 7.288977, 
    7.264961, 7.304605, 7.270858, 7.329367, 7.224547, 7.269897, 7.187921, 
    7.196721, 7.212644, 7.2493, 7.229509, 7.252666, 7.201579, 7.175167, 
    7.168364, 7.155654, 7.168654, 7.167597, 7.180052, 7.176049, 7.206001, 
    7.1899, 7.235716, 7.252487, 7.300031, 7.329284, 7.359179, 7.372397, 
    7.376426, 7.378109 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002557228, 0.0002556718, 0.0002556815, 0.000255641, 0.0002556631, 
    0.0002556368, 0.000255712, 0.0002556702, 0.0002556967, 0.0002557177, 
    0.0002555636, 0.0002556391, 0.0002554817, 0.0002555302, 0.0002554072, 
    0.0002554898, 0.0002553904, 0.0002554086, 0.0002553515, 0.0002553678, 
    0.0002552967, 0.000255344, 0.0002552585, 0.0002553075, 0.0002553002, 
    0.0002553457, 0.000255623, 0.0002555732, 0.0002556262, 0.000255619, 
    0.000255622, 0.000255663, 0.0002556842, 0.0002557261, 0.0002557183, 
    0.0002556872, 0.0002556158, 0.0002556394, 0.0002555781, 0.0002555795, 
    0.000255512, 0.0002555424, 0.0002554285, 0.0002554606, 0.0002553671, 
    0.0002553907, 0.0002553684, 0.0002553751, 0.0002553683, 0.0002554029, 
    0.0002553881, 0.0002554183, 0.0002555369, 0.0002555023, 0.0002556061, 
    0.00025567, 0.0002557104, 0.0002557397, 0.0002557356, 0.0002557278, 
    0.0002556871, 0.000255648, 0.0002556186, 0.000255599, 0.0002555797, 
    0.0002555235, 0.0002554918, 0.0002554224, 0.0002554342, 0.0002554137, 
    0.0002553931, 0.0002553595, 0.0002553649, 0.0002553503, 0.0002554137, 
    0.0002553718, 0.0002554411, 0.0002554222, 0.0002555775, 0.0002556329, 
    0.0002556591, 0.0002556798, 0.0002557324, 0.0002556962, 0.0002557106, 
    0.0002556758, 0.0002556542, 0.0002556648, 0.0002555985, 0.0002556244, 
    0.0002554899, 0.0002555477, 0.0002553955, 0.0002554317, 0.0002553867, 
    0.0002554095, 0.0002553707, 0.0002554056, 0.0002553446, 0.0002553317, 
    0.0002553406, 0.0002553054, 0.0002554076, 0.0002553687, 0.0002556652, 
    0.0002556635, 0.0002556552, 0.0002556918, 0.0002556938, 0.0002557265, 
    0.0002556971, 0.0002556849, 0.0002556527, 0.0002556343, 0.0002556165, 
    0.0002555775, 0.0002555345, 0.0002554736, 0.0002554294, 0.0002554, 
    0.0002554178, 0.0002554021, 0.0002554198, 0.0002554279, 0.0002553367, 
    0.0002553882, 0.0002553104, 0.0002553146, 0.0002553501, 0.0002553141, 
    0.0002556622, 0.0002556721, 0.0002557076, 0.0002556798, 0.0002557299, 
    0.0002557023, 0.0002556866, 0.0002556245, 0.0002556101, 0.0002555978, 
    0.0002555727, 0.0002555409, 0.0002554853, 0.0002554366, 0.0002553917, 
    0.000255395, 0.0002553939, 0.0002553842, 0.0002554086, 0.0002553801, 
    0.0002553756, 0.0002553878, 0.0002553152, 0.0002553359, 0.0002553147, 
    0.0002553281, 0.0002556689, 0.000255652, 0.0002556612, 0.0002556442, 
    0.0002556564, 0.000255603, 0.000255587, 0.0002555114, 0.0002555416, 
    0.0002554927, 0.0002555364, 0.0002555289, 0.0002554924, 0.0002555339, 
    0.0002554399, 0.0002555047, 0.0002553838, 0.0002554496, 0.0002553797, 
    0.0002553919, 0.0002553714, 0.0002553534, 0.0002553301, 0.0002552881, 
    0.0002552978, 0.0002552622, 0.0002556267, 0.0002556052, 0.0002556065, 
    0.0002555837, 0.0002555669, 0.0002555298, 0.0002554712, 0.000255493, 
    0.0002554523, 0.0002554443, 0.0002555059, 0.0002554686, 0.0002555904, 
    0.0002555713, 0.0002555822, 0.0002556254, 0.0002554888, 0.0002555591, 
    0.0002554288, 0.0002554667, 0.000255356, 0.0002554116, 0.0002553032, 
    0.0002552584, 0.0002552136, 0.0002551645, 0.0002555929, 0.0002556075, 
    0.0002555808, 0.0002555449, 0.0002555099, 0.0002554645, 0.0002554595, 
    0.0002554512, 0.0002554289, 0.0002554104, 0.0002554491, 0.0002554057, 
    0.000255568, 0.0002554824, 0.0002556136, 0.0002555748, 0.0002555467, 
    0.0002555585, 0.0002554954, 0.0002554807, 0.0002554215, 0.0002554518, 
    0.0002552699, 0.0002553504, 0.0002551252, 0.0002551884, 0.0002556128, 
    0.0002555927, 0.0002555235, 0.0002555563, 0.0002554611, 0.000255438, 
    0.0002554187, 0.000255395, 0.000255392, 0.0002553779, 0.0002554011, 
    0.0002553786, 0.0002554644, 0.000255426, 0.0002555307, 0.0002555055, 
    0.0002555169, 0.0002555298, 0.00025549, 0.0002554486, 0.0002554468, 
    0.0002554337, 0.0002553984, 0.0002554607, 0.0002552612, 0.0002553859, 
    0.0002555708, 0.0002555333, 0.0002555268, 0.0002555415, 0.0002554404, 
    0.0002554771, 0.0002553782, 0.0002554047, 0.000255361, 0.0002553828, 
    0.000255386, 0.0002554138, 0.0002554314, 0.0002554756, 0.0002555114, 
    0.0002555393, 0.0002555327, 0.000255502, 0.0002554459, 0.0002553922, 
    0.0002554041, 0.0002553643, 0.0002554681, 0.000255425, 0.0002554419, 
    0.0002553976, 0.0002554938, 0.0002554146, 0.0002555144, 0.0002555055, 
    0.0002554778, 0.0002554227, 0.0002554091, 0.0002553963, 0.000255404, 
    0.0002554443, 0.0002554505, 0.0002554783, 0.0002554864, 0.0002555073, 
    0.0002555251, 0.0002555091, 0.0002554925, 0.0002554439, 0.0002554007, 
    0.0002553533, 0.0002553413, 0.0002552883, 0.0002553327, 0.0002552607, 
    0.0002553238, 0.0002552137, 0.0002554087, 0.0002553238, 0.0002554763, 
    0.0002554596, 0.0002554304, 0.0002553617, 0.0002553978, 0.0002553551, 
    0.0002554506, 0.0002555015, 0.0002555134, 0.0002555378, 0.0002555129, 
    0.0002555149, 0.0002554911, 0.0002554987, 0.0002554423, 0.0002554726, 
    0.0002553863, 0.0002553552, 0.0002552662, 0.0002552124, 0.0002551561, 
    0.0002551318, 0.0002551244, 0.0002551213 ;

 W_SCALAR =
  0.6253964, 0.6270571, 0.6267344, 0.6280729, 0.6273305, 0.6282067, 
    0.6257331, 0.6271231, 0.6262359, 0.6255459, 0.6306667, 0.6281325, 
    0.6332931, 0.6316808, 0.6357269, 0.6330425, 0.6362674, 0.6356493, 
    0.6375082, 0.6369759, 0.6393509, 0.6377538, 0.6405799, 0.6389696, 
    0.6392217, 0.6377011, 0.6286427, 0.6303515, 0.6285414, 0.6287853, 
    0.6286758, 0.6273459, 0.6266753, 0.6252692, 0.6255246, 0.6265572, 
    0.6288949, 0.6281016, 0.6300995, 0.6300544, 0.6322752, 0.6312743, 
    0.6350011, 0.633943, 0.6369982, 0.6362305, 0.6369621, 0.6367403, 
    0.636965, 0.635839, 0.6363216, 0.6353303, 0.6314619, 0.6326001, 
    0.6292027, 0.6271558, 0.6257942, 0.6248273, 0.624964, 0.6252246, 
    0.6265632, 0.6278204, 0.6287776, 0.6294177, 0.6300479, 0.6319543, 
    0.6329618, 0.6352151, 0.6348086, 0.635497, 0.6361542, 0.6372568, 
    0.6370754, 0.637561, 0.6354787, 0.6368631, 0.634577, 0.6352027, 
    0.6302198, 0.6283157, 0.627506, 0.6267965, 0.6250691, 0.6262622, 
    0.625792, 0.6269103, 0.6276205, 0.6272693, 0.6294351, 0.6285936, 
    0.6330215, 0.6311161, 0.6360775, 0.634892, 0.6363615, 0.6356118, 
    0.6368961, 0.6357403, 0.6377416, 0.638177, 0.6378795, 0.6390218, 
    0.6356763, 0.6369622, 0.6272594, 0.6273167, 0.6275835, 0.6264104, 
    0.6263385, 0.6252623, 0.6262199, 0.6266276, 0.6276616, 0.628273, 
    0.6288538, 0.6301301, 0.631554, 0.6335424, 0.6349689, 0.6359242, 
    0.6353385, 0.6358557, 0.6352775, 0.6350065, 0.6380139, 0.6363261, 
    0.6388575, 0.6387176, 0.6375725, 0.6387333, 0.6273569, 0.6270273, 
    0.6258821, 0.6267784, 0.625145, 0.6260596, 0.6265852, 0.6286113, 
    0.6290559, 0.6294681, 0.6302819, 0.6313256, 0.6331545, 0.6347436, 
    0.6361923, 0.6360862, 0.6361236, 0.6364471, 0.6356457, 0.6365786, 
    0.6367351, 0.6363259, 0.6386988, 0.6380213, 0.6387146, 0.6382735, 
    0.6271344, 0.6276891, 0.6273894, 0.6279529, 0.627556, 0.6293201, 
    0.6298485, 0.6323183, 0.6313051, 0.632917, 0.6314689, 0.6317256, 
    0.6329699, 0.6315472, 0.6346561, 0.6325494, 0.6364596, 0.6343591, 
    0.6365912, 0.6361861, 0.6368567, 0.6374571, 0.6382118, 0.6396034, 
    0.6392813, 0.640444, 0.6285154, 0.629234, 0.6291707, 0.6299223, 
    0.6304778, 0.6316811, 0.6336089, 0.6328843, 0.6342141, 0.6344809, 
    0.6324604, 0.6337014, 0.6297147, 0.6303598, 0.6299756, 0.6285722, 
    0.6330515, 0.6307546, 0.6349925, 0.6337506, 0.6373715, 0.6355722, 
    0.6391039, 0.6406109, 0.6420269, 0.6436802, 0.629626, 0.6291379, 
    0.6300116, 0.6312197, 0.6323393, 0.6338264, 0.6339784, 0.6342568, 
    0.6349776, 0.6355833, 0.634345, 0.635735, 0.6305096, 0.6332505, 
    0.6289534, 0.630249, 0.6311485, 0.6307539, 0.6328014, 0.6332836, 
    0.635241, 0.6342294, 0.6402392, 0.637584, 0.644937, 0.6428869, 0.6289673, 
    0.6296242, 0.6319082, 0.6308219, 0.6339256, 0.6346884, 0.6353081, 
    0.6361001, 0.6361854, 0.6366544, 0.6358859, 0.636624, 0.6338296, 
    0.6350791, 0.6316472, 0.6324834, 0.6320987, 0.6316767, 0.6329787, 
    0.6343645, 0.6343939, 0.634838, 0.6360888, 0.6339381, 0.6405819, 
    0.6364834, 0.6303402, 0.6316042, 0.6317844, 0.631295, 0.634612, 
    0.6334112, 0.6366429, 0.6357703, 0.6371997, 0.6364896, 0.6363851, 
    0.6354724, 0.6349038, 0.6334662, 0.6322954, 0.631366, 0.6315821, 
    0.6326028, 0.6344492, 0.6361933, 0.6358114, 0.6370911, 0.6337008, 
    0.6351237, 0.634574, 0.6360067, 0.6328651, 0.6355414, 0.6321801, 
    0.6324751, 0.6333873, 0.6352202, 0.6356251, 0.6360576, 0.6357907, 
    0.634496, 0.6342837, 0.6333651, 0.6331115, 0.6324109, 0.6318307, 
    0.6323609, 0.6329174, 0.6344965, 0.6359178, 0.6374656, 0.637844, 
    0.6396499, 0.6381803, 0.6406047, 0.6385442, 0.6421086, 0.6356961, 
    0.6384832, 0.6334288, 0.6339742, 0.6349604, 0.637219, 0.636, 0.6374254, 
    0.6342753, 0.6326381, 0.632214, 0.6314225, 0.632232, 0.6321662, 
    0.6329404, 0.6326916, 0.6345488, 0.6335515, 0.6363825, 0.6374141, 
    0.6403223, 0.6421017, 0.6439101, 0.6447076, 0.6449502, 0.6450517,
  0.5466837, 0.5487262, 0.5483293, 0.5499756, 0.5490624, 0.5501403, 
    0.5470979, 0.5488074, 0.5477161, 0.5468675, 0.5531667, 0.550049, 
    0.5563989, 0.5544147, 0.5593947, 0.5560904, 0.5600601, 0.5592992, 
    0.5615879, 0.5609326, 0.5638572, 0.5618904, 0.565371, 0.5633876, 
    0.5636981, 0.5618255, 0.5506766, 0.552779, 0.5505521, 0.550852, 
    0.5507174, 0.5490814, 0.5482566, 0.5465273, 0.5468413, 0.5481113, 
    0.5509868, 0.550011, 0.5524688, 0.5524134, 0.5551461, 0.5539145, 
    0.5585013, 0.5571988, 0.5609599, 0.5600148, 0.5609156, 0.5606425, 
    0.5609191, 0.5595328, 0.560127, 0.5589065, 0.5541453, 0.5555459, 
    0.5513654, 0.5488476, 0.5471729, 0.5459838, 0.5461519, 0.5464725, 
    0.5481187, 0.549665, 0.5508426, 0.55163, 0.5524054, 0.5547512, 0.5559911, 
    0.5587647, 0.5582643, 0.5591118, 0.5599208, 0.5612784, 0.561055, 
    0.561653, 0.5590892, 0.5607936, 0.5579792, 0.5587494, 0.552617, 
    0.5502743, 0.5492784, 0.5484056, 0.5462812, 0.5477486, 0.5471703, 
    0.5485456, 0.5494191, 0.5489872, 0.5516515, 0.5506161, 0.5560646, 
    0.5537197, 0.5598264, 0.558367, 0.560176, 0.5592531, 0.5608342, 
    0.5594113, 0.5618753, 0.5624115, 0.5620452, 0.5634518, 0.5593324, 
    0.5609156, 0.5489751, 0.5490455, 0.5493737, 0.5479307, 0.5478424, 
    0.5465187, 0.5476965, 0.5481979, 0.5494697, 0.5502217, 0.5509363, 
    0.5525064, 0.5542586, 0.5567057, 0.5584616, 0.5596377, 0.5589166, 
    0.5595533, 0.5588415, 0.5585079, 0.5622107, 0.5601325, 0.5632496, 
    0.5630772, 0.5616672, 0.5630966, 0.549095, 0.5486895, 0.5472811, 
    0.5483834, 0.5463746, 0.5474994, 0.5481458, 0.550638, 0.5511849, 
    0.5516921, 0.5526933, 0.5539775, 0.5562283, 0.5581842, 0.5599678, 
    0.5598372, 0.5598831, 0.5602815, 0.5592948, 0.5604433, 0.5606361, 
    0.5601322, 0.5630541, 0.5622199, 0.5630736, 0.5625304, 0.5488213, 
    0.5495035, 0.5491349, 0.549828, 0.5493398, 0.5515099, 0.5521601, 
    0.5551991, 0.5539523, 0.555936, 0.5541539, 0.5544698, 0.5560011, 
    0.5542502, 0.5580766, 0.5554836, 0.5602969, 0.557711, 0.5604588, 
    0.5599601, 0.5607857, 0.561525, 0.5624543, 0.5641682, 0.5637714, 
    0.5652035, 0.55052, 0.5514041, 0.5513262, 0.5522508, 0.5529345, 
    0.5544151, 0.5567876, 0.5558957, 0.5575324, 0.5578609, 0.5553741, 
    0.5569015, 0.5519955, 0.5527891, 0.5523165, 0.5505899, 0.5561014, 
    0.553275, 0.5584906, 0.556962, 0.5614196, 0.5592043, 0.563553, 0.5654091, 
    0.5671535, 0.5691905, 0.5518863, 0.5512857, 0.5523607, 0.5538473, 
    0.555225, 0.5570553, 0.5572424, 0.5575851, 0.5584723, 0.5592179, 
    0.5576936, 0.5594048, 0.5529734, 0.5563465, 0.5510588, 0.5526528, 
    0.5537596, 0.553274, 0.5557937, 0.5563871, 0.5587966, 0.5575513, 
    0.5649514, 0.5616813, 0.5707393, 0.568213, 0.5510759, 0.5518841, 
    0.5546944, 0.5533578, 0.5571774, 0.5581164, 0.5588793, 0.5598541, 
    0.5599593, 0.5605366, 0.5595905, 0.5604992, 0.5570592, 0.5585973, 
    0.5543733, 0.5554023, 0.554929, 0.5544096, 0.5560119, 0.5577176, 
    0.5577538, 0.5583004, 0.5598403, 0.5571928, 0.5653734, 0.5603262, 
    0.552765, 0.5543203, 0.5545421, 0.5539399, 0.5580223, 0.5565442, 
    0.5605225, 0.5594481, 0.5612081, 0.5603338, 0.5602051, 0.5590814, 
    0.5583815, 0.556612, 0.5551709, 0.5540273, 0.5542932, 0.5555493, 
    0.5578219, 0.5599689, 0.5594988, 0.5610744, 0.5569007, 0.5586521, 
    0.5579755, 0.5597392, 0.555872, 0.5591664, 0.5550291, 0.5553922, 
    0.5565148, 0.558771, 0.5592694, 0.5598019, 0.5594733, 0.5578794, 
    0.5576181, 0.5564875, 0.5561753, 0.5553131, 0.5545991, 0.5552515, 
    0.5559365, 0.55788, 0.5596299, 0.5615355, 0.5620015, 0.5642254, 
    0.5624156, 0.5654016, 0.5628638, 0.5672541, 0.5593567, 0.5627885, 
    0.5565658, 0.5572372, 0.5584512, 0.5612318, 0.5597309, 0.5614859, 
    0.5576078, 0.5555927, 0.5550707, 0.5540968, 0.555093, 0.555012, 
    0.5559647, 0.5556586, 0.5579445, 0.556717, 0.5602019, 0.5614721, 
    0.5650536, 0.5672457, 0.5694737, 0.5704566, 0.5707555, 0.5708805,
  0.5141778, 0.5164276, 0.5159903, 0.5178041, 0.516798, 0.5179855, 0.514634, 
    0.516517, 0.515315, 0.5143803, 0.521321, 0.517885, 0.5248847, 0.5226967, 
    0.5281894, 0.5245445, 0.5289236, 0.528084, 0.5306097, 0.5298863, 
    0.5331147, 0.5309434, 0.5347862, 0.5325962, 0.532939, 0.5308718, 
    0.5185766, 0.5208935, 0.5184393, 0.5187698, 0.5186214, 0.5168189, 
    0.5159103, 0.5140056, 0.5143514, 0.5157502, 0.5189184, 0.5178432, 
    0.5205517, 0.5204906, 0.5235032, 0.5221453, 0.5272037, 0.5257669, 
    0.5299165, 0.5288736, 0.5298676, 0.5295662, 0.5298715, 0.5283418, 
    0.5289973, 0.5276507, 0.5223997, 0.5239441, 0.5193356, 0.5165614, 
    0.5147166, 0.5134071, 0.5135922, 0.5139452, 0.5157584, 0.5174619, 
    0.5187595, 0.5196272, 0.5204818, 0.5230678, 0.524435, 0.5274943, 
    0.5269422, 0.5278772, 0.5287698, 0.530268, 0.5300214, 0.5306814, 
    0.5278524, 0.5297329, 0.5266278, 0.5274774, 0.5207149, 0.5181332, 
    0.5170359, 0.5160744, 0.5137346, 0.5153507, 0.5147138, 0.5162287, 
    0.517191, 0.516715, 0.5196509, 0.5185099, 0.524516, 0.5219306, 0.5286657, 
    0.5270555, 0.5290515, 0.5280331, 0.5297778, 0.5282077, 0.5309269, 
    0.5315187, 0.5311143, 0.5326671, 0.5281206, 0.5298676, 0.5167018, 
    0.5167794, 0.5171409, 0.5155513, 0.515454, 0.5139962, 0.5152933, 
    0.5158455, 0.5172467, 0.5180753, 0.5188627, 0.5205932, 0.5225247, 
    0.5252231, 0.5271599, 0.5284575, 0.5276619, 0.5283643, 0.5275791, 
    0.527211, 0.531297, 0.5290034, 0.5324438, 0.5322536, 0.5306971, 0.532275, 
    0.5168339, 0.5163872, 0.5148358, 0.5160499, 0.5138373, 0.5150762, 
    0.5157883, 0.5185339, 0.5191366, 0.5196956, 0.5207992, 0.5222148, 
    0.5246965, 0.5268539, 0.5288217, 0.5286775, 0.5287283, 0.5291678, 
    0.5280792, 0.5293465, 0.5295592, 0.5290031, 0.5322281, 0.5313071, 
    0.5322495, 0.5316499, 0.5165324, 0.5172839, 0.5168778, 0.5176415, 
    0.5171036, 0.5194948, 0.5202114, 0.5235617, 0.522187, 0.5243742, 
    0.5224092, 0.5227575, 0.524446, 0.5225154, 0.5267352, 0.5238753, 
    0.5291849, 0.5263319, 0.5293636, 0.5288132, 0.5297243, 0.5305401, 
    0.531566, 0.533458, 0.53302, 0.5346013, 0.5184039, 0.5193782, 0.5192923, 
    0.5203114, 0.5210649, 0.5226972, 0.5253133, 0.5243298, 0.526135, 
    0.5264972, 0.5237545, 0.525439, 0.5200299, 0.5209047, 0.5203838, 
    0.5184809, 0.5245567, 0.5214403, 0.5271919, 0.5255058, 0.5304238, 
    0.5279793, 0.5327788, 0.5348283, 0.5367549, 0.5390055, 0.5199096, 
    0.5192478, 0.5204325, 0.5220711, 0.5235902, 0.5256087, 0.525815, 
    0.526193, 0.5271717, 0.5279943, 0.5263127, 0.5282005, 0.5211079, 
    0.5248269, 0.5189977, 0.5207545, 0.5219745, 0.5214393, 0.5242173, 
    0.5248717, 0.5275294, 0.5261558, 0.5343228, 0.5307127, 0.5407171, 
    0.5379254, 0.5190166, 0.5199072, 0.5230052, 0.5215316, 0.5257433, 
    0.5267791, 0.5276207, 0.5286963, 0.5288123, 0.5294494, 0.5284054, 
    0.5294081, 0.525613, 0.5273096, 0.5226511, 0.5237857, 0.5232638, 
    0.5226912, 0.5244579, 0.5263392, 0.5263791, 0.5269821, 0.528681, 
    0.5257604, 0.5347888, 0.5292172, 0.5208782, 0.5225928, 0.5228373, 
    0.5221733, 0.5266752, 0.5250449, 0.5294338, 0.5282483, 0.5301904, 
    0.5292255, 0.5290835, 0.5278437, 0.5270716, 0.5251198, 0.5235305, 
    0.5222696, 0.5225628, 0.5239478, 0.5264542, 0.5288229, 0.5283043, 
    0.5300428, 0.5254381, 0.5273701, 0.5266236, 0.5285695, 0.5243037, 
    0.5279375, 0.5233742, 0.5237746, 0.5250126, 0.5275012, 0.5280511, 
    0.5286386, 0.5282761, 0.5265177, 0.5262294, 0.5249824, 0.5246381, 
    0.5236874, 0.5229001, 0.5236195, 0.5243748, 0.5265183, 0.5284488, 
    0.5305518, 0.5310661, 0.5335212, 0.5315232, 0.5348199, 0.5320178, 
    0.5368661, 0.5281475, 0.5319349, 0.5250688, 0.5258093, 0.5271484, 
    0.5302166, 0.5285603, 0.5304971, 0.5262181, 0.5239957, 0.5234201, 
    0.5223463, 0.5234446, 0.5233553, 0.5244059, 0.5240683, 0.5265895, 
    0.5252355, 0.5290801, 0.5304818, 0.5344357, 0.5368568, 0.5393184, 
    0.5404046, 0.5407351, 0.5408732,
  0.507082, 0.5094725, 0.5090078, 0.5109357, 0.5098662, 0.5111286, 0.5075666, 
    0.5095675, 0.5082902, 0.507297, 0.5146761, 0.5110217, 0.5184693, 
    0.5161401, 0.5219896, 0.5181071, 0.5227721, 0.5218773, 0.5245695, 
    0.5237983, 0.5272413, 0.5249254, 0.529025, 0.5266882, 0.5270539, 
    0.5248491, 0.511757, 0.5142213, 0.511611, 0.5119625, 0.5118047, 
    0.5098884, 0.5089227, 0.5068991, 0.5072665, 0.5087526, 0.5121205, 
    0.5109772, 0.5138577, 0.5137926, 0.5169985, 0.5155532, 0.5209394, 
    0.5194088, 0.5238305, 0.5227188, 0.5237783, 0.5234571, 0.5237826, 
    0.522152, 0.5228506, 0.5214156, 0.515824, 0.5174678, 0.5125642, 
    0.5096147, 0.5076544, 0.5062633, 0.50646, 0.5068349, 0.5087613, 
    0.5105719, 0.5119515, 0.5128742, 0.5137833, 0.516535, 0.5179905, 
    0.5212489, 0.5206608, 0.5216569, 0.5226082, 0.5242053, 0.5239424, 
    0.524646, 0.5216305, 0.5236348, 0.5203258, 0.521231, 0.5140313, 
    0.5112856, 0.5101191, 0.5090972, 0.5066112, 0.5083281, 0.5076513, 
    0.5092611, 0.5102839, 0.509778, 0.5128995, 0.5116861, 0.5180768, 
    0.5153247, 0.5224972, 0.5207815, 0.5229084, 0.5218231, 0.5236827, 
    0.5220091, 0.5249078, 0.5255389, 0.5251076, 0.5267639, 0.5219163, 
    0.5237784, 0.5097639, 0.5098464, 0.5102307, 0.5085412, 0.5084379, 
    0.506889, 0.5082671, 0.5088539, 0.5103431, 0.511224, 0.5120613, 
    0.5139018, 0.5159569, 0.5188296, 0.5208927, 0.5222753, 0.5214275, 
    0.522176, 0.5213393, 0.520947, 0.5253025, 0.5228572, 0.5265256, 
    0.5263227, 0.5246627, 0.5263456, 0.5099043, 0.5094295, 0.507781, 
    0.5090711, 0.5067203, 0.5080364, 0.5087931, 0.5117117, 0.5123526, 
    0.5129471, 0.5141209, 0.5156272, 0.5182689, 0.5205667, 0.5226635, 
    0.5225099, 0.5225639, 0.5230324, 0.5218721, 0.5232228, 0.5234496, 
    0.5228568, 0.5262955, 0.5253133, 0.5263184, 0.5256788, 0.5095838, 
    0.5103827, 0.5099511, 0.5107628, 0.510191, 0.5127335, 0.5134957, 
    0.5170608, 0.5155976, 0.5179258, 0.515834, 0.5162048, 0.5180022, 
    0.515947, 0.5204402, 0.5173946, 0.5230506, 0.5200107, 0.523241, 
    0.5226544, 0.5236256, 0.5244954, 0.5255893, 0.5276076, 0.5271403, 
    0.5288277, 0.5115735, 0.5126095, 0.5125181, 0.5136021, 0.5144036, 
    0.5161406, 0.5189257, 0.5178785, 0.5198008, 0.5201867, 0.5172661, 
    0.5190596, 0.5133026, 0.5142332, 0.513679, 0.5116553, 0.5181201, 
    0.5148031, 0.5209268, 0.5191307, 0.5243714, 0.5217657, 0.526883, 0.52907, 
    0.5311269, 0.5335307, 0.5131747, 0.5124708, 0.5137309, 0.5154743, 
    0.5170911, 0.5192403, 0.5194601, 0.5198627, 0.5209052, 0.5217817, 
    0.5199901, 0.5220014, 0.5144494, 0.5184078, 0.5122048, 0.5140734, 
    0.5153715, 0.5148019, 0.5177587, 0.5184555, 0.5212864, 0.519823, 
    0.5285304, 0.5246793, 0.5353599, 0.5323769, 0.5122249, 0.5131721, 
    0.5164683, 0.5149001, 0.5193837, 0.520487, 0.5213836, 0.5225298, 
    0.5226535, 0.5233325, 0.5222198, 0.5232885, 0.5192448, 0.5210521, 
    0.5160915, 0.5172992, 0.5167436, 0.5161341, 0.5180149, 0.5200184, 
    0.5200609, 0.5207033, 0.5225136, 0.5194018, 0.5290278, 0.523085, 
    0.514205, 0.5160294, 0.5162897, 0.515583, 0.5203764, 0.5186399, 0.523316, 
    0.5220524, 0.5241225, 0.5230939, 0.5229426, 0.5216212, 0.5207986, 
    0.5187196, 0.5170276, 0.5156855, 0.5159976, 0.5174718, 0.5201408, 
    0.5226648, 0.522112, 0.5239652, 0.5190586, 0.5211166, 0.5203214, 
    0.5223947, 0.5178507, 0.5217211, 0.5168611, 0.5172873, 0.5186055, 
    0.5212563, 0.5218423, 0.5224684, 0.522082, 0.5202085, 0.5199015, 
    0.5185733, 0.5182068, 0.5171945, 0.5163565, 0.5171223, 0.5179264, 
    0.5202093, 0.522266, 0.5245078, 0.5250562, 0.5276751, 0.5255436, 
    0.529061, 0.5260713, 0.5312455, 0.521945, 0.5259827, 0.5186654, 
    0.5194539, 0.5208804, 0.5241504, 0.5223849, 0.5244495, 0.5198894, 
    0.5175228, 0.51691, 0.5157672, 0.5169361, 0.5168411, 0.5179595, 
    0.5176001, 0.520285, 0.5188429, 0.5229388, 0.5244331, 0.5286509, 
    0.5312356, 0.5338652, 0.5350259, 0.5353791, 0.5355268,
  0.5310288, 0.5334982, 0.5330179, 0.5350106, 0.533905, 0.5352101, 0.5315292, 
    0.5335963, 0.5322765, 0.5312509, 0.5388809, 0.5350995, 0.5428115, 
    0.5403972, 0.5464646, 0.5424359, 0.5472774, 0.546348, 0.5491452, 
    0.5483436, 0.5519241, 0.5495151, 0.5537811, 0.5513485, 0.5517291, 
    0.5494357, 0.5358599, 0.53841, 0.535709, 0.5360725, 0.5359093, 0.5339279, 
    0.53293, 0.5308399, 0.5312192, 0.5327542, 0.5362359, 0.5350536, 
    0.5380336, 0.5379663, 0.5412867, 0.5397893, 0.5453742, 0.543786, 
    0.548377, 0.547222, 0.5483229, 0.547989, 0.5483272, 0.5466332, 0.5473589, 
    0.5458686, 0.5400697, 0.5417732, 0.536695, 0.533645, 0.5316198, 
    0.5301836, 0.5303866, 0.5307737, 0.5327632, 0.5346345, 0.5360612, 
    0.5370158, 0.5379566, 0.5408065, 0.5423151, 0.5456956, 0.5450851, 
    0.5461192, 0.5471071, 0.5487665, 0.5484933, 0.5492246, 0.5460917, 
    0.5481737, 0.5447374, 0.545677, 0.5382133, 0.5353725, 0.5341663, 
    0.5331103, 0.5305427, 0.5323157, 0.5316167, 0.5332797, 0.5343367, 
    0.5338138, 0.5370419, 0.5357866, 0.5424045, 0.5395526, 0.5469918, 
    0.5452104, 0.547419, 0.5462917, 0.5482234, 0.5464849, 0.5494968, 
    0.5501531, 0.5497046, 0.5514272, 0.5463886, 0.5483229, 0.5337992, 
    0.5338845, 0.5342818, 0.5325359, 0.5324291, 0.5308296, 0.5322527, 
    0.532859, 0.534398, 0.5353088, 0.5361747, 0.5380793, 0.5402075, 
    0.5431852, 0.5453258, 0.5467613, 0.545881, 0.5466582, 0.5457894, 
    0.5453822, 0.5499072, 0.5473658, 0.5511795, 0.5509683, 0.5492421, 
    0.5509921, 0.5339444, 0.5334537, 0.5317506, 0.5330834, 0.5306554, 
    0.5320144, 0.5327961, 0.5358131, 0.536476, 0.5370911, 0.5383061, 
    0.5398659, 0.5426038, 0.5449874, 0.5471645, 0.5470049, 0.5470611, 
    0.5475478, 0.5463426, 0.5477456, 0.5479812, 0.5473654, 0.55094, 
    0.5499184, 0.5509638, 0.5502986, 0.5336131, 0.5344389, 0.5339927, 
    0.5348319, 0.5342407, 0.5368702, 0.5376589, 0.5413513, 0.5398352, 
    0.542248, 0.5400802, 0.5404643, 0.5423271, 0.5401973, 0.5448561, 
    0.5416973, 0.5475667, 0.5444103, 0.5477645, 0.5471551, 0.5481641, 
    0.5490681, 0.5502055, 0.5523053, 0.551819, 0.5535756, 0.5356702, 
    0.5367419, 0.5366473, 0.537769, 0.5385988, 0.5403978, 0.5432849, 
    0.5421989, 0.5441927, 0.5445932, 0.541564, 0.5434238, 0.5374591, 
    0.5384223, 0.5378487, 0.5357548, 0.5424494, 0.5390124, 0.5453612, 
    0.5434975, 0.5489392, 0.5462322, 0.5515513, 0.5538279, 0.555971, 
    0.5584781, 0.5373267, 0.5365984, 0.5379024, 0.5397075, 0.5413827, 
    0.5436112, 0.5438392, 0.5442569, 0.5453388, 0.5462488, 0.5443891, 
    0.546477, 0.5386461, 0.5427478, 0.5363232, 0.5382569, 0.539601, 
    0.5390112, 0.5420747, 0.5427972, 0.5457345, 0.5442157, 0.553266, 
    0.5492593, 0.5603875, 0.5572744, 0.536344, 0.5373241, 0.5407374, 
    0.5391129, 0.5437599, 0.5449046, 0.5458354, 0.5470257, 0.5471541, 
    0.5478595, 0.5467036, 0.5478138, 0.5436159, 0.5454913, 0.5403469, 
    0.5415984, 0.5410226, 0.5403911, 0.5423403, 0.5444184, 0.5444626, 
    0.5451292, 0.5470088, 0.5437787, 0.553784, 0.5476024, 0.5383931, 
    0.5402825, 0.5405522, 0.5398202, 0.5447899, 0.5429885, 0.5478423, 
    0.5465299, 0.5486805, 0.5476117, 0.5474545, 0.5460821, 0.5452281, 
    0.5430711, 0.5413169, 0.5399263, 0.5402496, 0.5417773, 0.5445455, 
    0.5471659, 0.5465918, 0.548517, 0.5434228, 0.5455582, 0.5447328, 
    0.5468853, 0.5421701, 0.5461859, 0.5411444, 0.5415861, 0.5429527, 
    0.5457033, 0.5463117, 0.5469618, 0.5465606, 0.5446157, 0.5442971, 
    0.5429195, 0.5425393, 0.5414899, 0.5406215, 0.541415, 0.5422486, 
    0.5446165, 0.5467517, 0.549081, 0.5496511, 0.5523756, 0.550158, 
    0.5538185, 0.5507067, 0.5560948, 0.5464183, 0.5506147, 0.5430148, 
    0.5438328, 0.545313, 0.5487095, 0.5468752, 0.5490203, 0.5442846, 
    0.5418302, 0.541195, 0.5400109, 0.5412221, 0.5411236, 0.5422829, 
    0.5419103, 0.5446951, 0.5431989, 0.5474506, 0.5490034, 0.5533915, 
    0.5560843, 0.558827, 0.5600387, 0.5604075, 0.5605617,
  0.535215, 0.5380583, 0.537505, 0.5398022, 0.5385273, 0.5400323, 0.5357908, 
    0.5381714, 0.5366511, 0.5354705, 0.5442734, 0.5399048, 0.5488272, 
    0.5460286, 0.5530714, 0.5483914, 0.5540173, 0.5529358, 0.5561932, 
    0.555259, 0.5594366, 0.5566247, 0.5616078, 0.5587642, 0.5592087, 
    0.5565321, 0.5407823, 0.5437287, 0.5406081, 0.5410277, 0.5408393, 
    0.5385537, 0.5374036, 0.5349978, 0.5354341, 0.5372012, 0.5412164, 
    0.5398518, 0.5432935, 0.5432156, 0.5470591, 0.5453246, 0.5518034, 
    0.5499582, 0.555298, 0.5539528, 0.5552348, 0.5548459, 0.5552399, 
    0.5532677, 0.5541123, 0.5523782, 0.5456493, 0.5476229, 0.5417466, 
    0.5382276, 0.5358952, 0.5342429, 0.5344764, 0.5349216, 0.5372116, 
    0.5393683, 0.5410146, 0.5421172, 0.5432045, 0.5465026, 0.5482513, 
    0.552177, 0.5514672, 0.5526696, 0.5538191, 0.5557519, 0.5554335, 
    0.5562859, 0.5526377, 0.5550611, 0.5510632, 0.5521553, 0.5435013, 
    0.5402197, 0.5388285, 0.5376113, 0.5346559, 0.5366961, 0.5358915, 
    0.5378065, 0.539025, 0.5384222, 0.5421473, 0.5406978, 0.548355, 
    0.5450506, 0.5536849, 0.5516129, 0.5541821, 0.5528703, 0.555119, 
    0.553095, 0.5566033, 0.5573688, 0.5568456, 0.5588562, 0.5529829, 
    0.555235, 0.5384053, 0.5385036, 0.5389616, 0.5369498, 0.5368267, 
    0.5349858, 0.5366237, 0.5373218, 0.5390956, 0.5401462, 0.5411457, 
    0.5433463, 0.5458089, 0.5492609, 0.5517471, 0.5534167, 0.5523925, 
    0.5532967, 0.5522861, 0.5518126, 0.5570819, 0.5541202, 0.5585667, 
    0.5583202, 0.5563062, 0.558348, 0.5385727, 0.538007, 0.5360457, 
    0.5375804, 0.5347855, 0.5363493, 0.5372494, 0.5407283, 0.5414937, 
    0.5422042, 0.5436085, 0.5454133, 0.5485862, 0.5513538, 0.5538859, 
    0.5537002, 0.5537656, 0.5543321, 0.5529295, 0.5545625, 0.5548369, 
    0.5541198, 0.5582872, 0.557095, 0.558315, 0.5575385, 0.5381908, 
    0.5391428, 0.5386283, 0.539596, 0.5389143, 0.5419489, 0.5428603, 
    0.5471339, 0.5453779, 0.5481735, 0.5456614, 0.5461062, 0.5482653, 
    0.545797, 0.5512012, 0.5475349, 0.5543541, 0.5506833, 0.5545846, 
    0.553875, 0.55505, 0.5561034, 0.55743, 0.559882, 0.5593137, 0.5613673, 
    0.5405633, 0.5418007, 0.5416915, 0.5429876, 0.5439471, 0.5460292, 
    0.5493765, 0.5481166, 0.5504305, 0.5508956, 0.5473805, 0.5495377, 
    0.5426294, 0.543743, 0.5430797, 0.540661, 0.5484071, 0.5444255, 
    0.5517883, 0.5496233, 0.5559531, 0.552801, 0.559001, 0.5616626, 
    0.5641724, 0.5671141, 0.5424764, 0.541635, 0.5431418, 0.54523, 0.5471703, 
    0.5497553, 0.5500199, 0.550505, 0.5517622, 0.5528204, 0.5506586, 
    0.5530857, 0.5440018, 0.5487532, 0.5413172, 0.5435517, 0.5451067, 
    0.5444241, 0.5479726, 0.5488106, 0.5522222, 0.5504572, 0.5610052, 
    0.5563263, 0.5693585, 0.5657009, 0.5413412, 0.5424734, 0.5464225, 
    0.5445418, 0.5499279, 0.5512576, 0.5523396, 0.5537243, 0.5538738, 
    0.5546952, 0.5533496, 0.554642, 0.5497608, 0.5519395, 0.5459703, 
    0.5474204, 0.546753, 0.5460215, 0.5482807, 0.5506927, 0.5507439, 
    0.5515185, 0.5537046, 0.5499498, 0.5616112, 0.5543957, 0.5437092, 
    0.5458958, 0.546208, 0.5453604, 0.5511243, 0.5490325, 0.5546752, 
    0.5531473, 0.5556517, 0.5544065, 0.5542235, 0.5526266, 0.5516335, 
    0.5491284, 0.547094, 0.5454832, 0.5458576, 0.5476277, 0.5508403, 
    0.5538875, 0.5532194, 0.5554611, 0.5495365, 0.5520173, 0.5510579, 
    0.553561, 0.5480832, 0.5527471, 0.5468942, 0.5474061, 0.548991, 0.552186, 
    0.5528935, 0.5536501, 0.5531831, 0.5509219, 0.5505518, 0.5489524, 
    0.5485114, 0.5472946, 0.5462883, 0.5472078, 0.5481742, 0.5509228, 
    0.5534055, 0.5561185, 0.5567833, 0.5599641, 0.5573745, 0.5616516, 
    0.5580149, 0.5643175, 0.5530175, 0.5579075, 0.5490631, 0.5500126, 
    0.5517322, 0.5556855, 0.5535492, 0.5560478, 0.5505372, 0.547689, 
    0.5469528, 0.5455812, 0.5469842, 0.54687, 0.548214, 0.5477819, 0.5510141, 
    0.5492768, 0.554219, 0.5560279, 0.561152, 0.5643053, 0.567524, 0.5689483, 
    0.5693821, 0.5695636,
  0.5840928, 0.5875039, 0.586839, 0.5896026, 0.5880677, 0.5898799, 0.5847825, 
    0.5876399, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057424, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041865, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048915, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.58908, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046446, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052099, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834237, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924328, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.603953, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912229, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041979, 0.6106832, 0.6070316, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065955, 0.6072922, 0.6055682, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106994, 0.6122084, 0.6112477, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.592193, 0.593295, 0.598482, 0.5963469, 
    0.5997487, 0.5966913, 0.5972319, 0.5998606, 0.596856, 0.6034486, 
    0.5989705, 0.6073194, 0.6028146, 0.607603, 0.6067299, 0.6081761, 
    0.6094749, 0.6111134, 0.614151, 0.6134459, 0.6159967, 0.59052, 0.5920138, 
    0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 0.5996793, 
    0.6025052, 0.6030745, 0.5987824, 0.6014137, 0.5930157, 0.5943638, 
    0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 0.6015183, 
    0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 0.6231793, 
    0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 0.6016796, 
    0.6020032, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 0.5946774, 
    0.6004559, 0.5914299, 0.5941321, 0.5960177, 0.5951895, 0.5995038, 
    0.6005259, 0.6047001, 0.6025379, 0.6155463, 0.60975, 0.6260031, 
    0.6214069, 0.5914588, 0.592827, 0.5976165, 0.5953323, 0.6018906, 
    0.6035177, 0.604844, 0.6065448, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980185, 
    0.5971288, 0.5998793, 0.6028261, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073706, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039783, 0.6009138, 0.5984336, 0.5964749, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014124, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007462, 0.6046556, 0.6055239, 0.6064534, 
    0.6058796, 0.6031066, 0.6026536, 0.600699, 0.6001608, 0.5986778, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103142, 0.6142529, 0.6110448, 0.6163503, 0.6118369, 0.6196756, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040993, 0.6089594, 
    0.6063294, 0.6094063, 0.6026358, 0.5991582, 0.5982617, 0.5965938, 
    0.5982998, 0.5981609, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260328, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026052, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01193812, 0.01193812, 0.01193812, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01893771, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01193812, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 0.01193812, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 0.01193812, 
    0.01193812, 0.01193812 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.347731e-11, 3.362562e-11, 3.359671e-11, 3.371641e-11, 3.364996e-11, 
    3.37283e-11, 3.35072e-11, 3.363128e-11, 3.355201e-11, 3.349037e-11, 
    3.394868e-11, 3.372148e-11, 3.4185e-11, 3.40398e-11, 3.44046e-11, 
    3.416231e-11, 3.445347e-11, 3.439752e-11, 3.45658e-11, 3.451751e-11, 
    3.47329e-11, 3.458797e-11, 3.484461e-11, 3.469821e-11, 3.472106e-11, 
    3.458302e-11, 3.376742e-11, 3.392063e-11, 3.375828e-11, 3.378012e-11, 
    3.377029e-11, 3.365118e-11, 3.359121e-11, 3.346567e-11, 3.34884e-11, 
    3.358058e-11, 3.37897e-11, 3.371861e-11, 3.389765e-11, 3.389361e-11, 
    3.409313e-11, 3.400312e-11, 3.43389e-11, 3.424334e-11, 3.451949e-11, 
    3.444994e-11, 3.451615e-11, 3.449601e-11, 3.451632e-11, 3.441441e-11, 
    3.445799e-11, 3.436835e-11, 3.402038e-11, 3.412274e-11, 3.381747e-11, 
    3.363414e-11, 3.351249e-11, 3.342627e-11, 3.343838e-11, 3.346163e-11, 
    3.358105e-11, 3.369341e-11, 3.377912e-11, 3.383643e-11, 3.389293e-11, 
    3.406421e-11, 3.415489e-11, 3.435814e-11, 3.432142e-11, 3.438356e-11, 
    3.444299e-11, 3.454277e-11, 3.452632e-11, 3.457027e-11, 3.438174e-11, 
    3.450699e-11, 3.430023e-11, 3.435673e-11, 3.390865e-11, 3.373793e-11, 
    3.366542e-11, 3.360195e-11, 3.344773e-11, 3.355419e-11, 3.351217e-11, 
    3.3612e-11, 3.367549e-11, 3.364403e-11, 3.383796e-11, 3.376248e-11, 
    3.416022e-11, 3.398877e-11, 3.44361e-11, 3.432888e-11, 3.446169e-11, 
    3.439389e-11, 3.451002e-11, 3.440544e-11, 3.458657e-11, 3.462607e-11, 
    3.459901e-11, 3.470269e-11, 3.439943e-11, 3.451581e-11, 3.364335e-11, 
    3.364848e-11, 3.36723e-11, 3.356736e-11, 3.356094e-11, 3.346484e-11, 
    3.355025e-11, 3.358666e-11, 3.367908e-11, 3.373374e-11, 3.378572e-11, 
    3.390019e-11, 3.402807e-11, 3.420706e-11, 3.433578e-11, 3.442209e-11, 
    3.436912e-11, 3.441581e-11, 3.436353e-11, 3.433899e-11, 3.461117e-11, 
    3.445827e-11, 3.468767e-11, 3.467497e-11, 3.457104e-11, 3.467631e-11, 
    3.3652e-11, 3.362248e-11, 3.352017e-11, 3.360016e-11, 3.345432e-11, 
    3.353592e-11, 3.358281e-11, 3.376401e-11, 3.380381e-11, 3.384078e-11, 
    3.391376e-11, 3.400746e-11, 3.417206e-11, 3.431534e-11, 3.44463e-11, 
    3.443665e-11, 3.444001e-11, 3.446923e-11, 3.439672e-11, 3.448107e-11, 
    3.449519e-11, 3.445816e-11, 3.467317e-11, 3.46117e-11, 3.467457e-11, 
    3.463448e-11, 3.363202e-11, 3.368157e-11, 3.365472e-11, 3.370513e-11, 
    3.366954e-11, 3.382753e-11, 3.387488e-11, 3.409679e-11, 3.400562e-11, 
    3.415068e-11, 3.402028e-11, 3.404337e-11, 3.41553e-11, 3.402723e-11, 
    3.430735e-11, 3.411732e-11, 3.447033e-11, 3.42804e-11, 3.448217e-11, 
    3.444545e-11, 3.450611e-11, 3.456051e-11, 3.462888e-11, 3.475524e-11, 
    3.47259e-11, 3.483163e-11, 3.37555e-11, 3.381984e-11, 3.381416e-11, 
    3.388151e-11, 3.393134e-11, 3.403949e-11, 3.421304e-11, 3.414769e-11, 
    3.426755e-11, 3.429164e-11, 3.410941e-11, 3.422123e-11, 3.386259e-11, 
    3.392042e-11, 3.388594e-11, 3.376005e-11, 3.416245e-11, 3.395575e-11, 
    3.43375e-11, 3.422537e-11, 3.455265e-11, 3.438978e-11, 3.470976e-11, 
    3.484677e-11, 3.497575e-11, 3.51266e-11, 3.385495e-11, 3.381114e-11, 
    3.388946e-11, 3.399796e-11, 3.409861e-11, 3.423262e-11, 3.424629e-11, 
    3.427135e-11, 3.433637e-11, 3.439112e-11, 3.427921e-11, 3.440475e-11, 
    3.393381e-11, 3.418038e-11, 3.379414e-11, 3.391035e-11, 3.399108e-11, 
    3.395564e-11, 3.413978e-11, 3.418317e-11, 3.435975e-11, 3.426844e-11, 
    3.481284e-11, 3.457174e-11, 3.52415e-11, 3.505408e-11, 3.379581e-11, 
    3.385466e-11, 3.405977e-11, 3.396214e-11, 3.424147e-11, 3.431032e-11, 
    3.436622e-11, 3.443782e-11, 3.444548e-11, 3.448793e-11, 3.441832e-11, 
    3.448511e-11, 3.423253e-11, 3.434532e-11, 3.403593e-11, 3.411112e-11, 
    3.407649e-11, 3.403847e-11, 3.415563e-11, 3.428059e-11, 3.428322e-11, 
    3.432323e-11, 3.443622e-11, 3.424196e-11, 3.484385e-11, 3.447181e-11, 
    3.391887e-11, 3.403237e-11, 3.404856e-11, 3.400456e-11, 3.430332e-11, 
    3.419499e-11, 3.448689e-11, 3.440788e-11, 3.453722e-11, 3.447292e-11, 
    3.446339e-11, 3.438084e-11, 3.432939e-11, 3.419968e-11, 3.409412e-11, 
    3.401054e-11, 3.40299e-11, 3.412174e-11, 3.428813e-11, 3.444576e-11, 
    3.441116e-11, 3.452695e-11, 3.422049e-11, 3.434891e-11, 3.42992e-11, 
    3.442868e-11, 3.414581e-11, 3.438727e-11, 3.408411e-11, 3.411061e-11, 
    3.419274e-11, 3.435814e-11, 3.439469e-11, 3.44338e-11, 3.440959e-11, 
    3.429262e-11, 3.427341e-11, 3.419051e-11, 3.41676e-11, 3.410452e-11, 
    3.405223e-11, 3.409994e-11, 3.414998e-11, 3.42924e-11, 3.442077e-11, 
    3.456086e-11, 3.459515e-11, 3.475901e-11, 3.462555e-11, 3.484575e-11, 
    3.465845e-11, 3.498272e-11, 3.440117e-11, 3.465367e-11, 3.419648e-11, 
    3.424562e-11, 3.43346e-11, 3.453887e-11, 3.442849e-11, 3.455754e-11, 
    3.427264e-11, 3.412497e-11, 3.408675e-11, 3.401557e-11, 3.408832e-11, 
    3.40824e-11, 3.415206e-11, 3.412961e-11, 3.429702e-11, 3.420706e-11, 
    3.446269e-11, 3.455611e-11, 3.482015e-11, 3.498217e-11, 3.514729e-11, 
    3.522018e-11, 3.524237e-11, 3.525162e-11,
  1.906691e-11, 1.921087e-11, 1.918285e-11, 1.929919e-11, 1.923463e-11, 
    1.931085e-11, 1.909607e-11, 1.921659e-11, 1.913962e-11, 1.907986e-11, 
    1.952568e-11, 1.930439e-11, 1.975655e-11, 1.96147e-11, 1.997174e-11, 
    1.973444e-11, 2.001971e-11, 1.996488e-11, 2.013007e-11, 2.00827e-11, 
    2.029451e-11, 2.015195e-11, 2.040462e-11, 2.026043e-11, 2.028296e-11, 
    2.014726e-11, 1.934885e-11, 1.949808e-11, 1.934002e-11, 1.936127e-11, 
    1.935174e-11, 1.923596e-11, 1.91777e-11, 1.905593e-11, 1.907802e-11, 
    1.916747e-11, 1.937083e-11, 1.930171e-11, 1.947609e-11, 1.947215e-11, 
    1.966693e-11, 1.957902e-11, 1.990746e-11, 1.981392e-11, 2.008468e-11, 
    2.001646e-11, 2.008147e-11, 2.006175e-11, 2.008173e-11, 1.998171e-11, 
    2.002454e-11, 1.993661e-11, 1.959547e-11, 1.969551e-11, 1.93977e-11, 
    1.921941e-11, 1.910135e-11, 1.901773e-11, 1.902954e-11, 1.905207e-11, 
    1.916799e-11, 1.927723e-11, 1.936062e-11, 1.941648e-11, 1.947158e-11, 
    1.963868e-11, 1.972735e-11, 1.992639e-11, 1.989042e-11, 1.995138e-11, 
    2.000968e-11, 2.010769e-11, 2.009154e-11, 2.013477e-11, 1.994977e-11, 
    2.007265e-11, 1.986995e-11, 1.992531e-11, 1.948655e-11, 1.932035e-11, 
    1.924985e-11, 1.918824e-11, 1.903863e-11, 1.91419e-11, 1.910116e-11, 
    1.919813e-11, 1.925984e-11, 1.922931e-11, 1.941801e-11, 1.934457e-11, 
    1.973261e-11, 1.956513e-11, 2.000287e-11, 1.98978e-11, 2.002809e-11, 
    1.996157e-11, 2.007559e-11, 1.997296e-11, 2.015086e-11, 2.018967e-11, 
    2.016315e-11, 2.026511e-11, 1.996728e-11, 2.008147e-11, 1.922845e-11, 
    1.923343e-11, 1.925663e-11, 1.915474e-11, 1.914851e-11, 1.905533e-11, 
    1.913823e-11, 1.917358e-11, 1.926342e-11, 1.931663e-11, 1.936726e-11, 
    1.947876e-11, 1.960355e-11, 1.977855e-11, 1.990461e-11, 1.998928e-11, 
    1.993735e-11, 1.998319e-11, 1.993194e-11, 1.990794e-11, 2.017513e-11, 
    2.002494e-11, 2.025043e-11, 2.023793e-11, 2.013579e-11, 2.023934e-11, 
    1.923693e-11, 1.920829e-11, 1.910897e-11, 1.918668e-11, 1.904519e-11, 
    1.912434e-11, 1.91699e-11, 1.93461e-11, 1.938489e-11, 1.942089e-11, 
    1.949205e-11, 1.958352e-11, 1.974434e-11, 1.988466e-11, 2.001307e-11, 
    2.000365e-11, 2.000697e-11, 2.003569e-11, 1.996457e-11, 2.004737e-11, 
    2.006128e-11, 2.002492e-11, 2.023626e-11, 2.01758e-11, 2.023767e-11, 
    2.01983e-11, 1.92176e-11, 1.92658e-11, 1.923975e-11, 1.928875e-11, 
    1.925422e-11, 1.940794e-11, 1.945411e-11, 1.967071e-11, 1.958171e-11, 
    1.972342e-11, 1.959609e-11, 1.961863e-11, 1.972804e-11, 1.960297e-11, 
    1.987691e-11, 1.969103e-11, 2.003681e-11, 1.985064e-11, 2.004849e-11, 
    2.001251e-11, 2.00721e-11, 2.012551e-11, 2.019278e-11, 2.031712e-11, 
    2.02883e-11, 2.039244e-11, 1.933776e-11, 1.940044e-11, 1.939492e-11, 
    1.946059e-11, 1.95092e-11, 1.961473e-11, 1.978442e-11, 1.972055e-11, 
    1.983786e-11, 1.986144e-11, 1.968324e-11, 1.979258e-11, 1.944243e-11, 
    1.949884e-11, 1.946525e-11, 1.93427e-11, 1.973526e-11, 1.953343e-11, 
    1.990669e-11, 1.979693e-11, 2.011789e-11, 1.995803e-11, 2.027245e-11, 
    2.040738e-11, 2.053468e-11, 2.068377e-11, 1.943468e-11, 1.939205e-11, 
    1.94684e-11, 1.957421e-11, 1.967257e-11, 1.980362e-11, 1.981705e-11, 
    1.984164e-11, 1.990538e-11, 1.995904e-11, 1.984941e-11, 1.997249e-11, 
    1.951193e-11, 1.975281e-11, 1.937594e-11, 1.948914e-11, 1.956797e-11, 
    1.953338e-11, 1.971325e-11, 1.975573e-11, 1.992869e-11, 1.983922e-11, 
    2.037405e-11, 2.01368e-11, 2.079755e-11, 2.061214e-11, 1.937717e-11, 
    1.943453e-11, 1.963466e-11, 1.953935e-11, 1.981238e-11, 1.98798e-11, 
    1.993466e-11, 2.000487e-11, 2.001246e-11, 2.00541e-11, 1.998587e-11, 
    2.005141e-11, 1.98039e-11, 1.991437e-11, 1.961175e-11, 1.968525e-11, 
    1.965143e-11, 1.961435e-11, 1.972887e-11, 1.985113e-11, 1.985375e-11, 
    1.989301e-11, 2.000379e-11, 1.981349e-11, 2.040473e-11, 2.003885e-11, 
    1.949716e-11, 1.960795e-11, 1.96238e-11, 1.958084e-11, 1.987303e-11, 
    1.976698e-11, 2.005309e-11, 1.997562e-11, 2.010261e-11, 2.003947e-11, 
    2.003018e-11, 1.994921e-11, 1.989885e-11, 1.977184e-11, 1.966871e-11, 
    1.958707e-11, 1.960604e-11, 1.969576e-11, 1.985862e-11, 2.001314e-11, 
    1.997925e-11, 2.009295e-11, 1.979254e-11, 1.99183e-11, 1.986966e-11, 
    1.999659e-11, 1.971885e-11, 1.995525e-11, 1.965858e-11, 1.968453e-11, 
    1.976488e-11, 1.992684e-11, 1.996274e-11, 2.00011e-11, 1.997743e-11, 
    1.986276e-11, 1.9844e-11, 1.976292e-11, 1.974055e-11, 1.967888e-11, 
    1.962787e-11, 1.967448e-11, 1.972346e-11, 1.986282e-11, 1.998869e-11, 
    2.012627e-11, 2.015999e-11, 2.032124e-11, 2.018994e-11, 2.040677e-11, 
    2.022236e-11, 2.054197e-11, 1.996899e-11, 2.021695e-11, 1.976854e-11, 
    1.981667e-11, 1.990384e-11, 2.010429e-11, 1.999599e-11, 2.012267e-11, 
    1.984327e-11, 1.969885e-11, 1.966156e-11, 1.959203e-11, 1.966315e-11, 
    1.965736e-11, 1.972549e-11, 1.970359e-11, 1.986745e-11, 1.977937e-11, 
    2.002995e-11, 2.012167e-11, 2.038152e-11, 2.054139e-11, 2.070458e-11, 
    2.077677e-11, 2.079876e-11, 2.080795e-11,
  1.783523e-11, 1.799288e-11, 1.796219e-11, 1.808968e-11, 1.801891e-11, 
    1.810246e-11, 1.786714e-11, 1.799915e-11, 1.791483e-11, 1.78494e-11, 
    1.833818e-11, 1.809538e-11, 1.859185e-11, 1.843594e-11, 1.882863e-11, 
    1.856754e-11, 1.888147e-11, 1.882109e-11, 1.900307e-11, 1.895086e-11, 
    1.918441e-11, 1.902719e-11, 1.930595e-11, 1.914682e-11, 1.917167e-11, 
    1.902201e-11, 1.814414e-11, 1.830787e-11, 1.813445e-11, 1.815776e-11, 
    1.81473e-11, 1.802037e-11, 1.795655e-11, 1.78232e-11, 1.784738e-11, 
    1.794533e-11, 1.816824e-11, 1.809245e-11, 1.828374e-11, 1.827941e-11, 
    1.849333e-11, 1.839675e-11, 1.875787e-11, 1.865494e-11, 1.895304e-11, 
    1.887788e-11, 1.894951e-11, 1.892778e-11, 1.894979e-11, 1.883962e-11, 
    1.888679e-11, 1.878996e-11, 1.841482e-11, 1.852474e-11, 1.819771e-11, 
    1.800225e-11, 1.787292e-11, 1.778139e-11, 1.779432e-11, 1.781898e-11, 
    1.794591e-11, 1.806561e-11, 1.815705e-11, 1.821832e-11, 1.827878e-11, 
    1.846229e-11, 1.855974e-11, 1.877871e-11, 1.873912e-11, 1.880622e-11, 
    1.887041e-11, 1.89784e-11, 1.896061e-11, 1.900824e-11, 1.880445e-11, 
    1.893979e-11, 1.871659e-11, 1.877752e-11, 1.829522e-11, 1.811288e-11, 
    1.80356e-11, 1.796809e-11, 1.780426e-11, 1.791733e-11, 1.787272e-11, 
    1.797892e-11, 1.804655e-11, 1.801309e-11, 1.822e-11, 1.813944e-11, 
    1.856553e-11, 1.838149e-11, 1.886292e-11, 1.874724e-11, 1.889069e-11, 
    1.881744e-11, 1.894303e-11, 1.882998e-11, 1.902598e-11, 1.906877e-11, 
    1.903953e-11, 1.915198e-11, 1.882372e-11, 1.89495e-11, 1.801215e-11, 
    1.80176e-11, 1.804303e-11, 1.793139e-11, 1.792457e-11, 1.782254e-11, 
    1.791331e-11, 1.795203e-11, 1.805047e-11, 1.81088e-11, 1.816433e-11, 
    1.828666e-11, 1.842369e-11, 1.861603e-11, 1.875473e-11, 1.884795e-11, 
    1.879077e-11, 1.884125e-11, 1.878482e-11, 1.87584e-11, 1.905274e-11, 
    1.888723e-11, 1.913579e-11, 1.9122e-11, 1.900937e-11, 1.912355e-11, 
    1.802144e-11, 1.799005e-11, 1.788127e-11, 1.796638e-11, 1.781145e-11, 
    1.78981e-11, 1.7948e-11, 1.814112e-11, 1.818367e-11, 1.822316e-11, 
    1.830125e-11, 1.840169e-11, 1.857843e-11, 1.873278e-11, 1.887415e-11, 
    1.886378e-11, 1.886743e-11, 1.889907e-11, 1.882074e-11, 1.891194e-11, 
    1.892726e-11, 1.888721e-11, 1.912015e-11, 1.905348e-11, 1.91217e-11, 
    1.907828e-11, 1.800025e-11, 1.805308e-11, 1.802453e-11, 1.807824e-11, 
    1.804039e-11, 1.820895e-11, 1.825961e-11, 1.849748e-11, 1.839971e-11, 
    1.855542e-11, 1.84155e-11, 1.844026e-11, 1.85605e-11, 1.842305e-11, 
    1.872425e-11, 1.851982e-11, 1.89003e-11, 1.869534e-11, 1.891317e-11, 
    1.887354e-11, 1.893918e-11, 1.899804e-11, 1.907221e-11, 1.920936e-11, 
    1.917757e-11, 1.929251e-11, 1.813197e-11, 1.820072e-11, 1.819466e-11, 
    1.826672e-11, 1.832008e-11, 1.843598e-11, 1.862249e-11, 1.855226e-11, 
    1.868128e-11, 1.870723e-11, 1.851125e-11, 1.863147e-11, 1.824679e-11, 
    1.830871e-11, 1.827184e-11, 1.813739e-11, 1.856843e-11, 1.834669e-11, 
    1.875703e-11, 1.863626e-11, 1.898964e-11, 1.881355e-11, 1.916007e-11, 
    1.9309e-11, 1.944961e-11, 1.961445e-11, 1.823829e-11, 1.819152e-11, 
    1.82753e-11, 1.839146e-11, 1.849953e-11, 1.864361e-11, 1.865838e-11, 
    1.868543e-11, 1.875558e-11, 1.881465e-11, 1.869399e-11, 1.882947e-11, 
    1.832308e-11, 1.858773e-11, 1.817385e-11, 1.829806e-11, 1.838461e-11, 
    1.834663e-11, 1.854424e-11, 1.859095e-11, 1.878124e-11, 1.868277e-11, 
    1.927219e-11, 1.901048e-11, 1.974035e-11, 1.953524e-11, 1.817519e-11, 
    1.823813e-11, 1.845787e-11, 1.835318e-11, 1.865325e-11, 1.872742e-11, 
    1.878781e-11, 1.886512e-11, 1.887347e-11, 1.891935e-11, 1.88442e-11, 
    1.891638e-11, 1.864392e-11, 1.876547e-11, 1.84327e-11, 1.851347e-11, 
    1.847629e-11, 1.843555e-11, 1.856141e-11, 1.869588e-11, 1.869877e-11, 
    1.874197e-11, 1.886394e-11, 1.865447e-11, 1.930607e-11, 1.890255e-11, 
    1.830686e-11, 1.842852e-11, 1.844594e-11, 1.839875e-11, 1.871998e-11, 
    1.860332e-11, 1.891823e-11, 1.883291e-11, 1.89728e-11, 1.890323e-11, 
    1.8893e-11, 1.880383e-11, 1.87484e-11, 1.860866e-11, 1.849528e-11, 
    1.840559e-11, 1.842643e-11, 1.852501e-11, 1.870412e-11, 1.887423e-11, 
    1.883691e-11, 1.896215e-11, 1.863142e-11, 1.876981e-11, 1.871627e-11, 
    1.8856e-11, 1.85504e-11, 1.881049e-11, 1.848416e-11, 1.851267e-11, 
    1.8601e-11, 1.87792e-11, 1.881873e-11, 1.886097e-11, 1.88349e-11, 
    1.870868e-11, 1.868804e-11, 1.859886e-11, 1.857426e-11, 1.850647e-11, 
    1.845041e-11, 1.850162e-11, 1.855546e-11, 1.870874e-11, 1.884731e-11, 
    1.899888e-11, 1.903605e-11, 1.921391e-11, 1.906907e-11, 1.930833e-11, 
    1.910482e-11, 1.945767e-11, 1.882561e-11, 1.909886e-11, 1.860503e-11, 
    1.865797e-11, 1.875388e-11, 1.897466e-11, 1.885534e-11, 1.899491e-11, 
    1.868723e-11, 1.852841e-11, 1.848742e-11, 1.841103e-11, 1.848917e-11, 
    1.848281e-11, 1.85577e-11, 1.853362e-11, 1.871383e-11, 1.861694e-11, 
    1.889274e-11, 1.899381e-11, 1.928044e-11, 1.945703e-11, 1.963747e-11, 
    1.971735e-11, 1.974168e-11, 1.975186e-11,
  1.829495e-11, 1.846857e-11, 1.843476e-11, 1.857525e-11, 1.849725e-11, 
    1.858933e-11, 1.833008e-11, 1.847548e-11, 1.83826e-11, 1.831054e-11, 
    1.884935e-11, 1.858153e-11, 1.912948e-11, 1.895725e-11, 1.939132e-11, 
    1.910263e-11, 1.944978e-11, 1.938296e-11, 1.95844e-11, 1.952659e-11, 
    1.978533e-11, 1.961111e-11, 1.99201e-11, 1.974366e-11, 1.977121e-11, 
    1.960538e-11, 1.863527e-11, 1.881591e-11, 1.86246e-11, 1.86503e-11, 
    1.863876e-11, 1.849886e-11, 1.842855e-11, 1.828171e-11, 1.830832e-11, 
    1.841619e-11, 1.866186e-11, 1.857829e-11, 1.878925e-11, 1.878447e-11, 
    1.902064e-11, 1.891398e-11, 1.931303e-11, 1.919921e-11, 1.9529e-11, 
    1.944581e-11, 1.952509e-11, 1.950103e-11, 1.952541e-11, 1.940346e-11, 
    1.945566e-11, 1.934853e-11, 1.893393e-11, 1.905534e-11, 1.869436e-11, 
    1.84789e-11, 1.833645e-11, 1.823568e-11, 1.824991e-11, 1.827705e-11, 
    1.841683e-11, 1.85487e-11, 1.864951e-11, 1.871709e-11, 1.878378e-11, 
    1.898637e-11, 1.909401e-11, 1.933609e-11, 1.929229e-11, 1.936651e-11, 
    1.943754e-11, 1.955708e-11, 1.953738e-11, 1.959013e-11, 1.936455e-11, 
    1.951433e-11, 1.926737e-11, 1.933477e-11, 1.880194e-11, 1.860082e-11, 
    1.851565e-11, 1.844125e-11, 1.826086e-11, 1.838535e-11, 1.833622e-11, 
    1.845319e-11, 1.85277e-11, 1.849083e-11, 1.871893e-11, 1.863009e-11, 
    1.91004e-11, 1.889714e-11, 1.942925e-11, 1.930128e-11, 1.945999e-11, 
    1.937892e-11, 1.951792e-11, 1.93928e-11, 1.960978e-11, 1.965718e-11, 
    1.962478e-11, 1.974937e-11, 1.938588e-11, 1.952509e-11, 1.84898e-11, 
    1.849581e-11, 1.852382e-11, 1.840083e-11, 1.839332e-11, 1.828098e-11, 
    1.838092e-11, 1.842356e-11, 1.853202e-11, 1.859632e-11, 1.865754e-11, 
    1.879248e-11, 1.894374e-11, 1.915621e-11, 1.930956e-11, 1.941268e-11, 
    1.934942e-11, 1.940527e-11, 1.934284e-11, 1.931361e-11, 1.963942e-11, 
    1.945615e-11, 1.973143e-11, 1.971615e-11, 1.959139e-11, 1.971787e-11, 
    1.850003e-11, 1.846545e-11, 1.834564e-11, 1.843937e-11, 1.826876e-11, 
    1.836417e-11, 1.841913e-11, 1.863195e-11, 1.867886e-11, 1.872242e-11, 
    1.880858e-11, 1.891943e-11, 1.911465e-11, 1.928528e-11, 1.944168e-11, 
    1.94302e-11, 1.943424e-11, 1.946926e-11, 1.938258e-11, 1.948351e-11, 
    1.950047e-11, 1.945613e-11, 1.97141e-11, 1.964024e-11, 1.971582e-11, 
    1.966771e-11, 1.847669e-11, 1.85349e-11, 1.850343e-11, 1.856263e-11, 
    1.852092e-11, 1.870675e-11, 1.876264e-11, 1.902522e-11, 1.891725e-11, 
    1.908923e-11, 1.893468e-11, 1.896202e-11, 1.909486e-11, 1.894302e-11, 
    1.927586e-11, 1.90499e-11, 1.947062e-11, 1.924389e-11, 1.948487e-11, 
    1.9441e-11, 1.951365e-11, 1.957884e-11, 1.966098e-11, 1.981298e-11, 
    1.977774e-11, 1.990517e-11, 1.862186e-11, 1.869767e-11, 1.869099e-11, 
    1.877047e-11, 1.882936e-11, 1.895729e-11, 1.916335e-11, 1.908574e-11, 
    1.922833e-11, 1.925702e-11, 1.904043e-11, 1.917327e-11, 1.874849e-11, 
    1.881681e-11, 1.877612e-11, 1.862783e-11, 1.910361e-11, 1.885873e-11, 
    1.93121e-11, 1.917856e-11, 1.956954e-11, 1.937463e-11, 1.975835e-11, 
    1.992348e-11, 2.007949e-11, 2.026255e-11, 1.873911e-11, 1.868752e-11, 
    1.877993e-11, 1.890815e-11, 1.902748e-11, 1.918669e-11, 1.920302e-11, 
    1.923292e-11, 1.93105e-11, 1.937584e-11, 1.924239e-11, 1.939223e-11, 
    1.883268e-11, 1.912494e-11, 1.866804e-11, 1.880507e-11, 1.890058e-11, 
    1.885865e-11, 1.907688e-11, 1.912848e-11, 1.933888e-11, 1.922998e-11, 
    1.988266e-11, 1.959262e-11, 2.040246e-11, 2.017457e-11, 1.866952e-11, 
    1.873893e-11, 1.898147e-11, 1.886589e-11, 1.919734e-11, 1.927935e-11, 
    1.934614e-11, 1.943169e-11, 1.944093e-11, 1.949171e-11, 1.940853e-11, 
    1.948842e-11, 1.918703e-11, 1.932144e-11, 1.895367e-11, 1.904287e-11, 
    1.900181e-11, 1.895682e-11, 1.909584e-11, 1.924449e-11, 1.924766e-11, 
    1.929545e-11, 1.943041e-11, 1.919869e-11, 1.992025e-11, 1.947314e-11, 
    1.881476e-11, 1.894907e-11, 1.896829e-11, 1.891618e-11, 1.927112e-11, 
    1.914215e-11, 1.949047e-11, 1.939604e-11, 1.955088e-11, 1.947386e-11, 
    1.946254e-11, 1.936386e-11, 1.930255e-11, 1.914806e-11, 1.902279e-11, 
    1.892374e-11, 1.894675e-11, 1.905563e-11, 1.92536e-11, 1.944177e-11, 
    1.940047e-11, 1.953909e-11, 1.917322e-11, 1.932623e-11, 1.926702e-11, 
    1.942159e-11, 1.908368e-11, 1.937126e-11, 1.90105e-11, 1.9042e-11, 
    1.91396e-11, 1.933663e-11, 1.938035e-11, 1.942709e-11, 1.939825e-11, 
    1.925863e-11, 1.92358e-11, 1.913722e-11, 1.911005e-11, 1.903514e-11, 
    1.897323e-11, 1.902979e-11, 1.908928e-11, 1.925869e-11, 1.941198e-11, 
    1.957976e-11, 1.962093e-11, 1.981805e-11, 1.965752e-11, 1.992276e-11, 
    1.969715e-11, 2.008846e-11, 1.938798e-11, 1.969053e-11, 1.914404e-11, 
    1.920256e-11, 1.930863e-11, 1.955295e-11, 1.942086e-11, 1.957538e-11, 
    1.923491e-11, 1.905939e-11, 1.901411e-11, 1.892975e-11, 1.901604e-11, 
    1.900901e-11, 1.909174e-11, 1.906513e-11, 1.926433e-11, 1.915721e-11, 
    1.946226e-11, 1.957415e-11, 1.98918e-11, 2.008773e-11, 2.028811e-11, 
    2.037688e-11, 2.040394e-11, 2.041525e-11,
  1.973495e-11, 1.991889e-11, 1.988306e-11, 2.003198e-11, 1.994929e-11, 
    2.004692e-11, 1.977216e-11, 1.992622e-11, 1.982779e-11, 1.975146e-11, 
    2.032282e-11, 2.003864e-11, 2.062039e-11, 2.043737e-11, 2.08989e-11, 
    2.059186e-11, 2.096113e-11, 2.088999e-11, 2.110448e-11, 2.10429e-11, 
    2.131865e-11, 2.113293e-11, 2.146239e-11, 2.127421e-11, 2.130359e-11, 
    2.112682e-11, 2.009563e-11, 2.028732e-11, 2.008431e-11, 2.011157e-11, 
    2.009933e-11, 1.9951e-11, 1.987649e-11, 1.972093e-11, 1.974911e-11, 
    1.986339e-11, 2.012384e-11, 2.00352e-11, 2.025899e-11, 2.025392e-11, 
    2.050471e-11, 2.039141e-11, 2.081558e-11, 2.069451e-11, 2.104547e-11, 
    2.095689e-11, 2.104131e-11, 2.101569e-11, 2.104164e-11, 2.091181e-11, 
    2.096738e-11, 2.085334e-11, 2.041261e-11, 2.054158e-11, 2.015831e-11, 
    1.992986e-11, 1.977891e-11, 1.96722e-11, 1.968726e-11, 1.9716e-11, 
    1.986406e-11, 2.000383e-11, 2.011073e-11, 2.018241e-11, 2.025319e-11, 
    2.046832e-11, 2.058269e-11, 2.084012e-11, 2.079351e-11, 2.087249e-11, 
    2.094809e-11, 2.107538e-11, 2.105439e-11, 2.111059e-11, 2.08704e-11, 
    2.102985e-11, 2.076699e-11, 2.08387e-11, 2.02725e-11, 2.005909e-11, 
    1.996881e-11, 1.988994e-11, 1.969885e-11, 1.983071e-11, 1.977867e-11, 
    1.990259e-11, 1.998156e-11, 1.994248e-11, 2.018438e-11, 2.009014e-11, 
    2.058948e-11, 2.037353e-11, 2.093926e-11, 2.080307e-11, 2.097198e-11, 
    2.088569e-11, 2.103367e-11, 2.090046e-11, 2.113152e-11, 2.118203e-11, 
    2.11475e-11, 2.128029e-11, 2.089309e-11, 2.104131e-11, 1.994139e-11, 
    1.994776e-11, 1.997745e-11, 1.984712e-11, 1.983915e-11, 1.972015e-11, 
    1.982602e-11, 1.98712e-11, 1.998614e-11, 2.005432e-11, 2.011924e-11, 
    2.026242e-11, 2.042302e-11, 2.06488e-11, 2.081189e-11, 2.092162e-11, 
    2.085429e-11, 2.091373e-11, 2.084729e-11, 2.081619e-11, 2.11631e-11, 
    2.09679e-11, 2.126116e-11, 2.124487e-11, 2.111192e-11, 2.124671e-11, 
    1.995223e-11, 1.991558e-11, 1.978864e-11, 1.988794e-11, 1.970722e-11, 
    1.980827e-11, 1.986651e-11, 2.009211e-11, 2.014187e-11, 2.018808e-11, 
    2.027951e-11, 2.03972e-11, 2.060462e-11, 2.078606e-11, 2.095249e-11, 
    2.094027e-11, 2.094457e-11, 2.098185e-11, 2.088958e-11, 2.099702e-11, 
    2.101509e-11, 2.096787e-11, 2.124269e-11, 2.116396e-11, 2.124453e-11, 
    2.119324e-11, 1.992749e-11, 1.99892e-11, 1.995584e-11, 2.00186e-11, 
    1.997438e-11, 2.017147e-11, 2.023077e-11, 2.050959e-11, 2.039489e-11, 
    2.05776e-11, 2.04134e-11, 2.044244e-11, 2.05836e-11, 2.042225e-11, 
    2.077604e-11, 2.053582e-11, 2.09833e-11, 2.074205e-11, 2.099847e-11, 
    2.095177e-11, 2.102912e-11, 2.109855e-11, 2.118607e-11, 2.134813e-11, 
    2.131054e-11, 2.144647e-11, 2.00814e-11, 2.016183e-11, 2.015473e-11, 
    2.023907e-11, 2.030157e-11, 2.043741e-11, 2.065638e-11, 2.057388e-11, 
    2.072548e-11, 2.075599e-11, 2.052573e-11, 2.066694e-11, 2.021574e-11, 
    2.028826e-11, 2.024506e-11, 2.008774e-11, 2.059289e-11, 2.033275e-11, 
    2.081459e-11, 2.067255e-11, 2.108864e-11, 2.088113e-11, 2.128986e-11, 
    2.146602e-11, 2.163254e-11, 2.182814e-11, 2.020578e-11, 2.015105e-11, 
    2.024911e-11, 2.038524e-11, 2.051198e-11, 2.06812e-11, 2.069856e-11, 
    2.073037e-11, 2.081288e-11, 2.088241e-11, 2.074044e-11, 2.089985e-11, 
    2.030512e-11, 2.061555e-11, 2.013039e-11, 2.02758e-11, 2.037719e-11, 
    2.033267e-11, 2.056446e-11, 2.061932e-11, 2.084309e-11, 2.072723e-11, 
    2.142247e-11, 2.111324e-11, 2.197773e-11, 2.173411e-11, 2.013195e-11, 
    2.020559e-11, 2.046311e-11, 2.034035e-11, 2.069252e-11, 2.077975e-11, 
    2.08508e-11, 2.094185e-11, 2.095169e-11, 2.100576e-11, 2.09172e-11, 
    2.100225e-11, 2.068156e-11, 2.082452e-11, 2.043357e-11, 2.052833e-11, 
    2.04847e-11, 2.043691e-11, 2.058462e-11, 2.074267e-11, 2.074604e-11, 
    2.079687e-11, 2.094054e-11, 2.069396e-11, 2.14626e-11, 2.098602e-11, 
    2.028607e-11, 2.04287e-11, 2.04491e-11, 2.039375e-11, 2.077099e-11, 
    2.063385e-11, 2.100444e-11, 2.09039e-11, 2.106877e-11, 2.098675e-11, 
    2.09747e-11, 2.086966e-11, 2.080443e-11, 2.064013e-11, 2.0507e-11, 
    2.040177e-11, 2.042621e-11, 2.054189e-11, 2.075236e-11, 2.095259e-11, 
    2.090863e-11, 2.105621e-11, 2.066687e-11, 2.082963e-11, 2.076664e-11, 
    2.093111e-11, 2.057169e-11, 2.087757e-11, 2.049393e-11, 2.05274e-11, 
    2.063113e-11, 2.08407e-11, 2.088721e-11, 2.093696e-11, 2.090625e-11, 
    2.075771e-11, 2.073343e-11, 2.06286e-11, 2.059972e-11, 2.052011e-11, 
    2.045434e-11, 2.051443e-11, 2.057765e-11, 2.075777e-11, 2.092088e-11, 
    2.109954e-11, 2.114339e-11, 2.135355e-11, 2.11824e-11, 2.146528e-11, 
    2.122467e-11, 2.164215e-11, 2.089535e-11, 2.121759e-11, 2.063585e-11, 
    2.069807e-11, 2.08109e-11, 2.107099e-11, 2.093033e-11, 2.109488e-11, 
    2.073248e-11, 2.05459e-11, 2.049776e-11, 2.040816e-11, 2.049982e-11, 
    2.049235e-11, 2.058026e-11, 2.055198e-11, 2.076377e-11, 2.064985e-11, 
    2.09744e-11, 2.109357e-11, 2.14322e-11, 2.164136e-11, 2.185545e-11, 
    2.195037e-11, 2.19793e-11, 2.199141e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
