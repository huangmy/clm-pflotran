netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/20/14 16:23:17" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/20/14" ;

 time_written =
  "16:23:17" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.485607e-14, 4.497747e-14, 4.495389e-14, 4.505172e-14, 4.499748e-14, 
    4.506151e-14, 4.488071e-14, 4.498227e-14, 4.491746e-14, 4.486703e-14, 
    4.524128e-14, 4.505608e-14, 4.54335e-14, 4.53156e-14, 4.561158e-14, 
    4.541514e-14, 4.565116e-14, 4.560596e-14, 4.574206e-14, 4.570309e-14, 
    4.58769e-14, 4.576004e-14, 4.596696e-14, 4.584903e-14, 4.586747e-14, 
    4.575618e-14, 4.509342e-14, 4.521822e-14, 4.508601e-14, 4.510382e-14, 
    4.509583e-14, 4.499858e-14, 4.494952e-14, 4.484682e-14, 4.486548e-14, 
    4.494092e-14, 4.511182e-14, 4.505386e-14, 4.519997e-14, 4.519667e-14, 
    4.535908e-14, 4.528588e-14, 4.555852e-14, 4.548112e-14, 4.570472e-14, 
    4.564851e-14, 4.570207e-14, 4.568584e-14, 4.570228e-14, 4.561985e-14, 
    4.565517e-14, 4.558262e-14, 4.529958e-14, 4.538283e-14, 4.513434e-14, 
    4.498462e-14, 4.488516e-14, 4.481451e-14, 4.48245e-14, 4.484354e-14, 
    4.494136e-14, 4.50333e-14, 4.51033e-14, 4.51501e-14, 4.519619e-14, 
    4.53355e-14, 4.540926e-14, 4.557415e-14, 4.554444e-14, 4.559479e-14, 
    4.564292e-14, 4.572364e-14, 4.571036e-14, 4.57459e-14, 4.559349e-14, 
    4.569479e-14, 4.552753e-14, 4.557328e-14, 4.520858e-14, 4.506951e-14, 
    4.501023e-14, 4.495842e-14, 4.483218e-14, 4.491936e-14, 4.4885e-14, 
    4.496677e-14, 4.501868e-14, 4.499301e-14, 4.515138e-14, 4.508983e-14, 
    4.541363e-14, 4.527427e-14, 4.563731e-14, 4.555054e-14, 4.56581e-14, 
    4.560324e-14, 4.569722e-14, 4.561264e-14, 4.575914e-14, 4.579099e-14, 
    4.576922e-14, 4.585288e-14, 4.560794e-14, 4.570206e-14, 4.499229e-14, 
    4.499647e-14, 4.501599e-14, 4.493019e-14, 4.492494e-14, 4.48463e-14, 
    4.491629e-14, 4.494607e-14, 4.50217e-14, 4.506638e-14, 4.510885e-14, 
    4.520218e-14, 4.53063e-14, 4.545177e-14, 4.555617e-14, 4.56261e-14, 
    4.558323e-14, 4.562108e-14, 4.557876e-14, 4.555893e-14, 4.577905e-14, 
    4.565549e-14, 4.584085e-14, 4.583061e-14, 4.574674e-14, 4.583176e-14, 
    4.499941e-14, 4.497533e-14, 4.48916e-14, 4.495713e-14, 4.483773e-14, 
    4.490456e-14, 4.494296e-14, 4.509108e-14, 4.512364e-14, 4.515377e-14, 
    4.52133e-14, 4.528963e-14, 4.54234e-14, 4.553966e-14, 4.564573e-14, 
    4.563796e-14, 4.56407e-14, 4.566436e-14, 4.560571e-14, 4.567399e-14, 
    4.568543e-14, 4.565549e-14, 4.582924e-14, 4.577963e-14, 4.583039e-14, 
    4.57981e-14, 4.498316e-14, 4.50237e-14, 4.500179e-14, 4.504297e-14, 
    4.501395e-14, 4.51429e-14, 4.518154e-14, 4.536219e-14, 4.528812e-14, 
    4.540601e-14, 4.530011e-14, 4.531887e-14, 4.54098e-14, 4.530584e-14, 
    4.553325e-14, 4.537907e-14, 4.566528e-14, 4.551147e-14, 4.567491e-14, 
    4.564527e-14, 4.569436e-14, 4.57383e-14, 4.579357e-14, 4.589544e-14, 
    4.587187e-14, 4.595703e-14, 4.508411e-14, 4.513663e-14, 4.513204e-14, 
    4.5187e-14, 4.522762e-14, 4.531564e-14, 4.545666e-14, 4.540366e-14, 
    4.550097e-14, 4.552048e-14, 4.537265e-14, 4.546342e-14, 4.517179e-14, 
    4.521893e-14, 4.519088e-14, 4.508824e-14, 4.541584e-14, 4.524782e-14, 
    4.555789e-14, 4.546704e-14, 4.573203e-14, 4.560028e-14, 4.585888e-14, 
    4.596918e-14, 4.607301e-14, 4.619408e-14, 4.516532e-14, 4.512964e-14, 
    4.519354e-14, 4.528184e-14, 4.536377e-14, 4.547258e-14, 4.548372e-14, 
    4.550408e-14, 4.555682e-14, 4.560114e-14, 4.551049e-14, 4.561226e-14, 
    4.52298e-14, 4.543042e-14, 4.511612e-14, 4.521082e-14, 4.527664e-14, 
    4.52478e-14, 4.53976e-14, 4.543288e-14, 4.557605e-14, 4.550209e-14, 
    4.594194e-14, 4.574753e-14, 4.628626e-14, 4.613596e-14, 4.511717e-14, 
    4.516521e-14, 4.533221e-14, 4.525279e-14, 4.547985e-14, 4.553566e-14, 
    4.558101e-14, 4.563894e-14, 4.564522e-14, 4.567953e-14, 4.56233e-14, 
    4.567732e-14, 4.547281e-14, 4.556424e-14, 4.531317e-14, 4.537431e-14, 
    4.53462e-14, 4.531533e-14, 4.541057e-14, 4.551191e-14, 4.551412e-14, 
    4.554656e-14, 4.563793e-14, 4.548077e-14, 4.596693e-14, 4.566685e-14, 
    4.521757e-14, 4.530994e-14, 4.532318e-14, 4.528741e-14, 4.553007e-14, 
    4.54422e-14, 4.56787e-14, 4.561483e-14, 4.571947e-14, 4.566748e-14, 
    4.565983e-14, 4.559303e-14, 4.555141e-14, 4.544622e-14, 4.536055e-14, 
    4.52926e-14, 4.530841e-14, 4.538304e-14, 4.551812e-14, 4.564577e-14, 
    4.56178e-14, 4.571152e-14, 4.54634e-14, 4.556747e-14, 4.552726e-14, 
    4.563213e-14, 4.540224e-14, 4.55979e-14, 4.535215e-14, 4.537373e-14, 
    4.544045e-14, 4.55745e-14, 4.56042e-14, 4.563583e-14, 4.561633e-14, 
    4.552156e-14, 4.550604e-14, 4.543884e-14, 4.542026e-14, 4.536904e-14, 
    4.532659e-14, 4.536536e-14, 4.540605e-14, 4.552161e-14, 4.56256e-14, 
    4.573892e-14, 4.576664e-14, 4.589875e-14, 4.579116e-14, 4.596859e-14, 
    4.581767e-14, 4.607883e-14, 4.560929e-14, 4.581332e-14, 4.54435e-14, 
    4.548341e-14, 4.55555e-14, 4.57208e-14, 4.563163e-14, 4.573593e-14, 
    4.550543e-14, 4.538559e-14, 4.535462e-14, 4.529672e-14, 4.535594e-14, 
    4.535113e-14, 4.540777e-14, 4.538958e-14, 4.552545e-14, 4.545249e-14, 
    4.565962e-14, 4.573512e-14, 4.59481e-14, 4.607843e-14, 4.621101e-14, 
    4.626946e-14, 4.628725e-14, 4.629468e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.859499e-14, -1.861845e-14, -1.861388e-14, -1.863279e-14, -1.862229e-14, 
    -1.863468e-14, -1.859973e-14, -1.861939e-14, -1.860684e-14, 
    -1.859708e-14, -1.866941e-14, -1.863363e-14, -1.870627e-14, 
    -1.868359e-14, -1.874048e-14, -1.870277e-14, -1.874807e-14, 
    -1.873936e-14, -1.876545e-14, -1.875799e-14, -1.879134e-14, -1.87689e-14, 
    -1.880853e-14, -1.878597e-14, -1.878952e-14, -1.876816e-14, 
    -1.864081e-14, -1.866497e-14, -1.863938e-14, -1.864283e-14, 
    -1.864128e-14, -1.862252e-14, -1.861308e-14, -1.859317e-14, 
    -1.859678e-14, -1.861139e-14, -1.864438e-14, -1.863317e-14, 
    -1.866132e-14, -1.866069e-14, -1.869194e-14, -1.867787e-14, 
    -1.873025e-14, -1.871536e-14, -1.87583e-14, -1.874752e-14, -1.87578e-14, 
    -1.875468e-14, -1.875784e-14, -1.874203e-14, -1.874881e-14, 
    -1.873487e-14, -1.868051e-14, -1.869652e-14, -1.864871e-14, 
    -1.861988e-14, -1.86006e-14, -1.858692e-14, -1.858886e-14, -1.859255e-14, 
    -1.861148e-14, -1.86292e-14, -1.86427e-14, -1.865172e-14, -1.86606e-14, 
    -1.868749e-14, -1.870162e-14, -1.873328e-14, -1.872754e-14, 
    -1.873724e-14, -1.874645e-14, -1.876194e-14, -1.875938e-14, 
    -1.876621e-14, -1.873696e-14, -1.875642e-14, -1.872427e-14, 
    -1.873308e-14, -1.866313e-14, -1.863619e-14, -1.862482e-14, 
    -1.861477e-14, -1.859035e-14, -1.860722e-14, -1.860058e-14, 
    -1.861636e-14, -1.862638e-14, -1.862142e-14, -1.865197e-14, 
    -1.864011e-14, -1.870246e-14, -1.867566e-14, -1.874538e-14, 
    -1.872871e-14, -1.874936e-14, -1.873883e-14, -1.875688e-14, 
    -1.874063e-14, -1.876874e-14, -1.877486e-14, -1.877068e-14, 
    -1.878668e-14, -1.873973e-14, -1.875781e-14, -1.862129e-14, -1.86221e-14, 
    -1.862586e-14, -1.860932e-14, -1.86083e-14, -1.859308e-14, -1.860661e-14, 
    -1.861238e-14, -1.862696e-14, -1.863559e-14, -1.864378e-14, 
    -1.866176e-14, -1.868182e-14, -1.870976e-14, -1.87298e-14, -1.874321e-14, 
    -1.873498e-14, -1.874225e-14, -1.873413e-14, -1.873031e-14, 
    -1.877257e-14, -1.874888e-14, -1.878438e-14, -1.878242e-14, 
    -1.876637e-14, -1.878264e-14, -1.862266e-14, -1.8618e-14, -1.860184e-14, 
    -1.861449e-14, -1.859141e-14, -1.860436e-14, -1.861179e-14, 
    -1.864038e-14, -1.864662e-14, -1.865244e-14, -1.86639e-14, -1.867859e-14, 
    -1.870431e-14, -1.872664e-14, -1.874698e-14, -1.874549e-14, 
    -1.874601e-14, -1.875057e-14, -1.873931e-14, -1.875241e-14, 
    -1.875462e-14, -1.874886e-14, -1.878215e-14, -1.877265e-14, 
    -1.878238e-14, -1.877619e-14, -1.861952e-14, -1.862735e-14, 
    -1.862312e-14, -1.863108e-14, -1.862548e-14, -1.865038e-14, 
    -1.865783e-14, -1.869258e-14, -1.86783e-14, -1.870098e-14, -1.86806e-14, 
    -1.868422e-14, -1.870176e-14, -1.86817e-14, -1.872543e-14, -1.869584e-14, 
    -1.875074e-14, -1.872127e-14, -1.875259e-14, -1.874689e-14, 
    -1.875631e-14, -1.876475e-14, -1.877533e-14, -1.879485e-14, 
    -1.879033e-14, -1.880661e-14, -1.863901e-14, -1.864915e-14, 
    -1.864824e-14, -1.865883e-14, -1.866666e-14, -1.868358e-14, 
    -1.871068e-14, -1.870049e-14, -1.871917e-14, -1.872293e-14, 
    -1.869453e-14, -1.871199e-14, -1.865592e-14, -1.866503e-14, 
    -1.865959e-14, -1.863982e-14, -1.870287e-14, -1.867058e-14, 
    -1.873013e-14, -1.871266e-14, -1.876355e-14, -1.87383e-14, -1.878784e-14, 
    -1.880899e-14, -1.882875e-14, -1.885189e-14, -1.865466e-14, 
    -1.864778e-14, -1.866009e-14, -1.867713e-14, -1.869284e-14, 
    -1.871373e-14, -1.871586e-14, -1.871978e-14, -1.872991e-14, 
    -1.873843e-14, -1.872104e-14, -1.874056e-14, -1.866718e-14, 
    -1.870566e-14, -1.864519e-14, -1.866347e-14, -1.867611e-14, 
    -1.867055e-14, -1.869932e-14, -1.87061e-14, -1.873364e-14, -1.871938e-14, 
    -1.88038e-14, -1.876656e-14, -1.88694e-14, -1.88408e-14, -1.864537e-14, 
    -1.865463e-14, -1.86868e-14, -1.86715e-14, -1.871511e-14, -1.872585e-14, 
    -1.873455e-14, -1.87457e-14, -1.874689e-14, -1.875348e-14, -1.874268e-14, 
    -1.875305e-14, -1.871378e-14, -1.873134e-14, -1.86831e-14, -1.869487e-14, 
    -1.868945e-14, -1.868352e-14, -1.870181e-14, -1.872132e-14, -1.87217e-14, 
    -1.872797e-14, -1.874565e-14, -1.871529e-14, -1.880866e-14, 
    -1.875118e-14, -1.866471e-14, -1.868254e-14, -1.868504e-14, 
    -1.867815e-14, -1.872478e-14, -1.87079e-14, -1.875331e-14, -1.874105e-14, 
    -1.876113e-14, -1.875116e-14, -1.874969e-14, -1.873687e-14, 
    -1.872888e-14, -1.870868e-14, -1.869223e-14, -1.867914e-14, 
    -1.868218e-14, -1.869655e-14, -1.87225e-14, -1.874701e-14, -1.874165e-14, 
    -1.87596e-14, -1.871196e-14, -1.873198e-14, -1.872426e-14, -1.874438e-14, 
    -1.870023e-14, -1.873794e-14, -1.869059e-14, -1.869474e-14, 
    -1.870756e-14, -1.873337e-14, -1.873901e-14, -1.874511e-14, 
    -1.874134e-14, -1.872316e-14, -1.872016e-14, -1.870724e-14, 
    -1.870369e-14, -1.869383e-14, -1.868568e-14, -1.869314e-14, 
    -1.870097e-14, -1.872315e-14, -1.874314e-14, -1.876487e-14, 
    -1.877017e-14, -1.879556e-14, -1.877494e-14, -1.880898e-14, 
    -1.878012e-14, -1.882998e-14, -1.874007e-14, -1.87792e-14, -1.870813e-14, 
    -1.871579e-14, -1.87297e-14, -1.876144e-14, -1.874428e-14, -1.876433e-14, 
    -1.872004e-14, -1.869706e-14, -1.869107e-14, -1.867995e-14, 
    -1.869132e-14, -1.86904e-14, -1.870127e-14, -1.869778e-14, -1.872389e-14, 
    -1.870986e-14, -1.874967e-14, -1.876416e-14, -1.880492e-14, 
    -1.882983e-14, -1.885506e-14, -1.886619e-14, -1.886957e-14, -1.887098e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.52139e-11, 1.520956e-11, 1.521047e-11, 1.520648e-11, 1.520877e-11, 
    1.520605e-11, 1.521309e-11, 1.520937e-11, 1.521181e-11, 1.521354e-11, 
    1.519693e-11, 1.520629e-11, 1.518437e-11, 1.519247e-11, 1.508232e-11, 
    1.518571e-11, 1.508282e-11, 1.508223e-11, 1.508284e-11, 1.508303e-11, 
    1.507981e-11, 1.508265e-11, 1.507563e-11, 1.508075e-11, 1.508015e-11, 
    1.50827e-11, 1.52046e-11, 1.519823e-11, 1.520494e-11, 1.520411e-11, 
    1.520449e-11, 1.520872e-11, 1.521063e-11, 1.52142e-11, 1.52136e-11, 
    1.521095e-11, 1.520373e-11, 1.520639e-11, 1.519925e-11, 1.519943e-11, 
    1.518963e-11, 1.519432e-11, 1.508121e-11, 1.507868e-11, 1.508303e-11, 
    1.50828e-11, 1.508303e-11, 1.508302e-11, 1.508303e-11, 1.508245e-11, 
    1.508286e-11, 1.508178e-11, 1.519347e-11, 1.518801e-11, 1.520264e-11, 
    1.520927e-11, 1.521294e-11, 1.521521e-11, 1.52149e-11, 1.52143e-11, 
    1.521094e-11, 1.520728e-11, 1.520414e-11, 1.520186e-11, 1.519946e-11, 
    1.519118e-11, 1.518614e-11, 1.508159e-11, 1.508083e-11, 1.508203e-11, 
    1.508275e-11, 1.508297e-11, 1.508302e-11, 1.508281e-11, 1.5082e-11, 
    1.508303e-11, 1.508032e-11, 1.508157e-11, 1.519876e-11, 1.52057e-11, 
    1.520824e-11, 1.52103e-11, 1.521466e-11, 1.521174e-11, 1.521294e-11, 
    1.520998e-11, 1.52079e-11, 1.520895e-11, 1.520179e-11, 1.520477e-11, 
    1.518582e-11, 1.519501e-11, 1.508268e-11, 1.5081e-11, 1.508288e-11, 
    1.508219e-11, 1.508303e-11, 1.508235e-11, 1.508266e-11, 1.508218e-11, 
    1.508253e-11, 1.508063e-11, 1.508227e-11, 1.508303e-11, 1.520897e-11, 
    1.520881e-11, 1.520801e-11, 1.521135e-11, 1.521154e-11, 1.521422e-11, 
    1.521185e-11, 1.521076e-11, 1.520777e-11, 1.520584e-11, 1.520388e-11, 
    1.519913e-11, 1.519305e-11, 1.5183e-11, 1.508115e-11, 1.508254e-11, 
    1.508179e-11, 1.508247e-11, 1.508169e-11, 1.508122e-11, 1.508238e-11, 
    1.508286e-11, 1.508099e-11, 1.508128e-11, 1.50828e-11, 1.508125e-11, 
    1.520869e-11, 1.520965e-11, 1.521271e-11, 1.521035e-11, 1.521449e-11, 
    1.521226e-11, 1.521088e-11, 1.520471e-11, 1.520317e-11, 1.520167e-11, 
    1.519852e-11, 1.519409e-11, 1.518512e-11, 1.508069e-11, 1.508278e-11, 
    1.508269e-11, 1.508272e-11, 1.508293e-11, 1.508223e-11, 1.508298e-11, 
    1.508302e-11, 1.508286e-11, 1.508132e-11, 1.508237e-11, 1.508129e-11, 
    1.508204e-11, 1.520934e-11, 1.520769e-11, 1.520859e-11, 1.520686e-11, 
    1.520809e-11, 1.520221e-11, 1.520023e-11, 1.518941e-11, 1.519418e-11, 
    1.518637e-11, 1.519344e-11, 1.519226e-11, 1.518609e-11, 1.519308e-11, 
    1.508049e-11, 1.518826e-11, 1.508293e-11, 1.507979e-11, 1.508298e-11, 
    1.508277e-11, 1.508303e-11, 1.508287e-11, 1.508213e-11, 1.50791e-11, 
    1.507999e-11, 1.507619e-11, 1.520503e-11, 1.520253e-11, 1.520276e-11, 
    1.519995e-11, 1.519773e-11, 1.519247e-11, 1.518263e-11, 1.518654e-11, 
    1.507943e-11, 1.50801e-11, 1.518871e-11, 1.518211e-11, 1.520074e-11, 
    1.51982e-11, 1.519974e-11, 1.520484e-11, 1.518566e-11, 1.519657e-11, 
    1.508119e-11, 1.518184e-11, 1.508292e-11, 1.508213e-11, 1.508044e-11, 
    1.50755e-11, 1.506837e-11, 1.505679e-11, 1.520108e-11, 1.520288e-11, 
    1.51996e-11, 1.519456e-11, 1.518931e-11, 1.518141e-11, 1.507878e-11, 
    1.507954e-11, 1.508116e-11, 1.508215e-11, 1.507976e-11, 1.508234e-11, 
    1.519759e-11, 1.51846e-11, 1.520353e-11, 1.519865e-11, 1.519487e-11, 
    1.519657e-11, 1.518698e-11, 1.518442e-11, 1.508163e-11, 1.507947e-11, 
    1.507697e-11, 1.508279e-11, 1.504553e-11, 1.506279e-11, 1.520348e-11, 
    1.520109e-11, 1.51914e-11, 1.519629e-11, 1.507863e-11, 1.508057e-11, 
    1.508174e-11, 1.50827e-11, 1.508277e-11, 1.5083e-11, 1.50825e-11, 
    1.508299e-11, 1.518139e-11, 1.508135e-11, 1.519262e-11, 1.51886e-11, 
    1.519049e-11, 1.519249e-11, 1.518605e-11, 1.507981e-11, 1.507989e-11, 
    1.508088e-11, 1.508268e-11, 1.507867e-11, 1.507561e-11, 1.508293e-11, 
    1.519829e-11, 1.519282e-11, 1.519199e-11, 1.519422e-11, 1.50804e-11, 
    1.518373e-11, 1.5083e-11, 1.508238e-11, 1.508299e-11, 1.508295e-11, 
    1.50829e-11, 1.508199e-11, 1.508102e-11, 1.518342e-11, 1.518953e-11, 
    1.519391e-11, 1.519293e-11, 1.518799e-11, 1.508002e-11, 1.508277e-11, 
    1.508242e-11, 1.508302e-11, 1.518212e-11, 1.508143e-11, 1.508031e-11, 
    1.508262e-11, 1.518665e-11, 1.508208e-11, 1.51901e-11, 1.518864e-11, 
    1.518386e-11, 1.508159e-11, 1.50822e-11, 1.508267e-11, 1.50824e-11, 
    1.508013e-11, 1.507961e-11, 1.518398e-11, 1.518535e-11, 1.518896e-11, 
    1.519177e-11, 1.518921e-11, 1.518637e-11, 1.508013e-11, 1.508254e-11, 
    1.508287e-11, 1.508257e-11, 1.507895e-11, 1.508216e-11, 1.507552e-11, 
    1.508159e-11, 1.506787e-11, 1.508228e-11, 1.50817e-11, 1.518363e-11, 
    1.507877e-11, 1.508113e-11, 1.508298e-11, 1.508262e-11, 1.508289e-11, 
    1.507959e-11, 1.518781e-11, 1.518993e-11, 1.519365e-11, 1.518984e-11, 
    1.519016e-11, 1.518625e-11, 1.518754e-11, 1.508025e-11, 1.518295e-11, 
    1.508289e-11, 1.50829e-11, 1.507666e-11, 1.506792e-11, 1.50549e-11, 
    1.504775e-11, 1.50454e-11, 1.504439e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931945e-23, 1.931947e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.93194e-23, 1.931941e-23, 1.931939e-23, 1.93194e-23, 1.93194e-23, 
    1.931941e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931945e-23, 1.931944e-23, 1.931946e-23, 
    1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931945e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.931941e-23, 1.93194e-23, 1.931942e-23, 1.931941e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.93194e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931941e-23, 1.931942e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931941e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931944e-23, 1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.93194e-23, 
    1.93194e-23, 1.931939e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931943e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.93194e-23, 
    1.931939e-23, 1.931938e-23, 1.931937e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931945e-23, 1.931944e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 
    1.931939e-23, 1.931941e-23, 1.931936e-23, 1.931938e-23, 1.931946e-23, 
    1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931939e-23, 1.931942e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 
    1.931944e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 
    1.931942e-23, 1.931944e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931941e-23, 1.931941e-23, 1.93194e-23, 1.931941e-23, 1.931939e-23, 
    1.93194e-23, 1.931938e-23, 1.931942e-23, 1.93194e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 
    1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931941e-23, 1.931939e-23, 1.931938e-23, 1.931937e-23, 
    1.931937e-23, 1.931936e-23, 1.931936e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.975377e-24, 1.975379e-24, 1.975374e-24, 1.975376e-24, 1.975372e-24, 
    1.975375e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975371e-24, 
    1.975369e-24, 1.975371e-24, 1.975368e-24, 1.97537e-24, 1.975369e-24, 
    1.975371e-24, 1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975378e-24, 
    1.975378e-24, 1.975379e-24, 1.97538e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 
    1.975375e-24, 1.975376e-24, 1.975373e-24, 1.975374e-24, 1.975371e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 1.975378e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975377e-24, 
    1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975373e-24, 
    1.975371e-24, 1.975373e-24, 1.975373e-24, 1.975377e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975375e-24, 1.975376e-24, 1.975372e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 1.97537e-24, 
    1.975371e-24, 1.97537e-24, 1.975372e-24, 1.975371e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 1.975372e-24, 
    1.975373e-24, 1.975372e-24, 1.975373e-24, 1.975373e-24, 1.97537e-24, 
    1.975372e-24, 1.97537e-24, 1.97537e-24, 1.975371e-24, 1.97537e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975371e-24, 1.975372e-24, 1.97537e-24, 1.97537e-24, 1.97537e-24, 
    1.97537e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975375e-24, 1.975376e-24, 
    1.975375e-24, 1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975376e-24, 
    1.975373e-24, 1.975375e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.97537e-24, 1.975369e-24, 
    1.975369e-24, 1.975368e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975375e-24, 1.975374e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 
    1.975373e-24, 1.975374e-24, 1.975371e-24, 1.975372e-24, 1.975369e-24, 
    1.975368e-24, 1.975367e-24, 1.975365e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975377e-24, 1.975374e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975374e-24, 
    1.975368e-24, 1.975371e-24, 1.975365e-24, 1.975366e-24, 1.975378e-24, 
    1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975374e-24, 1.975373e-24, 
    1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975372e-24, 1.975374e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975368e-24, 1.975372e-24, 
    1.975377e-24, 1.975376e-24, 1.975376e-24, 1.975376e-24, 1.975373e-24, 
    1.975374e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975373e-24, 1.975374e-24, 1.975375e-24, 
    1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975374e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975375e-24, 1.975373e-24, 1.975375e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975373e-24, 1.975374e-24, 1.975374e-24, 1.975375e-24, 1.975375e-24, 
    1.975376e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975371e-24, 1.975371e-24, 1.975369e-24, 1.97537e-24, 1.975368e-24, 
    1.97537e-24, 1.975367e-24, 1.975372e-24, 1.97537e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 
    1.975374e-24, 1.975375e-24, 1.975375e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975374e-24, 
    1.975372e-24, 1.975371e-24, 1.975368e-24, 1.975367e-24, 1.975365e-24, 
    1.975365e-24, 1.975365e-24, 1.975364e-24 ;

 CONC_CH4_SAT =
  8.378757e-08, 8.389566e-08, 8.387463e-08, 8.396173e-08, 8.391338e-08, 
    8.397043e-08, 8.380944e-08, 8.389999e-08, 8.384217e-08, 8.379723e-08, 
    8.413043e-08, 8.39656e-08, 8.43004e-08, 8.419587e-08, 8.445806e-08, 
    8.428423e-08, 8.449302e-08, 8.445291e-08, 8.457318e-08, 8.453875e-08, 
    8.469247e-08, 8.458905e-08, 8.477171e-08, 8.466773e-08, 8.468406e-08, 
    8.458566e-08, 8.399869e-08, 8.410999e-08, 8.399212e-08, 8.4008e-08, 
    8.400085e-08, 8.391443e-08, 8.387091e-08, 8.377921e-08, 8.379584e-08, 
    8.386314e-08, 8.401514e-08, 8.396351e-08, 8.409324e-08, 8.409032e-08, 
    8.423437e-08, 8.416949e-08, 8.441094e-08, 8.434231e-08, 8.454019e-08, 
    8.449053e-08, 8.453788e-08, 8.452351e-08, 8.453807e-08, 8.446521e-08, 
    8.449645e-08, 8.443224e-08, 8.418166e-08, 8.425545e-08, 8.403509e-08, 
    8.390224e-08, 8.381344e-08, 8.375042e-08, 8.375934e-08, 8.377636e-08, 
    8.386353e-08, 8.394523e-08, 8.400743e-08, 8.404899e-08, 8.40899e-08, 
    8.42138e-08, 8.427895e-08, 8.442486e-08, 8.439843e-08, 8.444311e-08, 
    8.448558e-08, 8.455695e-08, 8.45452e-08, 8.457664e-08, 8.444184e-08, 
    8.453152e-08, 8.438339e-08, 8.442397e-08, 8.410147e-08, 8.397743e-08, 
    8.392499e-08, 8.387869e-08, 8.37662e-08, 8.384394e-08, 8.381332e-08, 
    8.388604e-08, 8.393224e-08, 8.390937e-08, 8.405013e-08, 8.399548e-08, 
    8.428281e-08, 8.415929e-08, 8.448063e-08, 8.440384e-08, 8.4499e-08, 
    8.445045e-08, 8.453364e-08, 8.445878e-08, 8.458829e-08, 8.46165e-08, 
    8.459724e-08, 8.467102e-08, 8.445463e-08, 8.453792e-08, 8.390875e-08, 
    8.391249e-08, 8.392982e-08, 8.385359e-08, 8.384889e-08, 8.377877e-08, 
    8.384113e-08, 8.386769e-08, 8.393488e-08, 8.397465e-08, 8.40124e-08, 
    8.409527e-08, 8.41877e-08, 8.431648e-08, 8.440883e-08, 8.447068e-08, 
    8.443273e-08, 8.446624e-08, 8.442881e-08, 8.441123e-08, 8.460596e-08, 
    8.449677e-08, 8.466041e-08, 8.465136e-08, 8.45774e-08, 8.465238e-08, 
    8.39151e-08, 8.389363e-08, 8.381915e-08, 8.387745e-08, 8.377112e-08, 
    8.383073e-08, 8.3865e-08, 8.399672e-08, 8.40255e-08, 8.405231e-08, 
    8.41051e-08, 8.417281e-08, 8.429135e-08, 8.439427e-08, 8.448804e-08, 
    8.448117e-08, 8.448359e-08, 8.450456e-08, 8.445266e-08, 8.451306e-08, 
    8.452324e-08, 8.44967e-08, 8.465015e-08, 8.460636e-08, 8.465117e-08, 
    8.462266e-08, 8.390059e-08, 8.393669e-08, 8.39172e-08, 8.395387e-08, 
    8.392807e-08, 8.404279e-08, 8.407712e-08, 8.423726e-08, 8.41715e-08, 
    8.4276e-08, 8.418209e-08, 8.419877e-08, 8.427959e-08, 8.418714e-08, 
    8.438869e-08, 8.425229e-08, 8.450537e-08, 8.436953e-08, 8.451388e-08, 
    8.448763e-08, 8.453103e-08, 8.45699e-08, 8.461868e-08, 8.470866e-08, 
    8.468782e-08, 8.476288e-08, 8.39904e-08, 8.403715e-08, 8.403295e-08, 
    8.408176e-08, 8.411785e-08, 8.419583e-08, 8.432073e-08, 8.427378e-08, 
    8.435988e-08, 8.437721e-08, 8.424631e-08, 8.432676e-08, 8.406834e-08, 
    8.411029e-08, 8.408526e-08, 8.399414e-08, 8.428472e-08, 8.41359e-08, 
    8.441037e-08, 8.432988e-08, 8.456438e-08, 8.4448e-08, 8.467637e-08, 
    8.477382e-08, 8.486492e-08, 8.497159e-08, 8.406255e-08, 8.403082e-08, 
    8.408754e-08, 8.416605e-08, 8.423851e-08, 8.433481e-08, 8.434461e-08, 
    8.436268e-08, 8.440936e-08, 8.444861e-08, 8.436848e-08, 8.445843e-08, 
    8.412019e-08, 8.429758e-08, 8.401889e-08, 8.410312e-08, 8.416139e-08, 
    8.413576e-08, 8.426839e-08, 8.429962e-08, 8.442652e-08, 8.436087e-08, 
    8.474986e-08, 8.457823e-08, 8.505233e-08, 8.492047e-08, 8.401975e-08, 
    8.40624e-08, 8.421063e-08, 8.414015e-08, 8.434118e-08, 8.439066e-08, 
    8.443077e-08, 8.448212e-08, 8.44876e-08, 8.451799e-08, 8.44682e-08, 
    8.451598e-08, 8.433501e-08, 8.441597e-08, 8.419361e-08, 8.424784e-08, 
    8.422287e-08, 8.419553e-08, 8.427988e-08, 8.436977e-08, 8.437154e-08, 
    8.440039e-08, 8.448182e-08, 8.434199e-08, 8.477222e-08, 8.45073e-08, 
    8.410887e-08, 8.4191e-08, 8.420255e-08, 8.417079e-08, 8.438571e-08, 
    8.430791e-08, 8.451723e-08, 8.446071e-08, 8.455323e-08, 8.450729e-08, 
    8.450053e-08, 8.444142e-08, 8.440461e-08, 8.431151e-08, 8.423567e-08, 
    8.417538e-08, 8.41894e-08, 8.42556e-08, 8.437523e-08, 8.448816e-08, 
    8.446347e-08, 8.45462e-08, 8.432664e-08, 8.441891e-08, 8.43833e-08, 
    8.447604e-08, 8.427256e-08, 8.44463e-08, 8.422814e-08, 8.424727e-08, 
    8.430637e-08, 8.442525e-08, 8.445132e-08, 8.447937e-08, 8.446204e-08, 
    8.437824e-08, 8.436444e-08, 8.43049e-08, 8.428854e-08, 8.424309e-08, 
    8.42055e-08, 8.423989e-08, 8.427599e-08, 8.437822e-08, 8.447034e-08, 
    8.457048e-08, 8.459489e-08, 8.471187e-08, 8.461686e-08, 8.477372e-08, 
    8.464069e-08, 8.487054e-08, 8.445615e-08, 8.46365e-08, 8.430901e-08, 
    8.434432e-08, 8.440838e-08, 8.455465e-08, 8.44756e-08, 8.456797e-08, 
    8.436388e-08, 8.425796e-08, 8.423034e-08, 8.417907e-08, 8.423152e-08, 
    8.422725e-08, 8.427739e-08, 8.426127e-08, 8.438161e-08, 8.431697e-08, 
    8.450041e-08, 8.45672e-08, 8.475507e-08, 8.486989e-08, 8.49862e-08, 
    8.503752e-08, 8.505311e-08, 8.505963e-08,
  2.310813e-10, 2.316804e-10, 2.315638e-10, 2.320471e-10, 2.317787e-10, 
    2.320954e-10, 2.312024e-10, 2.317045e-10, 2.313838e-10, 2.311347e-10, 
    2.329852e-10, 2.320686e-10, 2.339321e-10, 2.333492e-10, 2.348123e-10, 
    2.338419e-10, 2.350076e-10, 2.347834e-10, 2.354558e-10, 2.352632e-10, 
    2.361242e-10, 2.355447e-10, 2.365685e-10, 2.359854e-10, 2.36077e-10, 
    2.355257e-10, 2.322523e-10, 2.328714e-10, 2.322158e-10, 2.323041e-10, 
    2.322643e-10, 2.317846e-10, 2.315433e-10, 2.310349e-10, 2.31127e-10, 
    2.315001e-10, 2.323438e-10, 2.32057e-10, 2.327779e-10, 2.327616e-10, 
    2.335637e-10, 2.332022e-10, 2.345489e-10, 2.341658e-10, 2.352712e-10, 
    2.349936e-10, 2.352584e-10, 2.35178e-10, 2.352594e-10, 2.348521e-10, 
    2.350267e-10, 2.346678e-10, 2.332701e-10, 2.336813e-10, 2.324546e-10, 
    2.317171e-10, 2.312246e-10, 2.308755e-10, 2.309249e-10, 2.310191e-10, 
    2.315023e-10, 2.319554e-10, 2.323008e-10, 2.325318e-10, 2.327592e-10, 
    2.334494e-10, 2.338124e-10, 2.346267e-10, 2.34479e-10, 2.347287e-10, 
    2.349659e-10, 2.353651e-10, 2.352993e-10, 2.354753e-10, 2.347215e-10, 
    2.352228e-10, 2.343951e-10, 2.346217e-10, 2.32824e-10, 2.321342e-10, 
    2.318433e-10, 2.315863e-10, 2.309629e-10, 2.313937e-10, 2.312239e-10, 
    2.31627e-10, 2.318833e-10, 2.317564e-10, 2.325381e-10, 2.322345e-10, 
    2.33834e-10, 2.331455e-10, 2.349383e-10, 2.345093e-10, 2.350409e-10, 
    2.347696e-10, 2.352347e-10, 2.348161e-10, 2.355405e-10, 2.356984e-10, 
    2.355905e-10, 2.360038e-10, 2.347929e-10, 2.352586e-10, 2.31753e-10, 
    2.317737e-10, 2.318699e-10, 2.314471e-10, 2.314211e-10, 2.310325e-10, 
    2.31378e-10, 2.315253e-10, 2.31898e-10, 2.321188e-10, 2.323285e-10, 
    2.327892e-10, 2.333037e-10, 2.340217e-10, 2.345371e-10, 2.348826e-10, 
    2.346706e-10, 2.348578e-10, 2.346486e-10, 2.345504e-10, 2.356395e-10, 
    2.350285e-10, 2.359443e-10, 2.358936e-10, 2.354796e-10, 2.358993e-10, 
    2.317882e-10, 2.316691e-10, 2.312563e-10, 2.315794e-10, 2.309901e-10, 
    2.313204e-10, 2.315104e-10, 2.322415e-10, 2.324013e-10, 2.325503e-10, 
    2.328439e-10, 2.332207e-10, 2.338815e-10, 2.344559e-10, 2.349796e-10, 
    2.349412e-10, 2.349548e-10, 2.35072e-10, 2.347819e-10, 2.351196e-10, 
    2.351765e-10, 2.350281e-10, 2.358868e-10, 2.356416e-10, 2.358926e-10, 
    2.357328e-10, 2.317078e-10, 2.31908e-10, 2.317999e-10, 2.320034e-10, 
    2.318603e-10, 2.324975e-10, 2.326884e-10, 2.3358e-10, 2.332135e-10, 
    2.337959e-10, 2.332724e-10, 2.333654e-10, 2.338161e-10, 2.333005e-10, 
    2.344248e-10, 2.336638e-10, 2.350765e-10, 2.34318e-10, 2.351241e-10, 
    2.349773e-10, 2.3522e-10, 2.354376e-10, 2.357106e-10, 2.362148e-10, 
    2.36098e-10, 2.365189e-10, 2.322062e-10, 2.324661e-10, 2.324426e-10, 
    2.32714e-10, 2.329148e-10, 2.33349e-10, 2.340454e-10, 2.337834e-10, 
    2.342638e-10, 2.343606e-10, 2.336303e-10, 2.340791e-10, 2.326394e-10, 
    2.328729e-10, 2.327335e-10, 2.322271e-10, 2.338446e-10, 2.330153e-10, 
    2.345458e-10, 2.340965e-10, 2.354066e-10, 2.34756e-10, 2.360338e-10, 
    2.365804e-10, 2.370918e-10, 2.376916e-10, 2.326072e-10, 2.324308e-10, 
    2.327461e-10, 2.331832e-10, 2.335868e-10, 2.34124e-10, 2.341786e-10, 
    2.342795e-10, 2.3454e-10, 2.347593e-10, 2.343119e-10, 2.348142e-10, 
    2.329281e-10, 2.339162e-10, 2.323646e-10, 2.32833e-10, 2.331572e-10, 
    2.330144e-10, 2.337534e-10, 2.339276e-10, 2.346359e-10, 2.342694e-10, 
    2.364461e-10, 2.354843e-10, 2.38146e-10, 2.374041e-10, 2.323693e-10, 
    2.326063e-10, 2.334315e-10, 2.330389e-10, 2.341595e-10, 2.344357e-10, 
    2.346596e-10, 2.349466e-10, 2.349772e-10, 2.351471e-10, 2.348687e-10, 
    2.351359e-10, 2.341251e-10, 2.345769e-10, 2.333365e-10, 2.336389e-10, 
    2.334996e-10, 2.333473e-10, 2.338174e-10, 2.343191e-10, 2.343289e-10, 
    2.3449e-10, 2.349453e-10, 2.34164e-10, 2.365717e-10, 2.350877e-10, 
    2.328648e-10, 2.333222e-10, 2.333864e-10, 2.332095e-10, 2.34408e-10, 
    2.339739e-10, 2.351428e-10, 2.348269e-10, 2.353442e-10, 2.350873e-10, 
    2.350495e-10, 2.347191e-10, 2.345136e-10, 2.33994e-10, 2.33571e-10, 
    2.33235e-10, 2.333131e-10, 2.336821e-10, 2.343496e-10, 2.349804e-10, 
    2.348424e-10, 2.353049e-10, 2.340783e-10, 2.345934e-10, 2.343946e-10, 
    2.349126e-10, 2.337767e-10, 2.347468e-10, 2.33529e-10, 2.336356e-10, 
    2.339653e-10, 2.34629e-10, 2.347744e-10, 2.349313e-10, 2.348343e-10, 
    2.343664e-10, 2.342893e-10, 2.33957e-10, 2.338658e-10, 2.336123e-10, 
    2.334028e-10, 2.335944e-10, 2.337958e-10, 2.343662e-10, 2.348808e-10, 
    2.354408e-10, 2.355774e-10, 2.362331e-10, 2.357006e-10, 2.365802e-10, 
    2.358344e-10, 2.371237e-10, 2.348016e-10, 2.358106e-10, 2.3398e-10, 
    2.34177e-10, 2.345348e-10, 2.353523e-10, 2.349101e-10, 2.354268e-10, 
    2.342862e-10, 2.336953e-10, 2.335413e-10, 2.332556e-10, 2.335478e-10, 
    2.33524e-10, 2.338035e-10, 2.337137e-10, 2.343852e-10, 2.340244e-10, 
    2.350488e-10, 2.354225e-10, 2.364751e-10, 2.371198e-10, 2.377737e-10, 
    2.380625e-10, 2.381504e-10, 2.381871e-10,
  1.303049e-13, 1.307562e-13, 1.306683e-13, 1.310326e-13, 1.308303e-13, 
    1.31069e-13, 1.303961e-13, 1.307743e-13, 1.305327e-13, 1.303451e-13, 
    1.317404e-13, 1.310488e-13, 1.324674e-13, 1.320154e-13, 1.331515e-13, 
    1.323973e-13, 1.333034e-13, 1.33129e-13, 1.336523e-13, 1.335024e-13, 
    1.341729e-13, 1.337215e-13, 1.345193e-13, 1.340647e-13, 1.341361e-13, 
    1.337067e-13, 1.311873e-13, 1.316545e-13, 1.311598e-13, 1.312264e-13, 
    1.311964e-13, 1.308347e-13, 1.306528e-13, 1.302699e-13, 1.303393e-13, 
    1.306203e-13, 1.312563e-13, 1.3104e-13, 1.315839e-13, 1.315716e-13, 
    1.321812e-13, 1.319043e-13, 1.329467e-13, 1.326491e-13, 1.335086e-13, 
    1.332925e-13, 1.334986e-13, 1.33436e-13, 1.334994e-13, 1.331825e-13, 
    1.333183e-13, 1.330392e-13, 1.319556e-13, 1.322725e-13, 1.3134e-13, 
    1.307838e-13, 1.304128e-13, 1.3015e-13, 1.301871e-13, 1.302581e-13, 
    1.306219e-13, 1.309635e-13, 1.312239e-13, 1.313982e-13, 1.315698e-13, 
    1.320924e-13, 1.323744e-13, 1.330072e-13, 1.328924e-13, 1.330865e-13, 
    1.33271e-13, 1.335816e-13, 1.335304e-13, 1.336674e-13, 1.330809e-13, 
    1.334709e-13, 1.328272e-13, 1.330033e-13, 1.316187e-13, 1.310983e-13, 
    1.308789e-13, 1.306852e-13, 1.302157e-13, 1.305401e-13, 1.304123e-13, 
    1.307159e-13, 1.309091e-13, 1.308135e-13, 1.31403e-13, 1.311739e-13, 
    1.323911e-13, 1.318615e-13, 1.332495e-13, 1.329159e-13, 1.333294e-13, 
    1.331183e-13, 1.334801e-13, 1.331545e-13, 1.337182e-13, 1.338412e-13, 
    1.337572e-13, 1.340791e-13, 1.331365e-13, 1.334988e-13, 1.308109e-13, 
    1.308265e-13, 1.30899e-13, 1.305804e-13, 1.305608e-13, 1.302681e-13, 
    1.305283e-13, 1.306393e-13, 1.309201e-13, 1.310867e-13, 1.312448e-13, 
    1.315924e-13, 1.31981e-13, 1.325371e-13, 1.329376e-13, 1.332062e-13, 
    1.330414e-13, 1.331869e-13, 1.330243e-13, 1.329479e-13, 1.337952e-13, 
    1.333197e-13, 1.340328e-13, 1.339932e-13, 1.336707e-13, 1.339977e-13, 
    1.308374e-13, 1.307476e-13, 1.304366e-13, 1.3068e-13, 1.302362e-13, 
    1.304849e-13, 1.306281e-13, 1.311791e-13, 1.312997e-13, 1.314121e-13, 
    1.316337e-13, 1.319183e-13, 1.324281e-13, 1.328744e-13, 1.332817e-13, 
    1.332518e-13, 1.332623e-13, 1.333535e-13, 1.331279e-13, 1.333906e-13, 
    1.334348e-13, 1.333194e-13, 1.33988e-13, 1.337969e-13, 1.339924e-13, 
    1.33868e-13, 1.307768e-13, 1.309277e-13, 1.308462e-13, 1.309996e-13, 
    1.308917e-13, 1.313722e-13, 1.315163e-13, 1.321938e-13, 1.319128e-13, 
    1.323616e-13, 1.319574e-13, 1.320276e-13, 1.323773e-13, 1.319786e-13, 
    1.328503e-13, 1.322589e-13, 1.333571e-13, 1.327672e-13, 1.333941e-13, 
    1.332799e-13, 1.334687e-13, 1.336381e-13, 1.338507e-13, 1.342435e-13, 
    1.341525e-13, 1.344806e-13, 1.311526e-13, 1.313486e-13, 1.313309e-13, 
    1.315357e-13, 1.316873e-13, 1.320152e-13, 1.325555e-13, 1.323519e-13, 
    1.327252e-13, 1.328004e-13, 1.322329e-13, 1.325816e-13, 1.314794e-13, 
    1.316556e-13, 1.315504e-13, 1.311683e-13, 1.323994e-13, 1.317632e-13, 
    1.329443e-13, 1.325952e-13, 1.33614e-13, 1.331078e-13, 1.341024e-13, 
    1.345287e-13, 1.349277e-13, 1.353963e-13, 1.314551e-13, 1.31322e-13, 
    1.315599e-13, 1.318899e-13, 1.321992e-13, 1.326165e-13, 1.32659e-13, 
    1.327374e-13, 1.329399e-13, 1.331103e-13, 1.327626e-13, 1.33153e-13, 
    1.316973e-13, 1.324551e-13, 1.31272e-13, 1.316255e-13, 1.318703e-13, 
    1.317625e-13, 1.323285e-13, 1.324639e-13, 1.330144e-13, 1.327295e-13, 
    1.344238e-13, 1.336744e-13, 1.357515e-13, 1.351716e-13, 1.312756e-13, 
    1.314544e-13, 1.320785e-13, 1.31781e-13, 1.326442e-13, 1.328588e-13, 
    1.330328e-13, 1.33256e-13, 1.332798e-13, 1.33412e-13, 1.331954e-13, 
    1.334033e-13, 1.326174e-13, 1.329685e-13, 1.320058e-13, 1.322396e-13, 
    1.321314e-13, 1.320139e-13, 1.323783e-13, 1.327682e-13, 1.327758e-13, 
    1.32901e-13, 1.33255e-13, 1.326477e-13, 1.345218e-13, 1.333657e-13, 
    1.316495e-13, 1.319949e-13, 1.320435e-13, 1.319098e-13, 1.328373e-13, 
    1.324999e-13, 1.334087e-13, 1.331629e-13, 1.335654e-13, 1.333654e-13, 
    1.333361e-13, 1.330791e-13, 1.329193e-13, 1.325155e-13, 1.321869e-13, 
    1.319291e-13, 1.319881e-13, 1.322732e-13, 1.327919e-13, 1.332823e-13, 
    1.331749e-13, 1.335348e-13, 1.325811e-13, 1.329814e-13, 1.328269e-13, 
    1.332296e-13, 1.323466e-13, 1.331005e-13, 1.321542e-13, 1.32237e-13, 
    1.324932e-13, 1.33009e-13, 1.331221e-13, 1.332441e-13, 1.331686e-13, 
    1.328049e-13, 1.32745e-13, 1.324868e-13, 1.324159e-13, 1.32219e-13, 
    1.320563e-13, 1.322051e-13, 1.323615e-13, 1.328048e-13, 1.332048e-13, 
    1.336406e-13, 1.337469e-13, 1.342577e-13, 1.338429e-13, 1.345284e-13, 
    1.33947e-13, 1.349526e-13, 1.331432e-13, 1.339285e-13, 1.325046e-13, 
    1.326578e-13, 1.329357e-13, 1.335717e-13, 1.332276e-13, 1.336297e-13, 
    1.327426e-13, 1.322834e-13, 1.321638e-13, 1.319447e-13, 1.321688e-13, 
    1.321504e-13, 1.323675e-13, 1.322977e-13, 1.328195e-13, 1.325391e-13, 
    1.333355e-13, 1.336263e-13, 1.344465e-13, 1.349496e-13, 1.354604e-13, 
    1.356862e-13, 1.357549e-13, 1.357837e-13,
  1.914467e-17, 1.921998e-17, 1.920532e-17, 1.926614e-17, 1.923236e-17, 
    1.927223e-17, 1.915989e-17, 1.922301e-17, 1.918269e-17, 1.915139e-17, 
    1.93849e-17, 1.926885e-17, 1.95112e-17, 1.943266e-17, 1.963016e-17, 
    1.949901e-17, 1.965661e-17, 1.962627e-17, 1.971736e-17, 1.969125e-17, 
    1.980808e-17, 1.972941e-17, 1.986852e-17, 1.978923e-17, 1.980167e-17, 
    1.972684e-17, 1.9292e-17, 1.937006e-17, 1.92874e-17, 1.929852e-17, 
    1.929351e-17, 1.923309e-17, 1.920272e-17, 1.913885e-17, 1.915043e-17, 
    1.91973e-17, 1.930352e-17, 1.926739e-17, 1.935829e-17, 1.935623e-17, 
    1.946147e-17, 1.941339e-17, 1.959455e-17, 1.95428e-17, 1.969234e-17, 
    1.965472e-17, 1.969059e-17, 1.96797e-17, 1.969073e-17, 1.963557e-17, 
    1.96592e-17, 1.961064e-17, 1.942229e-17, 1.947733e-17, 1.93175e-17, 
    1.922459e-17, 1.916268e-17, 1.911885e-17, 1.912504e-17, 1.913687e-17, 
    1.919758e-17, 1.92546e-17, 1.929811e-17, 1.932724e-17, 1.935594e-17, 
    1.944601e-17, 1.949503e-17, 1.960507e-17, 1.958511e-17, 1.961886e-17, 
    1.965098e-17, 1.970506e-17, 1.969614e-17, 1.971999e-17, 1.96179e-17, 
    1.968577e-17, 1.957377e-17, 1.96044e-17, 1.936408e-17, 1.927712e-17, 
    1.924047e-17, 1.920815e-17, 1.912981e-17, 1.918392e-17, 1.91626e-17, 
    1.921327e-17, 1.924553e-17, 1.922956e-17, 1.932804e-17, 1.928975e-17, 
    1.949794e-17, 1.940595e-17, 1.964723e-17, 1.95892e-17, 1.966113e-17, 
    1.96244e-17, 1.968738e-17, 1.96307e-17, 1.972884e-17, 1.975026e-17, 
    1.973563e-17, 1.979173e-17, 1.962757e-17, 1.969062e-17, 1.922912e-17, 
    1.923173e-17, 1.924384e-17, 1.919064e-17, 1.918737e-17, 1.913855e-17, 
    1.918196e-17, 1.920048e-17, 1.924737e-17, 1.927518e-17, 1.93016e-17, 
    1.935971e-17, 1.942669e-17, 1.952331e-17, 1.959296e-17, 1.96397e-17, 
    1.961102e-17, 1.963634e-17, 1.960805e-17, 1.959477e-17, 1.974226e-17, 
    1.965944e-17, 1.978366e-17, 1.977677e-17, 1.972057e-17, 1.977755e-17, 
    1.923356e-17, 1.921857e-17, 1.916666e-17, 1.920728e-17, 1.913323e-17, 
    1.917472e-17, 1.91986e-17, 1.929063e-17, 1.931078e-17, 1.932957e-17, 
    1.936662e-17, 1.941582e-17, 1.950437e-17, 1.958198e-17, 1.965283e-17, 
    1.964763e-17, 1.964947e-17, 1.966534e-17, 1.962608e-17, 1.967178e-17, 
    1.967949e-17, 1.965939e-17, 1.977585e-17, 1.974256e-17, 1.977663e-17, 
    1.975494e-17, 1.922343e-17, 1.924864e-17, 1.923502e-17, 1.926065e-17, 
    1.924262e-17, 1.93229e-17, 1.934698e-17, 1.946365e-17, 1.941486e-17, 
    1.94928e-17, 1.94226e-17, 1.943478e-17, 1.949552e-17, 1.942628e-17, 
    1.957776e-17, 1.947495e-17, 1.966596e-17, 1.956332e-17, 1.96724e-17, 
    1.965253e-17, 1.96854e-17, 1.971488e-17, 1.975192e-17, 1.982041e-17, 
    1.980453e-17, 1.986177e-17, 1.928619e-17, 1.931894e-17, 1.9316e-17, 
    1.935023e-17, 1.937572e-17, 1.943264e-17, 1.952652e-17, 1.949113e-17, 
    1.955604e-17, 1.95691e-17, 1.947046e-17, 1.953107e-17, 1.934081e-17, 
    1.937027e-17, 1.935268e-17, 1.928881e-17, 1.949938e-17, 1.938888e-17, 
    1.959413e-17, 1.953343e-17, 1.971069e-17, 1.962256e-17, 1.979581e-17, 
    1.987013e-17, 1.993982e-17, 2.002167e-17, 1.933675e-17, 1.93145e-17, 
    1.935428e-17, 1.941088e-17, 1.946459e-17, 1.953714e-17, 1.954453e-17, 
    1.955815e-17, 1.959336e-17, 1.962301e-17, 1.956252e-17, 1.963044e-17, 
    1.937743e-17, 1.950906e-17, 1.930615e-17, 1.936523e-17, 1.940748e-17, 
    1.938877e-17, 1.948707e-17, 1.95106e-17, 1.960632e-17, 1.955678e-17, 
    1.985184e-17, 1.97212e-17, 2.008381e-17, 1.99824e-17, 1.930674e-17, 
    1.933664e-17, 1.944362e-17, 1.939199e-17, 1.954195e-17, 1.957925e-17, 
    1.960953e-17, 1.964836e-17, 1.965251e-17, 1.967551e-17, 1.963782e-17, 
    1.9674e-17, 1.953729e-17, 1.959835e-17, 1.943101e-17, 1.947161e-17, 
    1.945283e-17, 1.943241e-17, 1.949573e-17, 1.956349e-17, 1.956483e-17, 
    1.958659e-17, 1.964813e-17, 1.954256e-17, 1.986891e-17, 1.966742e-17, 
    1.936926e-17, 1.942911e-17, 1.943755e-17, 1.941434e-17, 1.957552e-17, 
    1.951686e-17, 1.967494e-17, 1.963216e-17, 1.970223e-17, 1.966741e-17, 
    1.96623e-17, 1.961758e-17, 1.958978e-17, 1.951956e-17, 1.946246e-17, 
    1.941769e-17, 1.942793e-17, 1.947745e-17, 1.956761e-17, 1.965293e-17, 
    1.963425e-17, 1.96969e-17, 1.953098e-17, 1.960057e-17, 1.95737e-17, 
    1.964376e-17, 1.949021e-17, 1.962127e-17, 1.945679e-17, 1.947117e-17, 
    1.951569e-17, 1.960536e-17, 1.962506e-17, 1.964628e-17, 1.963316e-17, 
    1.956988e-17, 1.955947e-17, 1.951459e-17, 1.950225e-17, 1.946803e-17, 
    1.943977e-17, 1.946562e-17, 1.94928e-17, 1.956987e-17, 1.963944e-17, 
    1.971532e-17, 1.973385e-17, 1.982286e-17, 1.975055e-17, 1.987006e-17, 
    1.976866e-17, 1.994413e-17, 1.962871e-17, 1.976547e-17, 1.951768e-17, 
    1.954432e-17, 1.959263e-17, 1.970331e-17, 1.964343e-17, 1.971341e-17, 
    1.955906e-17, 1.947922e-17, 1.945844e-17, 1.942039e-17, 1.945933e-17, 
    1.945612e-17, 1.949385e-17, 1.948172e-17, 1.957243e-17, 1.952368e-17, 
    1.96622e-17, 1.971283e-17, 1.985581e-17, 1.994362e-17, 2.00329e-17, 
    2.00724e-17, 2.008441e-17, 2.008944e-17,
  8.06949e-22, 8.105278e-22, 8.098306e-22, 8.127231e-22, 8.111165e-22, 
    8.130125e-22, 8.076722e-22, 8.106716e-22, 8.087553e-22, 8.072685e-22, 
    8.183824e-22, 8.128518e-22, 8.244231e-22, 8.206834e-22, 8.300909e-22, 
    8.238425e-22, 8.313523e-22, 8.29906e-22, 8.342732e-22, 8.330054e-22, 
    8.387427e-22, 8.348669e-22, 8.417255e-22, 8.378141e-22, 8.384272e-22, 
    8.347399e-22, 8.139539e-22, 8.176692e-22, 8.137349e-22, 8.14264e-22, 
    8.140257e-22, 8.111511e-22, 8.097068e-22, 8.06673e-22, 8.072227e-22, 
    8.094495e-22, 8.145019e-22, 8.127828e-22, 8.171105e-22, 8.170125e-22, 
    8.220568e-22, 8.197556e-22, 8.283942e-22, 8.25929e-22, 8.330574e-22, 
    8.312629e-22, 8.329738e-22, 8.324543e-22, 8.329805e-22, 8.303492e-22, 
    8.314765e-22, 8.291612e-22, 8.201839e-22, 8.228114e-22, 8.151676e-22, 
    8.107458e-22, 8.078044e-22, 8.057229e-22, 8.060171e-22, 8.065787e-22, 
    8.094626e-22, 8.121746e-22, 8.14245e-22, 8.156317e-22, 8.169984e-22, 
    8.213201e-22, 8.236535e-22, 8.288952e-22, 8.279446e-22, 8.295524e-22, 
    8.310843e-22, 8.336668e-22, 8.332385e-22, 8.344023e-22, 8.295073e-22, 
    8.327435e-22, 8.274042e-22, 8.288637e-22, 8.17384e-22, 8.132457e-22, 
    8.115012e-22, 8.099651e-22, 8.062436e-22, 8.088136e-22, 8.078004e-22, 
    8.102089e-22, 8.117428e-22, 8.109834e-22, 8.156697e-22, 8.13847e-22, 
    8.23792e-22, 8.193969e-22, 8.309057e-22, 8.281394e-22, 8.315687e-22, 
    8.298174e-22, 8.328202e-22, 8.301174e-22, 8.348384e-22, 8.358936e-22, 
    8.351728e-22, 8.379382e-22, 8.299681e-22, 8.329751e-22, 8.109627e-22, 
    8.110867e-22, 8.116625e-22, 8.09133e-22, 8.089776e-22, 8.066586e-22, 
    8.087207e-22, 8.096006e-22, 8.118306e-22, 8.131534e-22, 8.144108e-22, 
    8.17178e-22, 8.203957e-22, 8.250004e-22, 8.283187e-22, 8.305468e-22, 
    8.291793e-22, 8.303866e-22, 8.290376e-22, 8.28405e-22, 8.354991e-22, 
    8.314878e-22, 8.375402e-22, 8.372006e-22, 8.344308e-22, 8.372389e-22, 
    8.111735e-22, 8.104609e-22, 8.079935e-22, 8.099242e-22, 8.064061e-22, 
    8.083763e-22, 8.09511e-22, 8.138881e-22, 8.148477e-22, 8.157423e-22, 
    8.17507e-22, 8.198725e-22, 8.240986e-22, 8.277949e-22, 8.311729e-22, 
    8.30925e-22, 8.310124e-22, 8.317692e-22, 8.29897e-22, 8.320766e-22, 
    8.32444e-22, 8.314856e-22, 8.371552e-22, 8.355146e-22, 8.371934e-22, 
    8.361247e-22, 8.106921e-22, 8.118907e-22, 8.112432e-22, 8.124618e-22, 
    8.116043e-22, 8.15424e-22, 8.165707e-22, 8.221601e-22, 8.198265e-22, 
    8.235478e-22, 8.20199e-22, 8.207856e-22, 8.236758e-22, 8.203767e-22, 
    8.275936e-22, 8.226976e-22, 8.317986e-22, 8.26905e-22, 8.32106e-22, 
    8.311583e-22, 8.327261e-22, 8.341508e-22, 8.359758e-22, 8.393517e-22, 
    8.385689e-22, 8.413929e-22, 8.136776e-22, 8.15236e-22, 8.150962e-22, 
    8.167264e-22, 8.179425e-22, 8.206825e-22, 8.251534e-22, 8.234688e-22, 
    8.265596e-22, 8.271816e-22, 8.224847e-22, 8.253698e-22, 8.162777e-22, 
    8.176802e-22, 8.168431e-22, 8.13802e-22, 8.238606e-22, 8.185753e-22, 
    8.283741e-22, 8.254824e-22, 8.339441e-22, 8.297286e-22, 8.381387e-22, 
    8.418044e-22, 8.452474e-22, 8.492929e-22, 8.160843e-22, 8.15025e-22, 
    8.169196e-22, 8.196344e-22, 8.222053e-22, 8.256592e-22, 8.260114e-22, 
    8.2666e-22, 8.283378e-22, 8.297509e-22, 8.268678e-22, 8.30105e-22, 
    8.180231e-22, 8.243219e-22, 8.146271e-22, 8.174402e-22, 8.194707e-22, 
    8.185707e-22, 8.232756e-22, 8.243957e-22, 8.289548e-22, 8.265952e-22, 
    8.409015e-22, 8.344613e-22, 8.52369e-22, 8.473513e-22, 8.146558e-22, 
    8.160794e-22, 8.212073e-22, 8.187253e-22, 8.258885e-22, 8.276653e-22, 
    8.291085e-22, 8.309593e-22, 8.311572e-22, 8.322543e-22, 8.304571e-22, 
    8.321823e-22, 8.256666e-22, 8.285753e-22, 8.206043e-22, 8.225394e-22, 
    8.216458e-22, 8.206718e-22, 8.236875e-22, 8.269138e-22, 8.269785e-22, 
    8.280149e-22, 8.30946e-22, 8.259176e-22, 8.417424e-22, 8.318663e-22, 
    8.176331e-22, 8.205116e-22, 8.209188e-22, 8.198017e-22, 8.274873e-22, 
    8.246934e-22, 8.322269e-22, 8.301872e-22, 8.335292e-22, 8.318682e-22, 
    8.316242e-22, 8.294921e-22, 8.28167e-22, 8.248222e-22, 8.221037e-22, 
    8.199631e-22, 8.204561e-22, 8.228172e-22, 8.271103e-22, 8.311771e-22, 
    8.302862e-22, 8.33275e-22, 8.253659e-22, 8.286809e-22, 8.274004e-22, 
    8.307401e-22, 8.234249e-22, 8.296657e-22, 8.218344e-22, 8.225189e-22, 
    8.246379e-22, 8.289089e-22, 8.298485e-22, 8.308601e-22, 8.302349e-22, 
    8.272186e-22, 8.267229e-22, 8.245853e-22, 8.239977e-22, 8.223695e-22, 
    8.210247e-22, 8.222545e-22, 8.235477e-22, 8.272181e-22, 8.305339e-22, 
    8.341721e-22, 8.350855e-22, 8.394713e-22, 8.359064e-22, 8.417986e-22, 
    8.367971e-22, 8.454579e-22, 8.300214e-22, 8.366414e-22, 8.247329e-22, 
    8.260013e-22, 8.283021e-22, 8.335798e-22, 8.307243e-22, 8.340775e-22, 
    8.267032e-22, 8.229011e-22, 8.219131e-22, 8.200929e-22, 8.219551e-22, 
    8.218023e-22, 8.235983e-22, 8.230207e-22, 8.2734e-22, 8.250186e-22, 
    8.316192e-22, 8.340491e-22, 8.410984e-22, 8.454343e-22, 8.498499e-22, 
    8.518045e-22, 8.523994e-22, 8.526483e-22,
  1.042531e-26, 1.047809e-26, 1.04678e-26, 1.051049e-26, 1.048678e-26, 
    1.051477e-26, 1.043597e-26, 1.048021e-26, 1.045194e-26, 1.043002e-26, 
    1.059401e-26, 1.051239e-26, 1.068201e-26, 1.062768e-26, 1.076445e-26, 
    1.067357e-26, 1.078282e-26, 1.076177e-26, 1.08255e-26, 1.080691e-26, 
    1.089144e-26, 1.083426e-26, 1.093551e-26, 1.087774e-26, 1.088679e-26, 
    1.083238e-26, 1.052868e-26, 1.058358e-26, 1.052544e-26, 1.053326e-26, 
    1.052974e-26, 1.048729e-26, 1.046597e-26, 1.042125e-26, 1.042935e-26, 
    1.046218e-26, 1.053677e-26, 1.051138e-26, 1.057534e-26, 1.057389e-26, 
    1.064765e-26, 1.061411e-26, 1.073977e-26, 1.070392e-26, 1.080766e-26, 
    1.078153e-26, 1.080644e-26, 1.079888e-26, 1.080654e-26, 1.076822e-26, 
    1.078463e-26, 1.075093e-26, 1.062038e-26, 1.06586e-26, 1.054661e-26, 
    1.048129e-26, 1.043792e-26, 1.040725e-26, 1.041158e-26, 1.041985e-26, 
    1.046237e-26, 1.05024e-26, 1.053298e-26, 1.055348e-26, 1.057369e-26, 
    1.063693e-26, 1.067083e-26, 1.074705e-26, 1.073323e-26, 1.075662e-26, 
    1.077892e-26, 1.081656e-26, 1.08103e-26, 1.08274e-26, 1.075597e-26, 
    1.080309e-26, 1.072537e-26, 1.07466e-26, 1.057935e-26, 1.051822e-26, 
    1.049244e-26, 1.046979e-26, 1.041492e-26, 1.04528e-26, 1.043786e-26, 
    1.047339e-26, 1.049602e-26, 1.048482e-26, 1.055404e-26, 1.05271e-26, 
    1.067284e-26, 1.060887e-26, 1.077632e-26, 1.073606e-26, 1.078598e-26, 
    1.076048e-26, 1.08042e-26, 1.076485e-26, 1.083384e-26, 1.08494e-26, 
    1.083876e-26, 1.087958e-26, 1.076267e-26, 1.080646e-26, 1.048451e-26, 
    1.048634e-26, 1.049484e-26, 1.045751e-26, 1.045522e-26, 1.042104e-26, 
    1.045143e-26, 1.046441e-26, 1.049732e-26, 1.051685e-26, 1.053543e-26, 
    1.057634e-26, 1.062347e-26, 1.069041e-26, 1.073867e-26, 1.07711e-26, 
    1.07512e-26, 1.076877e-26, 1.074913e-26, 1.073993e-26, 1.084358e-26, 
    1.07848e-26, 1.08737e-26, 1.086869e-26, 1.082782e-26, 1.086926e-26, 
    1.048762e-26, 1.047711e-26, 1.044071e-26, 1.046919e-26, 1.041731e-26, 
    1.044635e-26, 1.046308e-26, 1.05277e-26, 1.054189e-26, 1.055511e-26, 
    1.058121e-26, 1.061582e-26, 1.06773e-26, 1.073105e-26, 1.078022e-26, 
    1.077661e-26, 1.077788e-26, 1.07889e-26, 1.076164e-26, 1.079338e-26, 
    1.079872e-26, 1.078477e-26, 1.086802e-26, 1.084381e-26, 1.086859e-26, 
    1.085281e-26, 1.048052e-26, 1.049821e-26, 1.048865e-26, 1.050664e-26, 
    1.049398e-26, 1.05504e-26, 1.056735e-26, 1.064914e-26, 1.061515e-26, 
    1.06693e-26, 1.06206e-26, 1.062917e-26, 1.067115e-26, 1.06232e-26, 
    1.072811e-26, 1.065694e-26, 1.078933e-26, 1.071809e-26, 1.07938e-26, 
    1.078e-26, 1.080284e-26, 1.082369e-26, 1.085061e-26, 1.090044e-26, 
    1.088889e-26, 1.093061e-26, 1.05246e-26, 1.054762e-26, 1.054556e-26, 
    1.056966e-26, 1.058761e-26, 1.062767e-26, 1.069264e-26, 1.066816e-26, 
    1.071309e-26, 1.072213e-26, 1.065386e-26, 1.069578e-26, 1.056302e-26, 
    1.058376e-26, 1.057139e-26, 1.052643e-26, 1.067384e-26, 1.059685e-26, 
    1.073948e-26, 1.069742e-26, 1.082064e-26, 1.075918e-26, 1.088253e-26, 
    1.093667e-26, 1.098912e-26, 1.105081e-26, 1.056017e-26, 1.054451e-26, 
    1.057252e-26, 1.061233e-26, 1.06498e-26, 1.069999e-26, 1.070512e-26, 
    1.071454e-26, 1.073895e-26, 1.075951e-26, 1.071756e-26, 1.076467e-26, 
    1.058877e-26, 1.068055e-26, 1.053862e-26, 1.058021e-26, 1.060994e-26, 
    1.059679e-26, 1.066536e-26, 1.068163e-26, 1.074792e-26, 1.07136e-26, 
    1.092332e-26, 1.082826e-26, 1.109781e-26, 1.102119e-26, 1.053905e-26, 
    1.05601e-26, 1.063531e-26, 1.059905e-26, 1.070333e-26, 1.072916e-26, 
    1.075017e-26, 1.07771e-26, 1.077999e-26, 1.079596e-26, 1.076979e-26, 
    1.079492e-26, 1.07001e-26, 1.07424e-26, 1.062653e-26, 1.065466e-26, 
    1.064168e-26, 1.062752e-26, 1.067134e-26, 1.071823e-26, 1.071918e-26, 
    1.073425e-26, 1.077687e-26, 1.070375e-26, 1.093573e-26, 1.079028e-26, 
    1.058307e-26, 1.062516e-26, 1.063112e-26, 1.061479e-26, 1.072657e-26, 
    1.068595e-26, 1.079556e-26, 1.076587e-26, 1.081454e-26, 1.079034e-26, 
    1.078679e-26, 1.075575e-26, 1.073646e-26, 1.068782e-26, 1.064833e-26, 
    1.061715e-26, 1.062436e-26, 1.065869e-26, 1.072109e-26, 1.078027e-26, 
    1.07673e-26, 1.081083e-26, 1.069573e-26, 1.074394e-26, 1.072531e-26, 
    1.077391e-26, 1.066752e-26, 1.075824e-26, 1.064442e-26, 1.065436e-26, 
    1.068515e-26, 1.074725e-26, 1.076093e-26, 1.077566e-26, 1.076656e-26, 
    1.072266e-26, 1.071546e-26, 1.068438e-26, 1.067584e-26, 1.065219e-26, 
    1.063266e-26, 1.065052e-26, 1.06693e-26, 1.072266e-26, 1.077091e-26, 
    1.082401e-26, 1.083748e-26, 1.090219e-26, 1.084957e-26, 1.093656e-26, 
    1.086269e-26, 1.099229e-26, 1.076343e-26, 1.086041e-26, 1.068653e-26, 
    1.070497e-26, 1.073842e-26, 1.081526e-26, 1.077368e-26, 1.08226e-26, 
    1.071517e-26, 1.06599e-26, 1.064556e-26, 1.061905e-26, 1.064617e-26, 
    1.064396e-26, 1.067004e-26, 1.066165e-26, 1.072443e-26, 1.069068e-26, 
    1.078671e-26, 1.082219e-26, 1.092625e-26, 1.099196e-26, 1.105934e-26, 
    1.108919e-26, 1.109828e-26, 1.110208e-26,
  4.215264e-32, 4.240935e-32, 4.23593e-32, 4.256717e-32, 4.245169e-32, 
    4.2588e-32, 4.220451e-32, 4.241964e-32, 4.228216e-32, 4.217559e-32, 
    4.297897e-32, 4.257644e-32, 4.341546e-32, 4.314635e-32, 4.38247e-32, 
    4.33736e-32, 4.391607e-32, 4.381144e-32, 4.412808e-32, 4.403603e-32, 
    4.445318e-32, 4.417123e-32, 4.467102e-32, 4.438561e-32, 4.443025e-32, 
    4.416198e-32, 4.265586e-32, 4.292709e-32, 4.264008e-32, 4.267816e-32, 
    4.266103e-32, 4.245414e-32, 4.235031e-32, 4.213295e-32, 4.217231e-32, 
    4.233192e-32, 4.269529e-32, 4.257154e-32, 4.288589e-32, 4.287861e-32, 
    4.324526e-32, 4.307897e-32, 4.370211e-32, 4.352417e-32, 4.40398e-32, 
    4.39097e-32, 4.403371e-32, 4.399605e-32, 4.40342e-32, 4.384351e-32, 
    4.392514e-32, 4.375758e-32, 4.311006e-32, 4.32995e-32, 4.274331e-32, 
    4.242487e-32, 4.221396e-32, 4.206494e-32, 4.208598e-32, 4.212615e-32, 
    4.233285e-32, 4.252778e-32, 4.267686e-32, 4.277684e-32, 4.287757e-32, 
    4.319209e-32, 4.336004e-32, 4.373826e-32, 4.366965e-32, 4.37858e-32, 
    4.389676e-32, 4.408399e-32, 4.405293e-32, 4.413741e-32, 4.378262e-32, 
    4.401696e-32, 4.363065e-32, 4.373606e-32, 4.290585e-32, 4.260487e-32, 
    4.247918e-32, 4.236895e-32, 4.210218e-32, 4.228629e-32, 4.221365e-32, 
    4.23865e-32, 4.249672e-32, 4.244215e-32, 4.277958e-32, 4.264817e-32, 
    4.337001e-32, 4.305287e-32, 4.388381e-32, 4.368371e-32, 4.393185e-32, 
    4.380506e-32, 4.402254e-32, 4.382677e-32, 4.416912e-32, 4.42458e-32, 
    4.419341e-32, 4.439473e-32, 4.381596e-32, 4.403377e-32, 4.244065e-32, 
    4.244955e-32, 4.249096e-32, 4.23092e-32, 4.229807e-32, 4.21319e-32, 
    4.227968e-32, 4.234278e-32, 4.250306e-32, 4.259822e-32, 4.268878e-32, 
    4.289088e-32, 4.312539e-32, 4.345712e-32, 4.369667e-32, 4.385785e-32, 
    4.375892e-32, 4.384626e-32, 4.374866e-32, 4.370294e-32, 4.42171e-32, 
    4.392594e-32, 4.436573e-32, 4.434101e-32, 4.413946e-32, 4.434379e-32, 
    4.245579e-32, 4.240462e-32, 4.222752e-32, 4.236606e-32, 4.211383e-32, 
    4.225495e-32, 4.23363e-32, 4.265105e-32, 4.272029e-32, 4.278479e-32, 
    4.291537e-32, 4.308746e-32, 4.339216e-32, 4.365878e-32, 4.39032e-32, 
    4.388524e-32, 4.389157e-32, 4.394637e-32, 4.381081e-32, 4.396866e-32, 
    4.399525e-32, 4.392583e-32, 4.43377e-32, 4.421831e-32, 4.434048e-32, 
    4.426269e-32, 4.242123e-32, 4.250737e-32, 4.246081e-32, 4.254842e-32, 
    4.248673e-32, 4.276175e-32, 4.284561e-32, 4.325258e-32, 4.30841e-32, 
    4.335248e-32, 4.311118e-32, 4.315378e-32, 4.336154e-32, 4.312412e-32, 
    4.364417e-32, 4.32912e-32, 4.39485e-32, 4.359436e-32, 4.397079e-32, 
    4.390214e-32, 4.401578e-32, 4.411914e-32, 4.425184e-32, 4.449772e-32, 
    4.444066e-32, 4.464678e-32, 4.263598e-32, 4.274823e-32, 4.273822e-32, 
    4.285732e-32, 4.294737e-32, 4.314634e-32, 4.34682e-32, 4.334688e-32, 
    4.356967e-32, 4.361454e-32, 4.327608e-32, 4.348376e-32, 4.282391e-32, 
    4.292813e-32, 4.286597e-32, 4.264489e-32, 4.337498e-32, 4.299319e-32, 
    4.370066e-32, 4.349194e-32, 4.410412e-32, 4.379853e-32, 4.44093e-32, 
    4.467668e-32, 4.493897e-32, 4.52479e-32, 4.280957e-32, 4.273309e-32, 
    4.28717e-32, 4.307007e-32, 4.325594e-32, 4.350467e-32, 4.353011e-32, 
    4.357689e-32, 4.369808e-32, 4.380025e-32, 4.35918e-32, 4.382588e-32, 
    4.295296e-32, 4.340824e-32, 4.270436e-32, 4.291026e-32, 4.305823e-32, 
    4.299294e-32, 4.3333e-32, 4.341365e-32, 4.37426e-32, 4.357224e-32, 
    4.461068e-32, 4.414159e-32, 4.548771e-32, 4.509945e-32, 4.270646e-32, 
    4.280924e-32, 4.318416e-32, 4.300417e-32, 4.352125e-32, 4.364946e-32, 
    4.37538e-32, 4.388767e-32, 4.390205e-32, 4.398152e-32, 4.385136e-32, 
    4.397633e-32, 4.35052e-32, 4.371522e-32, 4.314067e-32, 4.327997e-32, 
    4.321577e-32, 4.314558e-32, 4.336264e-32, 4.359511e-32, 4.359989e-32, 
    4.367468e-32, 4.388631e-32, 4.352335e-32, 4.467188e-32, 4.395304e-32, 
    4.292477e-32, 4.313377e-32, 4.316348e-32, 4.308235e-32, 4.36366e-32, 
    4.343505e-32, 4.397955e-32, 4.383183e-32, 4.407403e-32, 4.395356e-32, 
    4.393587e-32, 4.378153e-32, 4.36857e-32, 4.344432e-32, 4.324862e-32, 
    4.309409e-32, 4.31299e-32, 4.329993e-32, 4.360931e-32, 4.390344e-32, 
    4.38389e-32, 4.405558e-32, 4.348355e-32, 4.37228e-32, 4.363027e-32, 
    4.387182e-32, 4.33437e-32, 4.379371e-32, 4.322933e-32, 4.327854e-32, 
    4.343106e-32, 4.37392e-32, 4.380731e-32, 4.388048e-32, 4.383528e-32, 
    4.361715e-32, 4.358141e-32, 4.34273e-32, 4.338492e-32, 4.326781e-32, 
    4.317113e-32, 4.32595e-32, 4.33525e-32, 4.361716e-32, 4.385686e-32, 
    4.412067e-32, 4.41871e-32, 4.450624e-32, 4.424659e-32, 4.467597e-32, 
    4.431113e-32, 4.495465e-32, 4.38196e-32, 4.430003e-32, 4.343794e-32, 
    4.352939e-32, 4.369537e-32, 4.407754e-32, 4.387068e-32, 4.411372e-32, 
    4.358e-32, 4.330591e-32, 4.323498e-32, 4.310349e-32, 4.323799e-32, 
    4.322702e-32, 4.335622e-32, 4.331466e-32, 4.362597e-32, 4.345852e-32, 
    4.393548e-32, 4.411169e-32, 4.462522e-32, 4.495309e-32, 4.529074e-32, 
    4.544331e-32, 4.549017e-32, 4.550978e-32,
  5.564283e-38, 5.61038e-38, 5.601381e-38, 5.63881e-38, 5.618005e-38, 
    5.642569e-38, 5.573585e-38, 5.612227e-38, 5.58752e-38, 5.568402e-38, 
    5.713426e-38, 5.640484e-38, 5.792536e-38, 5.743756e-38, 5.868961e-38, 
    5.784928e-38, 5.886184e-38, 5.866477e-38, 5.92613e-38, 5.908848e-38, 
    5.986996e-38, 5.93419e-38, 6.02801e-38, 5.974323e-38, 5.982694e-38, 
    5.932462e-38, 5.654827e-38, 5.704038e-38, 5.651976e-38, 5.658852e-38, 
    5.655761e-38, 5.618442e-38, 5.599752e-38, 5.560761e-38, 5.567814e-38, 
    5.596454e-38, 5.661947e-38, 5.639606e-38, 5.696555e-38, 5.695227e-38, 
    5.761668e-38, 5.731551e-38, 5.845918e-38, 5.812548e-38, 5.90956e-38, 
    5.884992e-38, 5.908408e-38, 5.901293e-38, 5.908501e-38, 5.872515e-38, 
    5.887904e-38, 5.856345e-38, 5.737179e-38, 5.771497e-38, 5.670635e-38, 
    5.613158e-38, 5.575278e-38, 5.548583e-38, 5.552349e-38, 5.559539e-38, 
    5.596622e-38, 5.631714e-38, 5.658625e-38, 5.676709e-38, 5.695036e-38, 
    5.75202e-38, 5.782472e-38, 5.852704e-38, 5.839824e-38, 5.861647e-38, 
    5.882553e-38, 5.917898e-38, 5.912042e-38, 5.927868e-38, 5.861055e-38, 
    5.905237e-38, 5.832507e-38, 5.852299e-38, 5.700159e-38, 5.645621e-38, 
    5.62294e-38, 5.603112e-38, 5.555247e-38, 5.588258e-38, 5.575221e-38, 
    5.606275e-38, 5.626116e-38, 5.61629e-38, 5.677204e-38, 5.65344e-38, 
    5.784283e-38, 5.726819e-38, 5.880111e-38, 5.842463e-38, 5.889173e-38, 
    5.86528e-38, 5.906294e-38, 5.869367e-38, 5.933794e-38, 5.948129e-38, 
    5.938331e-38, 5.976041e-38, 5.86733e-38, 5.908416e-38, 5.616019e-38, 
    5.61762e-38, 5.625079e-38, 5.592373e-38, 5.590374e-38, 5.560572e-38, 
    5.587075e-38, 5.598408e-38, 5.627262e-38, 5.64442e-38, 5.660778e-38, 
    5.69746e-38, 5.739953e-38, 5.800114e-38, 5.844897e-38, 5.875222e-38, 
    5.8566e-38, 5.873037e-38, 5.854669e-38, 5.846079e-38, 5.942758e-38, 
    5.888052e-38, 5.9706e-38, 5.965966e-38, 5.92825e-38, 5.966488e-38, 
    5.618744e-38, 5.609535e-38, 5.577712e-38, 5.602599e-38, 5.557336e-38, 
    5.582632e-38, 5.59724e-38, 5.653952e-38, 5.666478e-38, 5.678144e-38, 
    5.701933e-38, 5.733088e-38, 5.788311e-38, 5.837778e-38, 5.883769e-38, 
    5.880384e-38, 5.881576e-38, 5.891911e-38, 5.86636e-38, 5.896117e-38, 
    5.901136e-38, 5.888036e-38, 5.965346e-38, 5.942991e-38, 5.965867e-38, 
    5.951297e-38, 5.612524e-38, 5.628035e-38, 5.619649e-38, 5.635434e-38, 
    5.624314e-38, 5.673966e-38, 5.689193e-38, 5.762986e-38, 5.732477e-38, 
    5.781106e-38, 5.737385e-38, 5.745102e-38, 5.782733e-38, 5.739731e-38, 
    5.835028e-38, 5.769981e-38, 5.892313e-38, 5.825676e-38, 5.89652e-38, 
    5.88357e-38, 5.905021e-38, 5.924458e-38, 5.949265e-38, 5.995377e-38, 
    5.984659e-38, 6.023446e-38, 5.651238e-38, 5.671525e-38, 5.669721e-38, 
    5.691341e-38, 5.707744e-38, 5.743758e-38, 5.802131e-38, 5.780098e-38, 
    5.821072e-38, 5.829482e-38, 5.767259e-38, 5.804979e-38, 5.685247e-38, 
    5.704248e-38, 5.692916e-38, 5.652844e-38, 5.785188e-38, 5.716019e-38, 
    5.845645e-38, 5.806513e-38, 5.921655e-38, 5.864039e-38, 5.978772e-38, 
    6.029066e-38, 6.078079e-38, 6.136716e-38, 5.682636e-38, 5.668794e-38, 
    5.693967e-38, 5.72993e-38, 5.763604e-38, 5.808894e-38, 5.813662e-38, 
    5.822422e-38, 5.845165e-38, 5.864374e-38, 5.82521e-38, 5.869199e-38, 
    5.70873e-38, 5.791231e-38, 5.663591e-38, 5.700985e-38, 5.72779e-38, 
    5.715981e-38, 5.777582e-38, 5.792221e-38, 5.853522e-38, 5.821554e-38, 
    6.016622e-38, 5.928639e-38, 6.183349e-38, 6.108152e-38, 5.663977e-38, 
    5.68258e-38, 5.750601e-38, 5.718013e-38, 5.812002e-38, 5.836032e-38, 
    5.855637e-38, 5.880834e-38, 5.883551e-38, 5.898545e-38, 5.873999e-38, 
    5.897567e-38, 5.808994e-38, 5.848383e-38, 5.742733e-38, 5.76796e-38, 
    5.756332e-38, 5.743622e-38, 5.78296e-38, 5.825828e-38, 5.826736e-38, 
    5.840762e-38, 5.880538e-38, 5.812396e-38, 6.028134e-38, 5.893132e-38, 
    5.70365e-38, 5.741467e-38, 5.746865e-38, 5.732167e-38, 5.833618e-38, 
    5.796108e-38, 5.898176e-38, 5.870319e-38, 5.916035e-38, 5.893269e-38, 
    5.889929e-38, 5.860851e-38, 5.842838e-38, 5.797789e-38, 5.762278e-38, 
    5.734293e-38, 5.74078e-38, 5.771577e-38, 5.828494e-38, 5.883808e-38, 
    5.871643e-38, 5.912546e-38, 5.804947e-38, 5.849802e-38, 5.832427e-38, 
    5.877852e-38, 5.779519e-38, 5.863103e-38, 5.758789e-38, 5.767705e-38, 
    5.795382e-38, 5.852876e-38, 5.865703e-38, 5.879481e-38, 5.87097e-38, 
    5.829966e-38, 5.823269e-38, 5.794702e-38, 5.786999e-38, 5.76576e-38, 
    5.748253e-38, 5.764252e-38, 5.781113e-38, 5.829973e-38, 5.875028e-38, 
    5.924742e-38, 5.937157e-38, 5.996958e-38, 5.94826e-38, 6.028904e-38, 
    5.960314e-38, 6.08098e-38, 5.867994e-38, 5.95826e-38, 5.796637e-38, 
    5.813527e-38, 5.844643e-38, 5.916681e-38, 5.877637e-38, 5.923435e-38, 
    5.823004e-38, 5.772655e-38, 5.75981e-38, 5.735993e-38, 5.760357e-38, 
    5.758369e-38, 5.781795e-38, 5.774254e-38, 5.831625e-38, 5.800377e-38, 
    5.889852e-38, 5.92306e-38, 6.019376e-38, 6.080708e-38, 6.145031e-38, 
    6.174697e-38, 6.183837e-38, 6.187663e-38,
  2.662467e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 3.082857e-44, 3.082857e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 3.082857e-44, 3.082857e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 3.082857e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 3.082857e-44, 3.082857e-44, 
    3.082857e-44, 3.082857e-44, 3.082857e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  5.604323e-06, 5.328882e-06, 5.382194e-06, 5.161834e-06, 5.283812e-06, 
    5.139907e-06, 5.548251e-06, 5.318002e-06, 5.464747e-06, 5.579419e-06, 
    4.741034e-06, 5.152058e-06, 4.32516e-06, 4.579083e-06, 3.94948e-06, 
    4.364341e-06, 3.868341e-06, 3.961165e-06, 3.684557e-06, 3.762958e-06, 
    3.418476e-06, 3.648609e-06, 3.245915e-06, 3.47283e-06, 3.436848e-06, 
    3.656311e-06, 5.068629e-06, 4.791677e-06, 5.085164e-06, 5.045381e-06, 
    5.063227e-06, 5.281278e-06, 5.391978e-06, 5.62551e-06, 5.582963e-06, 
    5.41152e-06, 5.027519e-06, 5.157106e-06, 4.832254e-06, 4.839526e-06, 
    4.484953e-06, 4.643794e-06, 4.05938e-06, 4.221542e-06, 3.759672e-06, 
    3.873844e-06, 3.765e-06, 3.797873e-06, 3.764573e-06, 3.93258e-06, 
    3.860233e-06, 4.009395e-06, 4.613907e-06, 4.433758e-06, 4.977447e-06, 
    5.312607e-06, 5.538104e-06, 5.699292e-06, 5.676449e-06, 5.632947e-06, 
    5.41052e-06, 5.203248e-06, 5.046616e-06, 4.942537e-06, 4.840572e-06, 
    4.535704e-06, 4.376967e-06, 4.026867e-06, 4.088723e-06, 3.984161e-06, 
    3.88528e-06, 3.721504e-06, 3.748263e-06, 3.676823e-06, 3.98692e-06, 
    3.779674e-06, 4.12411e-06, 4.028742e-06, 4.812879e-06, 5.122067e-06, 
    5.254922e-06, 5.371934e-06, 5.658896e-06, 5.460381e-06, 5.53846e-06, 
    5.353121e-06, 5.236089e-06, 5.293898e-06, 4.939699e-06, 5.076653e-06, 
    4.367618e-06, 4.669067e-06, 3.896762e-06, 4.075999e-06, 3.854276e-06, 
    3.966815e-06, 3.77478e-06, 3.947439e-06, 3.650391e-06, 3.587005e-06, 
    3.630267e-06, 3.465366e-06, 3.957099e-06, 3.764994e-06, 5.295517e-06, 
    5.286077e-06, 5.242161e-06, 5.435834e-06, 5.447738e-06, 5.626674e-06, 
    5.467403e-06, 5.399871e-06, 5.22933e-06, 5.129061e-06, 5.034206e-06, 
    4.827329e-06, 4.599247e-06, 4.286303e-06, 4.064286e-06, 3.919768e-06, 
    4.00815e-06, 3.93008e-06, 4.01739e-06, 4.058568e-06, 3.610694e-06, 
    3.859556e-06, 3.488872e-06, 3.508957e-06, 3.675129e-06, 3.506692e-06, 
    5.279452e-06, 5.333809e-06, 5.523477e-06, 5.37492e-06, 5.646232e-06, 
    5.494005e-06, 5.406869e-06, 5.073764e-06, 5.00131e-06, 4.93435e-06, 
    4.802859e-06, 4.635621e-06, 4.346808e-06, 4.098653e-06, 3.87956e-06, 
    3.895454e-06, 3.889855e-06, 3.841502e-06, 3.961707e-06, 3.821911e-06, 
    3.798641e-06, 3.859595e-06, 3.511651e-06, 3.609609e-06, 3.509385e-06, 
    3.573013e-06, 5.316127e-06, 5.224816e-06, 5.274109e-06, 5.181504e-06, 
    5.246698e-06, 4.958379e-06, 4.87278e-06, 4.478156e-06, 4.638891e-06, 
    4.38398e-06, 4.612791e-06, 4.571965e-06, 4.375714e-06, 4.600334e-06, 
    4.112019e-06, 4.441737e-06, 3.839627e-06, 4.157515e-06, 3.820038e-06, 
    3.880498e-06, 3.780613e-06, 3.692065e-06, 3.581958e-06, 3.382689e-06, 
    3.428369e-06, 3.264791e-06, 5.089416e-06, 4.972346e-06, 4.982639e-06, 
    4.860856e-06, 4.771336e-06, 4.579028e-06, 4.275961e-06, 4.389114e-06, 
    4.179789e-06, 4.138831e-06, 4.455736e-06, 4.261573e-06, 4.894418e-06, 
    4.790336e-06, 4.85224e-06, 5.080147e-06, 4.36293e-06, 4.726911e-06, 
    4.060696e-06, 4.253934e-06, 3.704635e-06, 3.972805e-06, 3.453634e-06, 
    3.241624e-06, 3.048194e-06, 2.830005e-06, 4.908778e-06, 4.987972e-06, 
    4.846434e-06, 4.65252e-06, 4.474833e-06, 4.242173e-06, 4.216075e-06, 
    4.173216e-06, 4.062967e-06, 3.971128e-06, 4.159685e-06, 3.948234e-06, 
    4.76626e-06, 4.331799e-06, 5.017989e-06, 4.808167e-06, 4.663891e-06, 
    4.727035e-06, 4.402114e-06, 4.326643e-06, 4.022937e-06, 4.17743e-06, 
    3.293341e-06, 3.673457e-06, 2.669976e-06, 2.933644e-06, 5.015719e-06, 
    4.909057e-06, 4.54301e-06, 4.716122e-06, 4.224226e-06, 4.107071e-06, 
    4.012748e-06, 3.893386e-06, 3.880595e-06, 3.810646e-06, 3.925535e-06, 
    3.815163e-06, 4.241682e-06, 4.04752e-06, 4.58443e-06, 4.452121e-06, 
    4.512834e-06, 4.579731e-06, 4.374315e-06, 4.156687e-06, 4.15217e-06, 
    4.084243e-06, 3.895093e-06, 4.222289e-06, 3.245661e-06, 3.836103e-06, 
    4.793475e-06, 4.591271e-06, 4.562636e-06, 4.640496e-06, 4.118761e-06, 
    4.306741e-06, 3.812347e-06, 3.942931e-06, 3.729919e-06, 3.835165e-06, 
    3.850749e-06, 3.987885e-06, 4.074198e-06, 4.298154e-06, 4.48177e-06, 
    4.629181e-06, 4.594769e-06, 4.433324e-06, 4.143698e-06, 3.879427e-06, 
    3.936736e-06, 3.745937e-06, 4.26167e-06, 4.040751e-06, 4.124582e-06, 
    3.907387e-06, 4.392129e-06, 3.977471e-06, 4.499965e-06, 4.453417e-06, 
    4.310459e-06, 4.026091e-06, 3.964814e-06, 3.899752e-06, 3.939854e-06, 
    4.136524e-06, 4.169097e-06, 4.31392e-06, 4.353536e-06, 4.46354e-06, 
    4.555286e-06, 4.471431e-06, 4.383918e-06, 4.13645e-06, 3.920733e-06, 
    3.690808e-06, 3.635438e-06, 3.376128e-06, 3.586536e-06, 3.242497e-06, 
    3.533931e-06, 3.03723e-06, 3.954126e-06, 3.542722e-06, 4.304e-06, 
    4.216728e-06, 4.065587e-06, 3.727086e-06, 3.908398e-06, 3.69672e-06, 
    4.170377e-06, 4.427776e-06, 4.494624e-06, 4.620171e-06, 4.491767e-06, 
    4.502167e-06, 4.380322e-06, 4.419358e-06, 4.128426e-06, 4.284875e-06, 
    3.851135e-06, 3.698378e-06, 3.281747e-06, 3.038143e-06, 2.800344e-06, 
    2.698797e-06, 2.668325e-06, 2.655646e-06,
  8.252843e-06, 8.083784e-06, 8.116454e-06, 7.981572e-06, 8.056179e-06, 
    7.968172e-06, 8.218372e-06, 8.077121e-06, 8.167091e-06, 8.237527e-06, 
    7.725238e-06, 7.975597e-06, 7.473606e-06, 7.627021e-06, 6.964885e-06, 
    7.497236e-06, 6.926678e-06, 6.97039e-06, 6.840516e-06, 6.877205e-06, 
    6.716742e-06, 6.823726e-06, 6.637081e-06, 6.74193e-06, 6.725249e-06, 
    6.827322e-06, 7.924645e-06, 7.756001e-06, 7.934737e-06, 7.910461e-06, 
    7.921348e-06, 8.05463e-06, 8.12246e-06, 8.265868e-06, 8.239705e-06, 
    8.134439e-06, 7.899566e-06, 7.978677e-06, 7.780643e-06, 7.785065e-06, 
    7.570066e-06, 7.666224e-06, 7.016791e-06, 7.09373e-06, 6.875665e-06, 
    6.929261e-06, 6.878162e-06, 6.893575e-06, 6.877962e-06, 6.956913e-06, 
    6.922861e-06, 6.993156e-06, 7.648113e-06, 7.53913e-06, 7.869035e-06, 
    8.073825e-06, 8.21214e-06, 8.311275e-06, 8.297213e-06, 8.270446e-06, 
    8.133825e-06, 8.006883e-06, 7.91121e-06, 7.847761e-06, 7.7857e-06, 
    7.600778e-06, 7.50485e-06, 7.001417e-06, 7.030681e-06, 6.981243e-06, 
    6.93464e-06, 6.857795e-06, 6.870321e-06, 6.836904e-06, 6.982542e-06, 
    6.885043e-06, 7.047452e-06, 7.002299e-06, 7.768888e-06, 7.95727e-06, 
    8.038507e-06, 8.110165e-06, 8.286411e-06, 8.164415e-06, 8.212359e-06, 
    8.09863e-06, 8.026971e-06, 8.062352e-06, 7.846033e-06, 7.929541e-06, 
    7.499209e-06, 7.68155e-06, 6.940043e-06, 7.024656e-06, 6.92006e-06, 
    6.973053e-06, 6.882747e-06, 6.963915e-06, 6.824559e-06, 6.795005e-06, 
    6.815169e-06, 6.738464e-06, 6.968471e-06, 6.878161e-06, 8.063344e-06, 
    8.057565e-06, 8.030685e-06, 8.149354e-06, 8.156656e-06, 8.266586e-06, 
    8.168721e-06, 8.127293e-06, 8.022834e-06, 7.961542e-06, 7.903641e-06, 
    7.777649e-06, 7.639236e-06, 7.450189e-06, 7.019112e-06, 6.950875e-06, 
    6.992566e-06, 6.955733e-06, 6.996932e-06, 7.016404e-06, 6.806044e-06, 
    6.922545e-06, 6.749371e-06, 6.758698e-06, 6.836113e-06, 6.757645e-06, 
    8.053509e-06, 8.086797e-06, 8.203153e-06, 8.111991e-06, 8.278616e-06, 
    8.185054e-06, 8.131588e-06, 7.927783e-06, 7.883578e-06, 7.842777e-06, 
    7.762774e-06, 7.66127e-06, 7.486653e-06, 7.035389e-06, 6.931948e-06, 
    6.939426e-06, 6.936792e-06, 6.914058e-06, 6.970644e-06, 6.904856e-06, 
    6.893938e-06, 6.92256e-06, 6.759949e-06, 6.805535e-06, 6.758896e-06, 
    6.788486e-06, 8.075966e-06, 8.020074e-06, 8.050238e-06, 7.993591e-06, 
    8.033464e-06, 7.85742e-06, 7.805304e-06, 7.565963e-06, 7.663253e-06, 
    7.509078e-06, 7.647435e-06, 7.622712e-06, 7.504101e-06, 7.639887e-06, 
    7.041727e-06, 7.543958e-06, 6.913177e-06, 7.063315e-06, 6.903977e-06, 
    6.932389e-06, 6.885479e-06, 6.844027e-06, 6.792651e-06, 6.700176e-06, 
    6.721317e-06, 6.645767e-06, 7.937331e-06, 7.865928e-06, 7.872196e-06, 
    7.798039e-06, 7.743621e-06, 7.626984e-06, 7.443958e-06, 7.512171e-06, 
    7.07388e-06, 7.054436e-06, 7.552403e-06, 7.435297e-06, 7.818466e-06, 
    7.755171e-06, 7.7928e-06, 7.931676e-06, 7.496379e-06, 7.716651e-06, 
    7.017414e-06, 7.430695e-06, 6.849904e-06, 6.975885e-06, 6.733025e-06, 
    6.635112e-06, 6.546438e-06, 6.447261e-06, 7.827205e-06, 7.875446e-06, 
    7.789266e-06, 7.67152e-06, 7.563947e-06, 7.423617e-06, 7.09113e-06, 
    7.07076e-06, 7.018486e-06, 6.975088e-06, 7.064338e-06, 6.96429e-06, 
    7.740556e-06, 7.477603e-06, 7.893752e-06, 7.766009e-06, 7.678412e-06, 
    7.716719e-06, 7.520016e-06, 7.47449e-06, 6.999559e-06, 7.07276e-06, 
    6.65893e-06, 6.835337e-06, 6.375122e-06, 6.494257e-06, 7.892364e-06, 
    7.827372e-06, 7.605188e-06, 7.710095e-06, 7.095007e-06, 7.039376e-06, 
    6.994739e-06, 6.938456e-06, 6.932436e-06, 6.89957e-06, 6.953592e-06, 
    6.901688e-06, 7.423322e-06, 7.011178e-06, 7.630254e-06, 7.550221e-06, 
    7.586923e-06, 7.627409e-06, 7.503239e-06, 7.062916e-06, 7.060765e-06, 
    7.028562e-06, 6.93928e-06, 7.094086e-06, 6.636982e-06, 6.911541e-06, 
    7.757069e-06, 7.634408e-06, 7.617062e-06, 7.664223e-06, 7.044918e-06, 
    7.462498e-06, 6.900367e-06, 6.96179e-06, 6.861731e-06, 6.91108e-06, 
    6.918403e-06, 6.982996e-06, 7.023804e-06, 7.457325e-06, 7.568141e-06, 
    7.657364e-06, 7.636516e-06, 7.538867e-06, 7.05675e-06, 6.931888e-06, 
    6.958874e-06, 6.869231e-06, 7.435351e-06, 7.00798e-06, 7.047681e-06, 
    6.945045e-06, 7.513992e-06, 6.978101e-06, 7.579139e-06, 7.551002e-06, 
    7.464738e-06, 7.001052e-06, 6.972109e-06, 6.941453e-06, 6.960339e-06, 
    7.053345e-06, 7.068804e-06, 7.466822e-06, 7.490709e-06, 7.557118e-06, 
    7.61261e-06, 7.56189e-06, 7.509039e-06, 7.053307e-06, 6.951333e-06, 
    6.84344e-06, 6.81758e-06, 6.697152e-06, 6.794794e-06, 6.635527e-06, 
    6.770329e-06, 6.541447e-06, 6.96708e-06, 6.774404e-06, 7.460844e-06, 
    7.09144e-06, 7.019733e-06, 6.860414e-06, 6.945521e-06, 6.846208e-06, 
    7.069411e-06, 7.53552e-06, 7.57591e-06, 7.651905e-06, 7.574182e-06, 
    7.580471e-06, 7.506864e-06, 7.530427e-06, 7.049501e-06, 7.449323e-06, 
    6.918586e-06, 6.846982e-06, 6.65358e-06, 6.541855e-06, 6.433843e-06, 
    6.38807e-06, 6.374378e-06, 6.368688e-06,
  9.622186e-06, 9.637707e-06, 9.634876e-06, 9.646008e-06, 9.640034e-06, 
    9.647031e-06, 9.625523e-06, 9.638273e-06, 9.630326e-06, 9.623679e-06, 
    9.662735e-06, 9.646466e-06, 9.672489e-06, 9.667408e-06, 1.000887e-05, 
    9.671892e-06, 9.993944e-06, 1.0011e-05, 9.959222e-06, 9.974196e-06, 
    9.906439e-06, 9.952271e-06, 9.870403e-06, 9.917483e-06, 9.910188e-06, 
    9.953765e-06, 9.65025e-06, 9.661062e-06, 9.649519e-06, 9.651261e-06, 
    9.650486e-06, 9.640162e-06, 9.634345e-06, 9.620905e-06, 9.623468e-06, 
    9.633281e-06, 9.652026e-06, 9.646232e-06, 9.659659e-06, 9.659399e-06, 
    9.669624e-06, 9.665671e-06, 1.002872e-05, 1.005728e-05, 9.973573e-06, 
    9.994965e-06, 9.974582e-06, 9.980786e-06, 9.974501e-06, 1.000578e-05, 
    9.99244e-06, 1.001974e-05, 9.666494e-06, 9.670667e-06, 9.654113e-06, 
    9.63855e-06, 9.626116e-06, 9.616344e-06, 9.617771e-06, 9.62045e-06, 
    9.633336e-06, 9.644034e-06, 9.651209e-06, 9.655517e-06, 9.659362e-06, 
    9.668472e-06, 9.671686e-06, 1.002289e-05, 1.003395e-05, 1.001518e-05, 
    9.99708e-06, 9.966308e-06, 9.971408e-06, 9.957731e-06, 1.001568e-05, 
    9.977356e-06, 1.004022e-05, 1.002323e-05, 9.660333e-06, 9.647854e-06, 
    9.641488e-06, 9.635427e-06, 9.618859e-06, 9.63057e-06, 9.626095e-06, 
    9.636431e-06, 9.642428e-06, 9.639519e-06, 9.655629e-06, 9.649897e-06, 
    9.67184e-06, 9.664945e-06, 9.9992e-06, 1.003168e-05, 9.991333e-06, 
    1.001203e-05, 9.976432e-06, 1.00085e-05, 9.952617e-06, 9.940234e-06, 
    9.948704e-06, 9.915975e-06, 1.001026e-05, 9.974581e-06, 9.639436e-06, 
    9.639918e-06, 9.642128e-06, 9.631941e-06, 9.631279e-06, 9.620834e-06, 
    9.630176e-06, 9.633918e-06, 9.642762e-06, 9.647533e-06, 9.651742e-06, 
    9.659832e-06, 9.666885e-06, 9.673009e-06, 1.002959e-05, 1.000343e-05, 
    1.001952e-05, 1.000532e-05, 1.002118e-05, 1.002857e-05, 9.944883e-06, 
    9.992315e-06, 9.920715e-06, 9.924746e-06, 9.957404e-06, 9.924292e-06, 
    9.640255e-06, 9.637451e-06, 9.626968e-06, 9.635268e-06, 9.619638e-06, 
    9.628665e-06, 9.633535e-06, 9.650023e-06, 9.653131e-06, 9.655839e-06, 
    9.660686e-06, 9.665901e-06, 9.67217e-06, 1.003571e-05, 9.996023e-06, 
    9.998959e-06, 9.997926e-06, 9.988955e-06, 1.00111e-05, 9.985296e-06, 
    9.98093e-06, 9.992322e-06, 9.925286e-06, 9.944671e-06, 9.924832e-06, 
    9.937478e-06, 9.638373e-06, 9.642983e-06, 9.640527e-06, 9.645078e-06, 
    9.641902e-06, 9.654883e-06, 9.658185e-06, 9.669767e-06, 9.665809e-06, 
    9.671569e-06, 9.666525e-06, 9.667589e-06, 9.671705e-06, 9.666858e-06, 
    1.003808e-05, 9.67051e-06, 9.988606e-06, 1.00461e-05, 9.984945e-06, 
    9.996196e-06, 9.977534e-06, 9.960666e-06, 9.939241e-06, 9.89909e-06, 
    9.908461e-06, 9.874421e-06, 9.64933e-06, 9.654321e-06, 9.653902e-06, 
    9.658627e-06, 9.661752e-06, 9.667411e-06, 9.673136e-06, 9.671483e-06, 
    1.005001e-05, 1.004282e-05, 9.670234e-06, 9.673303e-06, 9.657378e-06, 
    9.661112e-06, 9.65894e-06, 9.649741e-06, 9.671917e-06, 9.663187e-06, 
    1.002895e-05, 9.673388e-06, 9.96308e-06, 1.001312e-05, 9.9136e-06, 
    9.869486e-06, 9.827098e-06, 9.776424e-06, 9.656831e-06, 9.653683e-06, 
    9.659151e-06, 9.665421e-06, 9.66984e-06, 9.673513e-06, 1.005633e-05, 
    1.004886e-05, 1.002936e-05, 1.001281e-05, 1.004648e-05, 1.000864e-05, 
    9.661915e-06, 9.672394e-06, 9.652431e-06, 9.6605e-06, 9.665096e-06, 
    9.663186e-06, 9.671256e-06, 9.672471e-06, 1.002218e-05, 1.004959e-05, 
    9.88046e-06, 9.957081e-06, 9.737024e-06, 9.800901e-06, 9.652527e-06, 
    9.656821e-06, 9.668302e-06, 9.663528e-06, 1.005775e-05, 1.003721e-05, 
    1.002035e-05, 9.998577e-06, 9.996214e-06, 9.983185e-06, 1.000449e-05, 
    9.984032e-06, 9.673518e-06, 1.00266e-05, 9.667273e-06, 9.670306e-06, 
    9.669008e-06, 9.667393e-06, 9.671733e-06, 1.004596e-05, 1.004516e-05, 
    1.003315e-05, 9.99889e-06, 1.005741e-05, 9.870347e-06, 9.987946e-06, 
    9.661008e-06, 9.667093e-06, 9.667823e-06, 9.665764e-06, 1.003927e-05, 
    9.672746e-06, 9.983504e-06, 1.000767e-05, 9.967916e-06, 9.987773e-06, 
    9.990677e-06, 1.001585e-05, 1.003136e-05, 9.672859e-06, 9.669692e-06, 
    9.66608e-06, 9.667005e-06, 9.670675e-06, 1.004367e-05, 9.995998e-06, 
    1.000654e-05, 9.970966e-06, 9.673303e-06, 1.002538e-05, 1.00403e-05, 
    1.000116e-05, 9.67143e-06, 1.001396e-05, 9.669297e-06, 9.670282e-06, 
    9.672696e-06, 1.002275e-05, 1.001166e-05, 9.999751e-06, 1.000711e-05, 
    1.004241e-05, 1.004813e-05, 9.672649e-06, 9.672067e-06, 9.670075e-06, 
    9.668005e-06, 9.669911e-06, 9.67157e-06, 1.00424e-05, 1.000361e-05, 
    9.960424e-06, 9.949712e-06, 9.897735e-06, 9.940141e-06, 9.869671e-06, 
    9.929729e-06, 9.824626e-06, 1.000972e-05, 9.931479e-06, 9.672784e-06, 
    1.005644e-05, 1.002983e-05, 9.967374e-06, 1.000134e-05, 9.96156e-06, 
    1.004836e-05, 9.67078e-06, 9.669415e-06, 9.666326e-06, 9.669478e-06, 
    9.669248e-06, 9.671633e-06, 9.670941e-06, 1.004098e-05, 9.673029e-06, 
    9.990749e-06, 9.961878e-06, 9.878014e-06, 9.824833e-06, 9.769275e-06, 
    9.744274e-06, 9.736606e-06, 9.733393e-06,
  4.406781e-06, 4.320459e-06, 4.337229e-06, 4.267696e-06, 4.306256e-06, 
    4.260744e-06, 4.389271e-06, 4.317032e-06, 4.363137e-06, 4.399009e-06, 
    4.133104e-06, 4.264597e-06, 3.997111e-06, 4.080551e-06, 3.871728e-06, 
    4.010074e-06, 3.843862e-06, 3.875726e-06, 3.779978e-06, 3.807367e-06, 
    3.685346e-06, 3.767349e-06, 3.622404e-06, 3.704904e-06, 3.691971e-06, 
    3.770059e-06, 4.238105e-06, 4.149445e-06, 4.243363e-06, 4.230706e-06, 
    4.236386e-06, 4.305457e-06, 4.340302e-06, 4.413391e-06, 4.400115e-06, 
    4.34644e-06, 4.225015e-06, 4.266199e-06, 4.162512e-06, 4.16485e-06, 
    4.049776e-06, 4.101608e-06, 3.909171e-06, 3.963829e-06, 3.806223e-06, 
    3.845759e-06, 3.808077e-06, 3.819498e-06, 3.807929e-06, 3.865941e-06, 
    3.841067e-06, 3.892183e-06, 4.091892e-06, 4.032961e-06, 4.209041e-06, 
    4.31533e-06, 4.386099e-06, 4.436374e-06, 4.429263e-06, 4.41571e-06, 
    4.346126e-06, 4.280809e-06, 4.2311e-06, 4.197884e-06, 4.165187e-06, 
    4.066389e-06, 4.014245e-06, 3.898128e-06, 3.919111e-06, 3.883581e-06, 
    3.849696e-06, 3.792911e-06, 3.802249e-06, 3.777265e-06, 3.884523e-06, 
    3.813179e-06, 3.93107e-06, 3.898766e-06, 4.156273e-06, 4.255085e-06, 
    4.297137e-06, 4.334004e-06, 4.423796e-06, 4.361767e-06, 4.38621e-06, 
    4.328088e-06, 4.291192e-06, 4.309437e-06, 4.196976e-06, 4.240658e-06, 
    4.011158e-06, 4.10981e-06, 3.853646e-06, 3.914804e-06, 3.839012e-06, 
    3.877658e-06, 3.811478e-06, 3.871031e-06, 3.767976e-06, 3.745597e-06, 
    3.760887e-06, 3.702227e-06, 3.874336e-06, 3.808075e-06, 4.309947e-06, 
    4.306971e-06, 4.29311e-06, 4.35407e-06, 4.357804e-06, 4.413754e-06, 
    4.363969e-06, 4.342783e-06, 4.289057e-06, 4.257305e-06, 4.227147e-06, 
    4.160927e-06, 4.08712e-06, 3.984222e-06, 3.910834e-06, 3.861548e-06, 
    3.89176e-06, 3.865085e-06, 3.894905e-06, 3.908896e-06, 3.753978e-06, 
    3.840833e-06, 3.710654e-06, 3.717837e-06, 3.77667e-06, 3.717027e-06, 
    4.304881e-06, 4.322011e-06, 4.381525e-06, 4.334943e-06, 4.419851e-06, 
    4.372301e-06, 4.34498e-06, 4.239738e-06, 4.21666e-06, 4.195264e-06, 
    4.153052e-06, 4.098953e-06, 4.004279e-06, 3.92247e-06, 3.847728e-06, 
    3.853197e-06, 3.851271e-06, 3.834601e-06, 3.875912e-06, 3.827827e-06, 
    3.819764e-06, 3.840847e-06, 3.718799e-06, 3.753596e-06, 3.71799e-06, 
    3.740639e-06, 4.316443e-06, 4.287629e-06, 4.303196e-06, 4.273927e-06, 
    4.294543e-06, 4.202948e-06, 4.17553e-06, 4.047545e-06, 4.100015e-06, 
    4.016561e-06, 4.09153e-06, 4.07823e-06, 4.01383e-06, 4.087476e-06, 
    3.926986e-06, 4.035584e-06, 3.833954e-06, 3.942325e-06, 3.827178e-06, 
    3.848051e-06, 3.813506e-06, 3.78261e-06, 3.74381e-06, 3.672404e-06, 
    3.688917e-06, 3.629357e-06, 4.244715e-06, 4.207412e-06, 4.2107e-06, 
    4.171704e-06, 4.14289e-06, 4.080533e-06, 3.980786e-06, 4.018256e-06, 
    3.94982e-06, 3.936034e-06, 4.040187e-06, 3.976e-06, 4.182472e-06, 
    4.149015e-06, 4.168935e-06, 4.241768e-06, 4.009609e-06, 4.128542e-06, 
    3.909617e-06, 3.973458e-06, 3.787012e-06, 3.879703e-06, 3.698012e-06, 
    3.62082e-06, 3.548496e-06, 3.464337e-06, 4.187075e-06, 4.212403e-06, 
    4.167071e-06, 4.10444e-06, 4.046457e-06, 3.969541e-06, 3.961998e-06, 
    3.94761e-06, 3.910387e-06, 3.879131e-06, 3.943057e-06, 3.871303e-06, 
    4.14125e-06, 3.999311e-06, 4.221979e-06, 4.154759e-06, 4.108131e-06, 
    4.128583e-06, 4.022543e-06, 3.997604e-06, 3.896792e-06, 3.949027e-06, 
    3.639837e-06, 3.776082e-06, 3.400579e-06, 3.504681e-06, 4.221255e-06, 
    4.187165e-06, 4.068778e-06, 4.125054e-06, 3.964729e-06, 3.925315e-06, 
    3.893325e-06, 3.852485e-06, 3.848084e-06, 3.823925e-06, 3.863526e-06, 
    3.825491e-06, 3.969377e-06, 3.905146e-06, 4.082295e-06, 4.038999e-06, 
    4.058911e-06, 4.080763e-06, 4.013371e-06, 3.942048e-06, 3.940529e-06, 
    3.917594e-06, 3.853067e-06, 3.96408e-06, 3.622305e-06, 3.832731e-06, 
    4.150029e-06, 4.084522e-06, 4.075187e-06, 4.100537e-06, 3.929264e-06, 
    3.991007e-06, 3.824515e-06, 3.869488e-06, 3.79585e-06, 3.832411e-06, 
    3.837795e-06, 3.884852e-06, 3.914194e-06, 3.988157e-06, 4.048732e-06, 
    4.09686e-06, 4.085663e-06, 4.032819e-06, 3.937674e-06, 3.847681e-06, 
    3.867364e-06, 3.801438e-06, 3.976033e-06, 3.902847e-06, 3.931228e-06, 
    3.857298e-06, 4.01925e-06, 3.881293e-06, 4.054697e-06, 4.039426e-06, 
    3.99224e-06, 3.897863e-06, 3.876974e-06, 3.854674e-06, 3.868434e-06, 
    3.935256e-06, 3.946225e-06, 3.993388e-06, 4.006505e-06, 4.04275e-06, 
    4.072789e-06, 4.045341e-06, 4.016541e-06, 3.935232e-06, 3.861878e-06, 
    3.782169e-06, 3.762711e-06, 3.670022e-06, 3.745429e-06, 3.621138e-06, 
    3.72674e-06, 3.544331e-06, 3.873316e-06, 3.729872e-06, 3.990098e-06, 
    3.962216e-06, 3.911274e-06, 3.794859e-06, 3.857645e-06, 3.78424e-06, 
    3.946655e-06, 4.030993e-06, 4.052946e-06, 4.09393e-06, 4.05201e-06, 
    4.055418e-06, 4.015355e-06, 4.028224e-06, 3.932525e-06, 3.983749e-06, 
    3.837928e-06, 3.784821e-06, 3.635587e-06, 3.544681e-06, 3.452662e-06, 
    3.412204e-06, 3.399912e-06, 3.394776e-06,
  4.550292e-07, 4.380054e-07, 4.412852e-07, 4.27773e-07, 4.352383e-07, 
    4.264347e-07, 4.515475e-07, 4.373368e-07, 4.46378e-07, 4.53482e-07, 
    4.022619e-07, 4.271762e-07, 3.773407e-07, 3.925299e-07, 3.550694e-07, 
    3.796794e-07, 3.502303e-07, 3.557667e-07, 3.392699e-07, 3.439463e-07, 
    3.233738e-07, 3.371251e-07, 3.130245e-07, 3.26626e-07, 3.244735e-07, 
    3.375847e-07, 4.220917e-07, 4.053142e-07, 4.230982e-07, 4.206774e-07, 
    4.21763e-07, 4.350827e-07, 4.418876e-07, 4.563473e-07, 4.537021e-07, 
    4.430923e-07, 4.195916e-07, 4.274846e-07, 4.07764e-07, 4.082032e-07, 
    3.868902e-07, 3.96414e-07, 3.616274e-07, 3.71316e-07, 3.437503e-07, 
    3.505588e-07, 3.44068e-07, 3.460284e-07, 3.440425e-07, 3.540617e-07, 
    3.49747e-07, 3.586443e-07, 3.946193e-07, 3.838275e-07, 4.165514e-07, 
    4.370052e-07, 4.509183e-07, 4.609465e-07, 4.595209e-07, 4.568101e-07, 
    4.430306e-07, 4.303039e-07, 4.207527e-07, 4.14435e-07, 4.082663e-07, 
    3.899291e-07, 3.804335e-07, 3.596867e-07, 3.633793e-07, 3.571385e-07, 
    3.512407e-07, 3.414738e-07, 3.430698e-07, 3.388085e-07, 3.573033e-07, 
    3.44943e-07, 3.654928e-07, 3.597988e-07, 4.065932e-07, 4.253468e-07, 
    4.334666e-07, 4.406534e-07, 4.584264e-07, 4.461081e-07, 4.509403e-07, 
    4.394959e-07, 4.323135e-07, 4.358572e-07, 4.14263e-07, 4.225802e-07, 
    3.798752e-07, 3.979325e-07, 3.519255e-07, 3.626196e-07, 3.493918e-07, 
    3.561039e-07, 3.446511e-07, 3.549481e-07, 3.372314e-07, 3.334479e-07, 
    3.360304e-07, 3.261798e-07, 3.555243e-07, 3.440675e-07, 4.359565e-07, 
    4.353773e-07, 4.326854e-07, 4.445922e-07, 4.453272e-07, 4.564197e-07, 
    4.465422e-07, 4.423742e-07, 4.318998e-07, 4.257733e-07, 4.199981e-07, 
    4.074664e-07, 3.937394e-07, 3.750229e-07, 3.619203e-07, 3.532976e-07, 
    3.5857e-07, 3.539126e-07, 3.591213e-07, 3.615791e-07, 3.348621e-07, 
    3.497066e-07, 3.275853e-07, 3.287859e-07, 3.387073e-07, 3.286505e-07, 
    4.349709e-07, 4.383084e-07, 4.500119e-07, 4.408374e-07, 4.576374e-07, 
    4.481871e-07, 4.428055e-07, 4.224041e-07, 4.179998e-07, 4.139389e-07, 
    4.059896e-07, 3.959231e-07, 3.786329e-07, 3.639722e-07, 3.508997e-07, 
    3.518475e-07, 3.515136e-07, 3.4863e-07, 3.557991e-07, 3.474618e-07, 
    3.46074e-07, 3.49709e-07, 3.289469e-07, 3.347975e-07, 3.288115e-07, 
    3.326126e-07, 4.37222e-07, 4.316234e-07, 4.346433e-07, 4.289746e-07, 
    4.329632e-07, 4.153949e-07, 4.102123e-07, 3.864832e-07, 3.961195e-07, 
    3.808526e-07, 3.945524e-07, 3.921031e-07, 3.803584e-07, 3.938049e-07, 
    3.647702e-07, 3.843043e-07, 3.485183e-07, 3.67488e-07, 3.473501e-07, 
    3.509556e-07, 3.449992e-07, 3.397178e-07, 3.331467e-07, 3.212311e-07, 
    3.239663e-07, 3.141589e-07, 4.233573e-07, 4.16242e-07, 4.168666e-07, 
    4.094919e-07, 4.040885e-07, 3.925268e-07, 3.744064e-07, 3.811594e-07, 
    3.688197e-07, 3.663721e-07, 3.851421e-07, 3.735485e-07, 4.115212e-07, 
    4.052338e-07, 4.089711e-07, 4.227927e-07, 3.795953e-07, 4.014121e-07, 
    3.61706e-07, 3.730933e-07, 3.404676e-07, 3.564609e-07, 3.254779e-07, 
    3.127663e-07, 3.01099e-07, 2.878165e-07, 4.123903e-07, 4.171903e-07, 
    4.086204e-07, 3.96938e-07, 3.862845e-07, 3.723923e-07, 3.709891e-07, 
    3.684268e-07, 3.618417e-07, 3.563611e-07, 3.676179e-07, 3.549955e-07, 
    4.037819e-07, 3.77737e-07, 4.190127e-07, 4.063095e-07, 3.976214e-07, 
    4.014197e-07, 3.819362e-07, 3.774296e-07, 3.594522e-07, 3.686787e-07, 
    3.158731e-07, 3.386074e-07, 2.779633e-07, 2.941445e-07, 4.188749e-07, 
    4.124073e-07, 3.903674e-07, 4.007629e-07, 3.714766e-07, 3.64475e-07, 
    3.588444e-07, 3.51724e-07, 3.509613e-07, 3.4679e-07, 3.536416e-07, 
    3.470594e-07, 3.723631e-07, 3.609195e-07, 3.928508e-07, 3.849257e-07, 
    3.885597e-07, 3.92569e-07, 3.802755e-07, 3.674387e-07, 3.671691e-07, 
    3.631117e-07, 3.518248e-07, 3.713607e-07, 3.130084e-07, 3.483072e-07, 
    4.054235e-07, 3.932607e-07, 3.915438e-07, 3.96216e-07, 3.651732e-07, 
    3.762421e-07, 3.468915e-07, 3.546792e-07, 3.419758e-07, 3.482522e-07, 
    3.491815e-07, 3.573608e-07, 3.625121e-07, 3.757298e-07, 3.866997e-07, 
    3.955365e-07, 3.93471e-07, 3.838015e-07, 3.666627e-07, 3.508916e-07, 
    3.543094e-07, 3.429311e-07, 3.735545e-07, 3.605154e-07, 3.655207e-07, 
    3.525591e-07, 3.813395e-07, 3.567386e-07, 3.87789e-07, 3.850034e-07, 
    3.764639e-07, 3.596402e-07, 3.559845e-07, 3.521037e-07, 3.544956e-07, 
    3.662342e-07, 3.681806e-07, 3.766704e-07, 3.790346e-07, 3.85609e-07, 
    3.911033e-07, 3.86081e-07, 3.808489e-07, 3.662298e-07, 3.53355e-07, 
    3.396428e-07, 3.363391e-07, 3.208376e-07, 3.334195e-07, 3.128181e-07, 
    3.302771e-07, 3.004342e-07, 3.553463e-07, 3.308028e-07, 3.760786e-07, 
    3.710282e-07, 3.619978e-07, 3.418065e-07, 3.526194e-07, 3.399952e-07, 
    3.682571e-07, 3.834697e-07, 3.874692e-07, 3.949955e-07, 3.872982e-07, 
    3.879209e-07, 3.806343e-07, 3.829668e-07, 3.657505e-07, 3.74938e-07, 
    3.492044e-07, 3.400942e-07, 3.151773e-07, 3.0049e-07, 2.859987e-07, 
    2.797463e-07, 2.778611e-07, 2.770755e-07,
  1.281292e-08, 1.207718e-08, 1.221775e-08, 1.164228e-08, 1.195902e-08, 
    1.15858e-08, 1.266122e-08, 1.204859e-08, 1.243714e-08, 1.274543e-08, 
    1.058242e-08, 1.161708e-08, 9.581546e-09, 1.018746e-08, 8.716812e-09, 
    9.673996e-09, 8.532719e-09, 8.743454e-09, 8.120853e-09, 8.295709e-09, 
    7.536279e-09, 8.04109e-09, 7.169221e-09, 7.654631e-09, 7.576226e-09, 
    8.058158e-09, 1.140321e-08, 1.070737e-08, 1.144544e-08, 1.134397e-08, 
    1.138943e-08, 1.195239e-08, 1.224362e-08, 1.287051e-08, 1.275502e-08, 
    1.229544e-08, 1.129855e-08, 1.16301e-08, 1.080802e-08, 1.08261e-08, 
    9.960978e-09, 1.034446e-08, 8.968478e-09, 9.344821e-09, 8.288356e-09, 
    8.545171e-09, 8.300279e-09, 8.373981e-09, 8.299321e-09, 8.678362e-09, 
    8.514407e-09, 8.853688e-09, 1.027181e-08, 9.838726e-09, 1.117175e-08, 
    1.203442e-08, 1.263387e-08, 1.307218e-08, 1.300955e-08, 1.289076e-08, 
    1.229278e-08, 1.174933e-08, 1.134712e-08, 1.108376e-08, 1.08287e-08, 
    1.008279e-08, 9.703873e-09, 8.893742e-09, 9.036128e-09, 8.795944e-09, 
    8.571044e-09, 8.203099e-09, 8.262838e-09, 8.103668e-09, 8.802258e-09, 
    8.333145e-09, 9.117977e-09, 8.898053e-09, 1.075988e-08, 1.153997e-08, 
    1.188358e-08, 1.219062e-08, 1.296154e-08, 1.242547e-08, 1.263483e-08, 
    1.214099e-08, 1.183457e-08, 1.198541e-08, 1.107662e-08, 1.14237e-08, 
    9.68175e-09, 1.040607e-08, 8.597052e-09, 9.00677e-09, 8.500959e-09, 
    8.756345e-09, 8.322178e-09, 8.71218e-09, 8.045037e-09, 7.90498e-09, 
    8.000486e-09, 7.638356e-09, 8.734187e-09, 8.30026e-09, 1.198965e-08, 
    1.196495e-08, 1.185037e-08, 1.236005e-08, 1.239176e-08, 1.287368e-08, 
    1.244423e-08, 1.226454e-08, 1.181701e-08, 1.155793e-08, 1.131555e-08, 
    1.079578e-08, 1.023626e-08, 9.490232e-09, 8.979776e-09, 8.649248e-09, 
    8.850839e-09, 8.67268e-09, 8.872012e-09, 8.966614e-09, 7.95723e-09, 
    8.512878e-09, 7.689666e-09, 7.733592e-09, 8.099904e-09, 7.728634e-09, 
    1.194762e-08, 1.209014e-08, 1.259451e-08, 1.219852e-08, 1.292697e-08, 
    1.25154e-08, 1.228309e-08, 1.141631e-08, 1.12321e-08, 1.106317e-08, 
    1.073509e-08, 1.032457e-08, 9.63259e-09, 9.059061e-09, 8.558102e-09, 
    8.594091e-09, 8.581407e-09, 8.472142e-09, 8.74469e-09, 8.428014e-09, 
    8.3757e-09, 8.512968e-09, 7.739488e-09, 7.954841e-09, 7.734528e-09, 
    7.874178e-09, 1.204369e-08, 1.180528e-08, 1.193367e-08, 1.169306e-08, 
    1.186218e-08, 1.112364e-08, 1.090894e-08, 9.944698e-09, 1.033253e-08, 
    9.720487e-09, 1.026911e-08, 1.017026e-08, 9.700893e-09, 1.023891e-08, 
    9.089964e-09, 9.857725e-09, 8.467916e-09, 9.195479e-09, 8.423799e-09, 
    8.560223e-09, 8.335258e-09, 8.137542e-09, 7.893868e-09, 7.458658e-09, 
    7.557793e-09, 7.204457e-09, 1.145632e-08, 1.115887e-08, 1.118487e-08, 
    1.087921e-08, 1.065713e-08, 1.018733e-08, 9.465992e-09, 9.732662e-09, 
    9.247338e-09, 9.152105e-09, 9.891137e-09, 9.432301e-09, 1.096303e-08, 
    1.070407e-08, 1.085774e-08, 1.143262e-08, 9.670666e-09, 1.054772e-08, 
    8.971508e-09, 9.414442e-09, 8.165511e-09, 8.770003e-09, 7.61278e-09, 
    7.159988e-09, 6.747238e-09, 6.288079e-09, 1.099899e-08, 1.119835e-08, 
    1.084329e-08, 1.036571e-08, 9.936761e-09, 9.386961e-09, 9.332034e-09, 
    9.232028e-09, 8.976742e-09, 8.766185e-09, 9.200535e-09, 8.71399e-09, 
    1.064458e-08, 9.597192e-09, 1.127437e-08, 1.074822e-08, 1.039344e-08, 
    1.054804e-08, 9.763501e-09, 9.585055e-09, 8.884728e-09, 9.241843e-09, 
    7.265785e-09, 8.096183e-09, 5.954996e-09, 6.505391e-09, 1.126862e-08, 
    1.09997e-08, 1.01004e-08, 1.052125e-08, 9.351103e-09, 9.078527e-09, 
    8.861375e-09, 8.589399e-09, 8.560441e-09, 8.402674e-09, 8.662351e-09, 
    8.412834e-09, 9.385816e-09, 8.941192e-09, 1.02004e-08, 9.882503e-09, 
    1.002784e-08, 1.018903e-08, 9.69761e-09, 9.193564e-09, 9.183077e-09, 
    9.025782e-09, 8.593227e-09, 9.34657e-09, 7.168644e-09, 8.459939e-09, 
    1.071186e-08, 1.021693e-08, 1.014773e-08, 1.033644e-08, 9.105582e-09, 
    9.538227e-09, 8.406502e-09, 8.701917e-09, 8.221871e-09, 8.45786e-09, 
    8.493e-09, 8.804463e-09, 9.002617e-09, 9.518049e-09, 9.953357e-09, 
    1.030892e-08, 1.022542e-08, 9.837695e-09, 9.163394e-09, 8.557794e-09, 
    8.687809e-09, 8.257641e-09, 9.432536e-09, 8.925627e-09, 9.119059e-09, 
    8.621143e-09, 9.739808e-09, 8.780631e-09, 9.996954e-09, 9.885602e-09, 
    9.546968e-09, 8.891955e-09, 8.75178e-09, 8.603826e-09, 8.694911e-09, 
    9.146748e-09, 9.222437e-09, 9.55511e-09, 9.648478e-09, 9.909773e-09, 
    1.013e-08, 9.928629e-09, 9.720344e-09, 9.14658e-09, 8.651434e-09, 
    8.134745e-09, 8.011929e-09, 7.444432e-09, 7.903934e-09, 7.16184e-09, 
    7.788269e-09, 6.723985e-09, 8.727389e-09, 7.807577e-09, 9.531788e-09, 
    9.333562e-09, 8.982764e-09, 8.215536e-09, 8.623437e-09, 8.147888e-09, 
    9.225417e-09, 9.824481e-09, 9.984149e-09, 1.028703e-08, 9.977303e-09, 
    1.000224e-08, 9.711834e-09, 9.804468e-09, 9.127974e-09, 9.486893e-09, 
    8.493868e-09, 8.15158e-09, 7.24087e-09, 6.725935e-09, 6.226141e-09, 
    6.01479e-09, 5.951578e-09, 5.925303e-09,
  8.841755e-11, 8.066264e-11, 8.212646e-11, 7.618853e-11, 7.943888e-11, 
    7.561373e-11, 8.679991e-11, 8.036601e-11, 8.442805e-11, 8.769666e-11, 
    6.564504e-11, 7.593193e-11, 5.618734e-11, 6.185275e-11, 4.843886e-11, 
    5.703953e-11, 4.684305e-11, 4.86714e-11, 4.33444e-11, 4.481748e-11, 
    3.855547e-11, 4.267855e-11, 3.241819e-11, 3.950777e-11, 3.88759e-11, 
    4.282069e-11, 7.376501e-11, 6.686059e-11, 7.41912e-11, 7.316841e-11, 
    7.36261e-11, 7.937038e-11, 8.239685e-11, 8.903422e-11, 8.779902e-11, 
    8.293913e-11, 7.271221e-11, 7.606447e-11, 6.784524e-11, 6.802262e-11, 
    5.971315e-11, 6.335109e-11, 5.065152e-11, 5.402578e-11, 4.475517e-11, 
    4.695037e-11, 4.485622e-11, 4.548277e-11, 4.48481e-11, 4.810394e-11, 
    4.668538e-11, 4.963788e-11, 6.265626e-11, 5.856904e-11, 7.144332e-11, 
    8.02191e-11, 8.650929e-11, 9.120418e-11, 9.052852e-11, 8.925128e-11, 
    8.291133e-11, 7.728209e-11, 7.320012e-11, 7.056726e-11, 6.804816e-11, 
    6.086076e-11, 5.731589e-11, 4.999073e-11, 5.125236e-11, 4.913075e-11, 
    4.717366e-11, 4.4035e-11, 4.453916e-11, 4.320061e-11, 4.918611e-11, 
    4.513523e-11, 5.198265e-11, 5.002877e-11, 6.737369e-11, 7.514828e-11, 
    7.86607e-11, 8.184336e-11, 9.001166e-11, 8.430517e-11, 8.651944e-11, 
    8.132606e-11, 7.815653e-11, 7.971171e-11, 7.049635e-11, 7.397168e-11, 
    5.711121e-11, 6.394235e-11, 4.739851e-11, 5.099131e-11, 4.656972e-11, 
    4.878407e-11, 4.504205e-11, 4.839846e-11, 4.271139e-11, 4.155125e-11, 
    4.234106e-11, 3.937629e-11, 4.859047e-11, 4.485607e-11, 7.975551e-11, 
    7.950008e-11, 7.831893e-11, 8.361703e-11, 8.395028e-11, 8.906814e-11, 
    8.450282e-11, 8.261569e-11, 7.797607e-11, 7.533055e-11, 7.288285e-11, 
    6.772524e-11, 6.231717e-11, 5.535002e-11, 5.07517e-11, 4.785092e-11, 
    4.961281e-11, 4.805453e-11, 4.979918e-11, 5.063502e-11, 4.198264e-11, 
    4.667222e-11, 3.979138e-11, 4.014805e-11, 4.316914e-11, 4.010773e-11, 
    7.932115e-11, 8.079729e-11, 8.609159e-11, 8.192574e-11, 8.964007e-11, 
    8.5254e-11, 8.280985e-11, 7.389712e-11, 7.204631e-11, 7.036279e-11, 
    6.713129e-11, 6.31606e-11, 5.66573e-11, 5.14566e-11, 4.706192e-11, 
    4.737289e-11, 4.72632e-11, 4.632221e-11, 4.86822e-11, 4.594415e-11, 
    4.549743e-11, 4.6673e-11, 4.019602e-11, 4.196289e-11, 4.015566e-11, 
    4.129772e-11, 8.031515e-11, 7.785564e-11, 7.917706e-11, 7.670667e-11, 
    7.844037e-11, 7.096383e-11, 6.883733e-11, 5.956036e-11, 6.323676e-11, 
    5.746978e-11, 6.263044e-11, 6.168934e-11, 5.728831e-11, 6.234238e-11, 
    5.17323e-11, 5.874634e-11, 4.628596e-11, 5.267755e-11, 4.59081e-11, 
    4.708023e-11, 4.515319e-11, 4.348421e-11, 4.145971e-11, 3.793578e-11, 
    3.872791e-11, 3.593382e-11, 7.430113e-11, 7.131485e-11, 7.157429e-11, 
    6.854457e-11, 6.637099e-11, 6.185154e-11, 5.512849e-11, 5.758263e-11, 
    5.314436e-11, 5.228825e-11, 5.905859e-11, 5.48211e-11, 6.937101e-11, 
    6.682846e-11, 6.833337e-11, 7.40617e-11, 5.700876e-11, 6.530887e-11, 
    5.067839e-11, 5.46584e-11, 4.371888e-11, 4.890354e-11, 3.917e-11, 
    3.236422e-11, 2.996439e-11, 2.732573e-11, 6.972664e-11, 7.170893e-11, 
    6.819138e-11, 6.355475e-11, 5.94859e-11, 5.440838e-11, 5.390987e-11, 
    5.300639e-11, 5.072479e-11, 4.887014e-11, 5.2723e-11, 4.841424e-11, 
    6.624882e-11, 5.633125e-11, 7.246963e-11, 6.725968e-11, 6.382097e-11, 
    6.531189e-11, 5.786884e-11, 5.621961e-11, 4.991124e-11, 5.309483e-11, 
    3.641291e-11, 4.313805e-11, 2.54335e-11, 2.857034e-11, 7.241199e-11, 
    6.973361e-11, 6.102729e-11, 6.505269e-11, 5.408276e-11, 5.163021e-11, 
    4.970552e-11, 4.73323e-11, 4.708211e-11, 4.572757e-11, 4.796474e-11, 
    4.581436e-11, 5.439797e-11, 5.040992e-11, 6.197579e-11, 5.897785e-11, 
    6.034209e-11, 6.186773e-11, 5.725792e-11, 5.266035e-11, 5.256614e-11, 
    5.11603e-11, 4.736541e-11, 5.404164e-11, 3.241481e-11, 4.621755e-11, 
    6.690441e-11, 6.213313e-11, 6.147558e-11, 6.327421e-11, 5.187183e-11, 
    5.578957e-11, 4.576026e-11, 4.830901e-11, 4.41932e-11, 4.619973e-11, 
    4.650131e-11, 4.920545e-11, 5.095441e-11, 5.560463e-11, 5.964161e-11, 
    6.301081e-11, 6.221395e-11, 5.855941e-11, 5.238947e-11, 4.705926e-11, 
    4.818615e-11, 4.449522e-11, 5.482324e-11, 5.027228e-11, 5.199234e-11, 
    4.760713e-11, 5.764891e-11, 4.899658e-11, 6.00513e-11, 5.900683e-11, 
    5.586974e-11, 4.997497e-11, 4.874416e-11, 4.745713e-11, 4.8248e-11, 
    5.224024e-11, 5.292003e-11, 5.594448e-11, 5.680386e-11, 5.923301e-11, 
    6.13075e-11, 5.940966e-11, 5.746844e-11, 5.223874e-11, 4.786991e-11, 
    4.346076e-11, 4.243607e-11, 3.782263e-11, 4.154262e-11, 3.237504e-11, 
    4.059371e-11, 2.982996e-11, 4.853113e-11, 4.075154e-11, 5.573052e-11, 
    5.392372e-11, 5.07782e-11, 4.413979e-11, 4.7627e-11, 4.357096e-11, 
    5.294686e-11, 5.843621e-11, 5.993087e-11, 6.280153e-11, 5.986651e-11, 
    6.010099e-11, 5.738962e-11, 5.82498e-11, 5.207211e-11, 5.531948e-11, 
    4.650877e-11, 4.360193e-11, 3.621798e-11, 2.984123e-11, 2.697242e-11, 
    2.577177e-11, 2.541418e-11, 2.526575e-11,
  8.52261e-14, 7.269577e-14, 7.502897e-14, 6.566399e-14, 7.075727e-14, 
    6.477193e-14, 8.257873e-14, 7.222487e-14, 7.872836e-14, 8.404422e-14, 
    4.975651e-14, 6.526543e-14, 3.643888e-14, 4.429571e-14, 2.637756e-14, 
    3.759587e-14, 2.441931e-14, 2.666643e-14, 2.028255e-14, 2.199697e-14, 
    1.501375e-14, 1.952133e-14, 1.202253e-14, 1.602173e-14, 1.535058e-14, 
    1.96831e-14, 6.192115e-14, 5.153815e-14, 6.257585e-14, 6.100727e-14, 
    6.17081e-14, 7.064909e-14, 7.546162e-14, 8.623977e-14, 8.421183e-14, 
    7.633094e-14, 6.031049e-14, 6.547122e-14, 5.2992e-14, 5.325489e-14, 
    4.12839e-14, 4.64351e-14, 2.91609e-14, 3.354657e-14, 2.192362e-14, 
    2.454966e-14, 2.204261e-14, 2.27845e-14, 2.203304e-14, 2.596307e-14, 
    2.422816e-14, 2.787629e-14, 4.543997e-14, 3.969514e-14, 5.838193e-14, 
    7.199188e-14, 8.210493e-14, 8.982569e-14, 8.8706e-14, 8.659713e-14, 
    7.628631e-14, 6.736841e-14, 6.105577e-14, 5.70587e-14, 5.329275e-14, 
    4.289287e-14, 3.797305e-14, 2.832167e-14, 2.992971e-14, 2.723961e-14, 
    2.48215e-14, 2.108118e-14, 2.166993e-14, 2.011743e-14, 2.730891e-14, 
    2.237209e-14, 3.08714e-14, 2.83698e-14, 5.229457e-14, 6.405155e-14, 
    6.953044e-14, 7.457651e-14, 8.785139e-14, 7.852992e-14, 8.212146e-14, 
    7.375127e-14, 6.873806e-14, 7.118848e-14, 5.695191e-14, 6.223843e-14, 
    3.769361e-14, 4.728595e-14, 2.509608e-14, 2.959501e-14, 2.408821e-14, 
    2.680671e-14, 2.22619e-14, 2.632747e-14, 1.955867e-14, 1.825284e-14, 
    1.913886e-14, 1.588132e-14, 2.65658e-14, 2.204242e-14, 7.125776e-14, 
    7.085395e-14, 6.899308e-14, 7.742055e-14, 7.795738e-14, 8.629559e-14, 
    7.884915e-14, 7.581219e-14, 6.845491e-14, 6.433344e-14, 6.057091e-14, 
    5.28143e-14, 4.495621e-14, 3.531116e-14, 2.92887e-14, 2.565115e-14, 
    2.784473e-14, 2.590207e-14, 2.807966e-14, 2.913985e-14, 1.87352e-14, 
    2.421222e-14, 1.632591e-14, 1.671101e-14, 2.008135e-14, 1.666733e-14, 
    7.057138e-14, 7.290972e-14, 8.142492e-14, 7.470811e-14, 8.723798e-14, 
    8.006485e-14, 7.61235e-14, 6.212394e-14, 5.929666e-14, 5.675084e-14, 
    5.193692e-14, 4.616177e-14, 3.70758e-14, 3.019229e-14, 2.468535e-14, 
    2.506475e-14, 2.493074e-14, 2.378952e-14, 2.667988e-14, 2.333534e-14, 
    2.280194e-14, 2.421317e-14, 1.676302e-14, 1.871303e-14, 1.671926e-14, 
    1.797116e-14, 7.214419e-14, 6.82661e-14, 7.034399e-14, 6.647037e-14, 
    6.918391e-14, 5.765685e-14, 5.446619e-14, 4.107084e-14, 4.627101e-14, 
    3.818347e-14, 4.540309e-14, 4.406386e-14, 3.793536e-14, 4.499214e-14, 
    3.05477e-14, 3.994033e-14, 2.374586e-14, 3.177465e-14, 2.329217e-14, 
    2.470764e-14, 2.239335e-14, 2.044349e-14, 1.815099e-14, 1.436923e-14, 
    1.519473e-14, 1.235161e-14, 6.274495e-14, 5.818746e-14, 5.858033e-14, 
    5.403021e-14, 5.081878e-14, 4.4294e-14, 3.501433e-14, 3.833798e-14, 
    3.238528e-14, 3.126777e-14, 4.037306e-14, 3.460354e-14, 5.526303e-14, 
    5.149087e-14, 5.371617e-14, 6.237675e-14, 3.755394e-14, 4.926638e-14, 
    2.919516e-14, 3.438662e-14, 2.071447e-14, 2.695568e-14, 1.566183e-14, 
    1.195312e-14, 9.047568e-15, 6.281996e-15, 5.57955e-14, 5.878446e-14, 
    5.350529e-14, 4.672777e-14, 4.096711e-14, 3.405398e-14, 3.339324e-14, 
    3.220448e-14, 2.925436e-14, 2.6914e-14, 3.183396e-14, 2.634704e-14, 
    5.063964e-14, 3.663362e-14, 5.994072e-14, 5.212628e-14, 4.711098e-14, 
    4.927077e-14, 3.873054e-14, 3.648252e-14, 2.822117e-14, 3.232034e-14, 
    1.282519e-14, 2.004571e-14, 4.594181e-15, 7.528408e-15, 5.985292e-14, 
    5.580594e-14, 4.31276e-14, 4.889364e-14, 3.362201e-14, 3.041596e-14, 
    2.796152e-14, 2.501514e-14, 2.470994e-14, 2.307629e-14, 2.579133e-14, 
    2.318e-14, 3.404014e-14, 2.885327e-14, 4.447046e-14, 4.026105e-14, 
    4.216382e-14, 4.431697e-14, 3.789386e-14, 3.175221e-14, 3.162936e-14, 
    2.981157e-14, 2.505561e-14, 3.356756e-14, 1.201818e-14, 2.366352e-14, 
    5.160265e-14, 4.469417e-14, 4.376103e-14, 4.632475e-14, 3.072799e-14, 
    3.590202e-14, 2.311533e-14, 2.621665e-14, 2.12654e-14, 2.36421e-14, 
    2.400555e-14, 2.733314e-14, 2.95478e-14, 3.565311e-14, 4.11841e-14, 
    4.594711e-14, 4.48092e-14, 3.968184e-14, 3.139936e-14, 2.468212e-14, 
    2.606464e-14, 2.161842e-14, 3.46064e-14, 2.867842e-14, 3.088395e-14, 
    2.535161e-14, 3.84288e-14, 2.707184e-14, 4.175643e-14, 4.030124e-14, 
    3.601007e-14, 2.830173e-14, 2.675699e-14, 2.516781e-14, 2.614113e-14, 
    3.120541e-14, 3.209146e-14, 3.611085e-14, 3.7275e-14, 4.061526e-14, 
    4.352328e-14, 4.086096e-14, 3.818165e-14, 3.120346e-14, 2.567452e-14, 
    2.041647e-14, 1.92463e-14, 1.425253e-14, 1.824323e-14, 1.196702e-14, 
    1.719611e-14, 8.895534e-15, 2.649208e-14, 1.736895e-14, 3.582251e-14, 
    3.341156e-14, 2.932254e-14, 2.120315e-14, 2.5376e-14, 2.054353e-14, 
    3.212656e-14, 3.95117e-14, 4.158798e-14, 4.564759e-14, 4.149804e-14, 
    4.182597e-14, 3.807382e-14, 3.925462e-14, 3.098729e-14, 3.527021e-14, 
    2.401455e-14, 2.057929e-14, 1.263177e-14, 8.908236e-15, 5.947607e-15, 
    4.877096e-15, 4.578276e-15, 4.456976e-15,
  2.880588e-19, 2.462415e-19, 2.540362e-19, 2.227254e-19, 2.397624e-19, 
    2.197393e-19, 2.792325e-19, 2.446678e-19, 2.663872e-19, 2.84119e-19, 
    1.693738e-19, 2.213913e-19, 1.245086e-19, 1.510022e-19, 9.045997e-20, 
    1.28415e-19, 8.381287e-20, 9.14399e-20, 6.974475e-20, 7.557968e-20, 
    5.17657e-20, 6.715174e-20, 4.156028e-20, 5.521134e-20, 5.291745e-20, 
    6.770291e-20, 2.101925e-19, 1.75361e-19, 2.123855e-19, 2.071306e-19, 
    2.094787e-19, 2.394007e-19, 2.554812e-19, 2.914372e-19, 2.846777e-19, 
    2.583841e-19, 2.047956e-19, 2.220802e-19, 1.802442e-19, 1.81127e-19, 
    1.408553e-19, 1.582036e-19, 9.98954e-20, 1.147361e-19, 7.533018e-20, 
    8.425557e-20, 7.57349e-20, 7.825775e-20, 7.570238e-20, 8.905366e-20, 
    8.316363e-20, 9.554236e-20, 1.548545e-19, 1.354983e-19, 1.983305e-19, 
    2.438892e-19, 2.776523e-19, 3.033834e-19, 2.996541e-19, 2.926281e-19, 
    2.582351e-19, 2.284289e-19, 2.072931e-19, 1.938928e-19, 1.812541e-19, 
    1.462774e-19, 1.296881e-19, 9.705191e-20, 1.024992e-19, 9.338379e-20, 
    8.517868e-20, 7.246368e-20, 7.446712e-20, 6.918241e-20, 9.361877e-20, 
    7.685548e-20, 1.056873e-19, 9.721501e-20, 1.779019e-19, 2.173275e-19, 
    2.356604e-19, 2.52525e-19, 2.968071e-19, 2.657249e-19, 2.777075e-19, 
    2.497681e-19, 2.330105e-19, 2.412038e-19, 1.935346e-19, 2.112553e-19, 
    1.287449e-19, 1.610662e-19, 8.611095e-20, 1.013658e-19, 8.268825e-20, 
    9.19157e-20, 7.648075e-20, 9.029005e-20, 6.727898e-20, 6.282756e-20, 
    6.584838e-20, 5.473156e-20, 9.109854e-20, 7.573429e-20, 2.414355e-19, 
    2.400856e-19, 2.338634e-19, 2.62022e-19, 2.63814e-19, 2.916232e-19, 
    2.667904e-19, 2.566519e-19, 2.320635e-19, 2.182713e-19, 2.056683e-19, 
    1.796474e-19, 1.532261e-19, 1.206993e-19, 1.003283e-19, 8.799511e-20, 
    9.543535e-20, 8.884667e-20, 9.623167e-20, 9.98241e-20, 6.447238e-20, 
    8.310949e-20, 5.625056e-20, 5.756582e-20, 6.905951e-20, 5.741666e-20, 
    2.391409e-19, 2.469564e-19, 2.753843e-19, 2.529645e-19, 2.947634e-19, 
    2.70847e-19, 2.576915e-19, 2.108718e-19, 2.013974e-19, 1.928601e-19, 
    1.767005e-19, 1.572838e-19, 1.266593e-19, 1.033883e-19, 8.471639e-20, 
    8.60046e-20, 8.554961e-20, 8.167349e-20, 9.14855e-20, 8.013014e-20, 
    7.831703e-20, 8.311272e-20, 5.774341e-20, 6.43968e-20, 5.759399e-20, 
    6.186676e-20, 2.443982e-19, 2.314319e-19, 2.383807e-19, 2.25424e-19, 
    2.345016e-19, 1.95899e-19, 1.851937e-19, 1.401371e-19, 1.576514e-19, 
    1.303983e-19, 1.547304e-19, 1.502215e-19, 1.295609e-19, 1.53347e-19, 
    1.045915e-19, 1.363252e-19, 8.152516e-20, 1.087438e-19, 7.998342e-20, 
    8.479207e-20, 7.692778e-20, 7.029279e-20, 6.248017e-20, 4.956078e-20, 
    5.238456e-20, 4.264938e-20, 2.129519e-19, 1.976784e-19, 1.989958e-19, 
    1.837301e-19, 1.729439e-19, 1.509965e-19, 1.196964e-19, 1.309197e-19, 
    1.108093e-19, 1.070287e-19, 1.377845e-19, 1.183082e-19, 1.878681e-19, 
    1.752021e-19, 1.826758e-19, 2.117187e-19, 1.282735e-19, 1.677262e-19, 
    1.000114e-19, 1.175752e-19, 7.121541e-20, 9.242094e-20, 5.398142e-20, 
    4.132196e-20, 3.132732e-20, 2.177435e-20, 1.896549e-19, 1.996802e-19, 
    1.819677e-19, 1.591883e-19, 1.397874e-19, 1.164511e-19, 1.142177e-19, 
    1.101978e-19, 1.00212e-19, 9.227958e-20, 1.089444e-19, 9.035643e-20, 
    1.723419e-19, 1.251662e-19, 2.035562e-19, 1.773366e-19, 1.604776e-19, 
    1.67741e-19, 1.322443e-19, 1.24656e-19, 9.67113e-20, 1.105897e-19, 
    4.427296e-20, 6.893813e-20, 1.591863e-20, 2.60852e-20, 2.03262e-19, 
    1.8969e-19, 1.470681e-19, 1.66473e-19, 1.14991e-19, 1.041456e-19, 
    9.583127e-20, 8.583616e-20, 8.479986e-20, 7.924967e-20, 8.847086e-20, 
    7.960218e-20, 1.164043e-19, 9.885323e-20, 1.515906e-19, 1.374068e-19, 
    1.438209e-19, 1.510738e-19, 1.294208e-19, 1.086678e-19, 1.082522e-19, 
    1.020992e-19, 8.597356e-20, 1.14807e-19, 4.154536e-20, 8.12454e-20, 
    1.755776e-19, 1.523439e-19, 1.492017e-19, 1.578323e-19, 1.052019e-19, 
    1.226954e-19, 7.938239e-20, 8.991404e-20, 7.309066e-20, 8.117259e-20, 
    8.240744e-20, 9.370092e-20, 1.012059e-19, 1.218546e-19, 1.405189e-19, 
    1.565614e-19, 1.527312e-19, 1.354534e-19, 1.07474e-19, 8.470539e-20, 
    8.939831e-20, 7.429188e-20, 1.183179e-19, 9.826082e-20, 1.057297e-19, 
    8.697842e-20, 1.312261e-19, 9.281487e-20, 1.42448e-19, 1.375423e-19, 
    1.230603e-19, 9.698434e-20, 9.174707e-20, 8.635449e-20, 8.965782e-20, 
    1.068177e-19, 1.098155e-19, 1.234008e-19, 1.273318e-19, 1.386012e-19, 
    1.484009e-19, 1.394295e-19, 1.303921e-19, 1.068111e-19, 8.807442e-20, 
    7.020079e-20, 6.621454e-20, 4.916142e-20, 6.27948e-20, 4.136969e-20, 
    5.922202e-20, 3.080326e-20, 9.084847e-20, 5.981192e-20, 1.224268e-19, 
    1.142796e-19, 1.004429e-19, 7.287881e-20, 8.70612e-20, 7.063344e-20, 
    1.099342e-19, 1.348796e-19, 1.418803e-19, 1.555534e-19, 1.415771e-19, 
    1.426824e-19, 1.300282e-19, 1.340124e-19, 1.060795e-19, 1.20561e-19, 
    8.243803e-20, 7.075518e-20, 4.360997e-20, 3.084704e-20, 2.061603e-20, 
    1.690187e-20, 1.586333e-20, 1.544152e-20,
  2.114394e-25, 1.808954e-25, 1.865904e-25, 1.637086e-25, 1.761609e-25, 
    1.615256e-25, 2.049942e-25, 1.797455e-25, 1.956128e-25, 2.085625e-25, 
    1.246823e-25, 1.627333e-25, 9.18155e-26, 1.112302e-25, 6.682711e-26, 
    9.46794e-26, 6.194308e-26, 6.754694e-26, 5.159874e-26, 5.589054e-26, 
    3.83599e-26, 4.969081e-26, 3.084301e-26, 4.089903e-26, 3.920875e-26, 
    5.00964e-26, 1.545454e-25, 1.290646e-25, 1.56149e-25, 1.523064e-25, 
    1.540235e-25, 1.758966e-25, 1.876461e-25, 2.139061e-25, 2.089706e-25, 
    1.897668e-25, 1.505988e-25, 1.632369e-25, 1.326383e-25, 1.332843e-25, 
    1.037968e-25, 1.165042e-25, 7.375645e-26, 8.46482e-26, 5.570706e-26, 
    6.226842e-26, 5.600468e-26, 5.78597e-26, 5.598077e-26, 6.579398e-26, 
    6.146592e-26, 7.056006e-26, 1.140516e-25, 9.987123e-26, 1.458704e-25, 
    1.791765e-25, 2.038403e-25, 2.226275e-25, 2.199051e-25, 2.147755e-25, 
    1.896579e-25, 1.678777e-25, 1.524252e-25, 1.426243e-25, 1.333773e-25, 
    1.077692e-25, 9.561265e-26, 7.16686e-26, 7.566805e-26, 6.897476e-26, 
    6.294679e-26, 5.359886e-26, 5.507237e-26, 5.118501e-26, 6.914735e-26, 
    5.682867e-26, 7.800814e-26, 7.178837e-26, 1.309242e-25, 1.597623e-25, 
    1.731632e-25, 1.854863e-25, 2.178267e-25, 1.951291e-25, 2.038806e-25, 
    1.834722e-25, 1.712265e-25, 1.772143e-25, 1.423622e-25, 1.553226e-25, 
    9.492126e-26, 1.186003e-25, 6.363186e-26, 7.483597e-26, 6.111654e-26, 
    6.789644e-26, 5.655314e-26, 6.670228e-26, 4.978444e-26, 4.65081e-26, 
    4.873164e-26, 4.054554e-26, 6.729619e-26, 5.600423e-26, 1.773835e-25, 
    1.763971e-25, 1.718498e-25, 1.924242e-25, 1.937332e-25, 2.140419e-25, 
    1.959073e-25, 1.885013e-25, 1.705343e-25, 1.604524e-25, 1.51237e-25, 
    1.322016e-25, 1.12859e-25, 8.902228e-26, 7.407429e-26, 6.501626e-26, 
    7.048149e-26, 6.564191e-26, 7.106628e-26, 7.370411e-26, 4.771888e-26, 
    6.142614e-26, 4.166464e-26, 4.26335e-26, 5.109458e-26, 4.252363e-26, 
    1.757067e-25, 1.814177e-25, 2.02184e-25, 1.858075e-25, 2.163346e-25, 
    1.988702e-25, 1.892608e-25, 1.550422e-25, 1.481135e-25, 1.418689e-25, 
    1.30045e-25, 1.158306e-25, 9.339229e-26, 7.632071e-26, 6.260707e-26, 
    6.355371e-26, 6.321937e-26, 6.037069e-26, 6.758044e-26, 5.923621e-26, 
    5.790328e-26, 6.142851e-26, 4.276431e-26, 4.766325e-26, 4.265425e-26, 
    4.580074e-26, 1.795485e-25, 1.700727e-25, 1.751512e-25, 1.656813e-25, 
    1.723163e-25, 1.440918e-25, 1.3626e-25, 1.032706e-25, 1.160998e-25, 
    9.613322e-26, 1.139607e-25, 1.106584e-25, 9.551941e-26, 1.129476e-25, 
    7.720391e-26, 1.004773e-25, 6.026165e-26, 8.025136e-26, 5.912835e-26, 
    6.266269e-26, 5.688183e-26, 5.200193e-26, 4.625235e-26, 3.673451e-26, 
    3.881602e-26, 3.163655e-26, 1.565632e-25, 1.453934e-25, 1.46357e-25, 
    1.351891e-25, 1.272955e-25, 1.11226e-25, 8.828677e-26, 9.651542e-26, 
    8.176712e-26, 7.899269e-26, 1.015467e-25, 8.72687e-26, 1.382168e-25, 
    1.289483e-25, 1.344177e-25, 1.556614e-25, 9.457564e-26, 1.234762e-25, 
    7.384165e-26, 8.673103e-26, 5.268066e-26, 6.826755e-26, 3.99928e-26, 
    3.066705e-26, 2.328101e-26, 1.620576e-26, 1.395241e-25, 1.468576e-25, 
    1.338995e-25, 1.172252e-25, 1.030143e-25, 8.590639e-26, 8.426792e-26, 
    8.131839e-26, 7.398888e-26, 6.816373e-26, 8.039861e-26, 6.675104e-26, 
    1.268549e-25, 9.229765e-26, 1.496924e-25, 1.305105e-25, 1.181693e-25, 
    1.23487e-25, 9.748635e-26, 9.192355e-26, 7.141849e-26, 8.160595e-26, 
    3.283458e-26, 5.100528e-26, 1.185808e-26, 1.940089e-26, 1.494772e-25, 
    1.395497e-25, 1.083485e-25, 1.225588e-25, 8.483527e-26, 7.687655e-26, 
    7.077223e-26, 6.342993e-26, 6.266842e-26, 5.858894e-26, 6.536581e-26, 
    5.884809e-26, 8.587209e-26, 7.299127e-26, 1.116612e-25, 1.012699e-25, 
    1.059696e-25, 1.112826e-25, 9.541672e-26, 8.019563e-26, 7.989062e-26, 
    7.537437e-26, 6.35309e-26, 8.470025e-26, 3.0832e-26, 6.005602e-26, 
    1.292232e-25, 1.122129e-25, 1.099113e-25, 1.162322e-25, 7.765187e-26, 
    9.048598e-26, 5.868652e-26, 6.642606e-26, 5.406003e-26, 6.00025e-26, 
    6.091014e-26, 6.920769e-26, 7.471857e-26, 8.986943e-26, 1.035503e-25, 
    1.153016e-25, 1.124965e-25, 9.983837e-26, 7.931948e-26, 6.2599e-26, 
    6.604718e-26, 5.494349e-26, 8.727577e-26, 7.255629e-26, 7.803931e-26, 
    6.426927e-26, 9.674007e-26, 6.855689e-26, 1.049637e-25, 1.013692e-25, 
    9.075359e-26, 7.161898e-26, 6.777258e-26, 6.381081e-26, 6.623783e-26, 
    7.883781e-26, 8.103784e-26, 9.10032e-26, 9.388533e-26, 1.021451e-25, 
    1.093248e-25, 1.027521e-25, 9.612872e-26, 7.883297e-26, 6.507454e-26, 
    5.193425e-26, 4.900112e-26, 3.644006e-26, 4.648398e-26, 3.07023e-26, 
    4.38533e-26, 2.289332e-26, 6.71125e-26, 4.428773e-26, 9.028904e-26, 
    8.431334e-26, 7.415844e-26, 5.390421e-26, 6.433008e-26, 5.225253e-26, 
    8.112496e-26, 9.94178e-26, 1.045478e-25, 1.145634e-25, 1.043257e-25, 
    1.051355e-25, 9.586197e-26, 9.878223e-26, 7.829603e-26, 8.892081e-26, 
    6.093263e-26, 5.234209e-26, 3.234541e-26, 2.292572e-26, 1.53465e-26, 
    1.258881e-26, 1.181697e-26, 1.150337e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.01117137, 0.01118577, 0.01118297, 0.01119457, 0.01118813, 0.01119573, 
    0.01117428, 0.01118634, 0.01117864, 0.01117266, 0.01121704, 0.01119508, 
    0.01123968, 0.01122576, 0.01126068, 0.01123753, 0.01126534, 0.01126, 
    0.01127602, 0.01127143, 0.01129191, 0.01127813, 0.01130246, 0.01128861, 
    0.01129079, 0.01127768, 0.01119949, 0.01121431, 0.01119862, 0.01120073, 
    0.01119978, 0.01118827, 0.01118247, 0.01117025, 0.01117247, 0.01118143, 
    0.01120168, 0.01119481, 0.01121209, 0.0112117, 0.01123089, 0.01122224, 
    0.0112544, 0.01124526, 0.01127162, 0.01126501, 0.01127131, 0.0112694, 
    0.01127134, 0.01126163, 0.0112658, 0.01125724, 0.01122386, 0.01123369, 
    0.01120434, 0.01118664, 0.01117481, 0.01116642, 0.01116761, 0.01116987, 
    0.01118149, 0.01119237, 0.01120065, 0.01120619, 0.01121164, 0.01122815, 
    0.01123682, 0.01125626, 0.01125274, 0.01125869, 0.01126435, 0.01127386, 
    0.01127229, 0.01127648, 0.01125852, 0.01127047, 0.01125074, 0.01125614, 
    0.01121318, 0.01119666, 0.01118967, 0.01118351, 0.01116852, 0.01117888, 
    0.0111748, 0.01118448, 0.01119064, 0.01118759, 0.01120634, 0.01119906, 
    0.01123734, 0.01122088, 0.01126369, 0.01125346, 0.01126614, 0.01125967, 
    0.01127075, 0.01126078, 0.01127803, 0.01128179, 0.01127922, 0.01128905, 
    0.01126023, 0.01127132, 0.01118751, 0.01118801, 0.01119032, 0.01118016, 
    0.01117954, 0.0111702, 0.0111785, 0.01118204, 0.01119099, 0.01119629, 
    0.01120132, 0.01121236, 0.01122467, 0.01124182, 0.01125413, 0.01126236, 
    0.01125731, 0.01126177, 0.01125679, 0.01125444, 0.01128038, 0.01126584, 
    0.01128764, 0.01128643, 0.01127658, 0.01128657, 0.01118836, 0.0111855, 
    0.01117558, 0.01118334, 0.01116918, 0.01117712, 0.01118168, 0.01119923, 
    0.01120306, 0.01120663, 0.01121367, 0.01122268, 0.01123848, 0.01125219, 
    0.01126468, 0.01126376, 0.01126408, 0.01126688, 0.01125996, 0.01126801, 
    0.01126936, 0.01126583, 0.01128627, 0.01128044, 0.01128641, 0.01128261, 
    0.01118642, 0.01119123, 0.01118864, 0.01119352, 0.01119008, 0.01120536, 
    0.01120994, 0.01123127, 0.01122251, 0.01123643, 0.01122392, 0.01122614, 
    0.01123691, 0.01122459, 0.01125144, 0.01123327, 0.01126698, 0.01124889, 
    0.01126812, 0.01126462, 0.0112704, 0.01127558, 0.01128208, 0.01129406, 
    0.01129129, 0.01130129, 0.01119839, 0.01120461, 0.01120405, 0.01121056, 
    0.01121536, 0.01122575, 0.01124239, 0.01123613, 0.0112476, 0.01124991, 
    0.01123248, 0.01124319, 0.01120877, 0.01121436, 0.01121102, 0.01119888, 
    0.01123759, 0.01121777, 0.01125433, 0.01124361, 0.01127484, 0.01125934, 
    0.01128976, 0.01130274, 0.01131488, 0.01132909, 0.011208, 0.01120377, 
    0.01121133, 0.01122178, 0.01123144, 0.01124426, 0.01124557, 0.01124798, 
    0.0112542, 0.01125942, 0.01124875, 0.01126073, 0.01121567, 0.0112393, 
    0.01120218, 0.0112134, 0.01122116, 0.01121775, 0.01123542, 0.01123958, 
    0.01125648, 0.01124774, 0.01129955, 0.01127669, 0.01133984, 0.01132228, 
    0.0112023, 0.01120798, 0.01122772, 0.01121834, 0.01124511, 0.0112517, 
    0.01125705, 0.01126389, 0.01126462, 0.01126866, 0.01126203, 0.0112684, 
    0.01124429, 0.01125508, 0.01122546, 0.01123268, 0.01122935, 0.01122571, 
    0.01123695, 0.01124892, 0.01124916, 0.011253, 0.01126384, 0.01124522, 
    0.01130253, 0.01126724, 0.01121417, 0.01122511, 0.01122665, 0.01122242, 
    0.01125105, 0.01124068, 0.01126856, 0.01126104, 0.01127336, 0.01126724, 
    0.01126634, 0.01125847, 0.01125356, 0.01124116, 0.01123106, 0.01122303, 
    0.01122489, 0.01123371, 0.01124965, 0.01126469, 0.0112614, 0.01127242, 
    0.01124318, 0.01125547, 0.01125072, 0.01126308, 0.01123597, 0.01125911, 
    0.01123006, 0.0112326, 0.01124048, 0.01125631, 0.01125978, 0.01126352, 
    0.01126121, 0.01125005, 0.01124821, 0.01124028, 0.0112381, 0.01123205, 
    0.01122704, 0.01123162, 0.01123643, 0.01125005, 0.01126232, 0.01127566, 
    0.01127891, 0.01129449, 0.01128183, 0.01130273, 0.01128501, 0.01131563, 
    0.01126043, 0.01128445, 0.01124083, 0.01124553, 0.01125406, 0.01127355, 
    0.01126302, 0.01127532, 0.01124814, 0.01123403, 0.01123035, 0.01122352, 
    0.01123051, 0.01122994, 0.01123662, 0.01123447, 0.0112505, 0.01124189, 
    0.01126632, 0.01127522, 0.01130025, 0.01131554, 0.01133103, 0.01133787, 
    0.01133995, 0.01134081,
  3.668333e-05, 3.677487e-05, 3.675705e-05, 3.68309e-05, 3.678989e-05, 
    3.683827e-05, 3.670184e-05, 3.677856e-05, 3.672956e-05, 3.669149e-05, 
    3.697417e-05, 3.683418e-05, 3.711874e-05, 3.702975e-05, 3.725308e-05, 
    3.710498e-05, 3.728289e-05, 3.724867e-05, 3.735128e-05, 3.73219e-05, 
    3.745326e-05, 3.736484e-05, 3.752103e-05, 3.743208e-05, 3.744606e-05, 
    3.736195e-05, 3.686224e-05, 3.69568e-05, 3.685667e-05, 3.687015e-05, 
    3.686407e-05, 3.679079e-05, 3.675392e-05, 3.667624e-05, 3.669032e-05, 
    3.674733e-05, 3.687621e-05, 3.683239e-05, 3.69425e-05, 3.694001e-05, 
    3.70625e-05, 3.70073e-05, 3.721288e-05, 3.715441e-05, 3.732312e-05, 
    3.728075e-05, 3.732116e-05, 3.730889e-05, 3.732132e-05, 3.725916e-05, 
    3.72858e-05, 3.723104e-05, 3.701767e-05, 3.708044e-05, 3.689314e-05, 
    3.678049e-05, 3.670523e-05, 3.665189e-05, 3.665943e-05, 3.667383e-05, 
    3.674766e-05, 3.681689e-05, 3.686964e-05, 3.690493e-05, 3.693966e-05, 
    3.704504e-05, 3.710047e-05, 3.722477e-05, 3.720222e-05, 3.724032e-05, 
    3.727653e-05, 3.733744e-05, 3.73274e-05, 3.735425e-05, 3.723923e-05, 
    3.731574e-05, 3.71894e-05, 3.722399e-05, 3.694956e-05, 3.684419e-05, 
    3.679976e-05, 3.67605e-05, 3.666524e-05, 3.673106e-05, 3.670513e-05, 
    3.676671e-05, 3.680587e-05, 3.678648e-05, 3.690589e-05, 3.685951e-05, 
    3.710376e-05, 3.699864e-05, 3.727231e-05, 3.720684e-05, 3.728797e-05, 
    3.724656e-05, 3.731754e-05, 3.725366e-05, 3.73642e-05, 3.73883e-05, 
    3.737184e-05, 3.743488e-05, 3.725013e-05, 3.73212e-05, 3.678596e-05, 
    3.678913e-05, 3.680382e-05, 3.673923e-05, 3.673525e-05, 3.667587e-05, 
    3.672867e-05, 3.675118e-05, 3.680811e-05, 3.684184e-05, 3.687387e-05, 
    3.694423e-05, 3.70228e-05, 3.713242e-05, 3.721109e-05, 3.726382e-05, 
    3.723146e-05, 3.726003e-05, 3.722811e-05, 3.721312e-05, 3.73793e-05, 
    3.728608e-05, 3.742582e-05, 3.741808e-05, 3.73549e-05, 3.741895e-05, 
    3.679135e-05, 3.677314e-05, 3.671007e-05, 3.675943e-05, 3.66694e-05, 
    3.671987e-05, 3.67489e-05, 3.686058e-05, 3.688498e-05, 3.690775e-05, 
    3.695258e-05, 3.701013e-05, 3.711101e-05, 3.719869e-05, 3.727862e-05, 
    3.727276e-05, 3.727482e-05, 3.729272e-05, 3.724845e-05, 3.729997e-05, 
    3.730866e-05, 3.728602e-05, 3.741704e-05, 3.737963e-05, 3.741791e-05, 
    3.739354e-05, 3.677905e-05, 3.680965e-05, 3.679312e-05, 3.682422e-05, 
    3.680235e-05, 3.689968e-05, 3.692884e-05, 3.706498e-05, 3.700902e-05, 
    3.709794e-05, 3.701802e-05, 3.703221e-05, 3.710104e-05, 3.702231e-05, 
    3.719394e-05, 3.707777e-05, 3.729341e-05, 3.717764e-05, 3.730067e-05, 
    3.727827e-05, 3.73153e-05, 3.73485e-05, 3.739015e-05, 3.746708e-05, 
    3.744925e-05, 3.751346e-05, 3.68552e-05, 3.689488e-05, 3.68913e-05, 
    3.693275e-05, 3.696341e-05, 3.702971e-05, 3.713603e-05, 3.709604e-05, 
    3.716937e-05, 3.718413e-05, 3.707265e-05, 3.714117e-05, 3.692136e-05, 
    3.695701e-05, 3.693573e-05, 3.685838e-05, 3.710538e-05, 3.697877e-05, 
    3.721241e-05, 3.714383e-05, 3.734378e-05, 3.72445e-05, 3.743946e-05, 
    3.752285e-05, 3.760082e-05, 3.769229e-05, 3.691644e-05, 3.688949e-05, 
    3.693765e-05, 3.70044e-05, 3.706602e-05, 3.714802e-05, 3.715636e-05, 
    3.717177e-05, 3.721153e-05, 3.724499e-05, 3.717672e-05, 3.725337e-05, 
    3.696545e-05, 3.711632e-05, 3.687938e-05, 3.695093e-05, 3.700043e-05, 
    3.697863e-05, 3.709144e-05, 3.711804e-05, 3.722617e-05, 3.717022e-05, 
    3.750236e-05, 3.735563e-05, 3.776155e-05, 3.764845e-05, 3.68801e-05, 
    3.69163e-05, 3.70423e-05, 3.698237e-05, 3.715345e-05, 3.71956e-05, 
    3.722978e-05, 3.727359e-05, 3.727825e-05, 3.730418e-05, 3.72617e-05, 
    3.730247e-05, 3.714819e-05, 3.721716e-05, 3.702781e-05, 3.707397e-05, 
    3.705271e-05, 3.702944e-05, 3.710123e-05, 3.717782e-05, 3.717931e-05, 
    3.72039e-05, 3.72734e-05, 3.715414e-05, 3.752153e-05, 3.729513e-05, 
    3.695577e-05, 3.702562e-05, 3.703542e-05, 3.700841e-05, 3.719138e-05, 
    3.712512e-05, 3.730353e-05, 3.725531e-05, 3.733426e-05, 3.729505e-05, 
    3.728929e-05, 3.723886e-05, 3.720749e-05, 3.712818e-05, 3.706361e-05, 
    3.701231e-05, 3.702423e-05, 3.708058e-05, 3.718247e-05, 3.727874e-05, 
    3.725768e-05, 3.732826e-05, 3.714106e-05, 3.721968e-05, 3.718934e-05, 
    3.726839e-05, 3.7095e-05, 3.72431e-05, 3.705719e-05, 3.707347e-05, 
    3.71238e-05, 3.722511e-05, 3.72473e-05, 3.727124e-05, 3.725644e-05, 
    3.718503e-05, 3.717326e-05, 3.712254e-05, 3.710861e-05, 3.706991e-05, 
    3.703793e-05, 3.706719e-05, 3.709793e-05, 3.7185e-05, 3.726353e-05, 
    3.7349e-05, 3.736983e-05, 3.746987e-05, 3.738864e-05, 3.752282e-05, 
    3.740906e-05, 3.76057e-05, 3.725146e-05, 3.740543e-05, 3.712604e-05, 
    3.715612e-05, 3.721072e-05, 3.73355e-05, 3.726802e-05, 3.734686e-05, 
    3.717279e-05, 3.708259e-05, 3.705906e-05, 3.701545e-05, 3.706006e-05, 
    3.705643e-05, 3.709911e-05, 3.708538e-05, 3.718789e-05, 3.713282e-05, 
    3.728918e-05, 3.73462e-05, 3.750678e-05, 3.76051e-05, 3.770479e-05, 
    3.774883e-05, 3.776221e-05, 3.776782e-05,
  8.811749e-10, 8.839173e-10, 8.833831e-10, 8.85597e-10, 8.843674e-10, 
    8.858181e-10, 8.81729e-10, 8.840278e-10, 8.825593e-10, 8.814192e-10, 
    8.898973e-10, 8.856952e-10, 8.943256e-10, 8.915667e-10, 8.985015e-10, 
    8.93898e-10, 8.994289e-10, 8.983642e-10, 9.015575e-10, 9.006425e-10, 
    9.047348e-10, 9.019797e-10, 9.068481e-10, 9.040745e-10, 9.045102e-10, 
    9.018895e-10, 8.86537e-10, 8.893756e-10, 8.863698e-10, 8.867744e-10, 
    8.865919e-10, 8.843943e-10, 8.832895e-10, 8.809624e-10, 8.813841e-10, 
    8.830917e-10, 8.869562e-10, 8.856417e-10, 8.889459e-10, 8.888711e-10, 
    8.925783e-10, 8.908921e-10, 8.972513e-10, 8.954342e-10, 9.006806e-10, 
    8.993621e-10, 9.006195e-10, 9.002377e-10, 9.006245e-10, 8.986903e-10, 
    8.995193e-10, 8.978159e-10, 8.912037e-10, 8.931357e-10, 8.874642e-10, 
    8.840856e-10, 8.818306e-10, 8.802333e-10, 8.804592e-10, 8.808905e-10, 
    8.831018e-10, 8.851768e-10, 8.86759e-10, 8.878179e-10, 8.888604e-10, 
    8.920365e-10, 8.93758e-10, 8.976209e-10, 8.969198e-10, 8.981045e-10, 
    8.992307e-10, 9.011265e-10, 9.008139e-10, 9.016499e-10, 8.980705e-10, 
    9.004509e-10, 8.965214e-10, 8.975968e-10, 8.891584e-10, 8.859957e-10, 
    8.846635e-10, 8.834864e-10, 8.806331e-10, 8.826044e-10, 8.818277e-10, 
    8.836724e-10, 8.848465e-10, 8.842652e-10, 8.878468e-10, 8.864551e-10, 
    8.9386e-10, 8.906321e-10, 8.990995e-10, 8.970634e-10, 8.995868e-10, 
    8.982985e-10, 9.00507e-10, 8.985194e-10, 9.019597e-10, 9.027104e-10, 
    9.021978e-10, 9.041618e-10, 8.984096e-10, 9.006209e-10, 8.842496e-10, 
    8.843445e-10, 8.847849e-10, 8.828492e-10, 8.8273e-10, 8.809515e-10, 
    8.825327e-10, 8.832072e-10, 8.849134e-10, 8.859252e-10, 8.86886e-10, 
    8.889978e-10, 8.913582e-10, 8.947507e-10, 8.971955e-10, 8.988352e-10, 
    8.978289e-10, 8.987174e-10, 8.977247e-10, 8.972587e-10, 9.024301e-10, 
    8.995279e-10, 9.038794e-10, 9.036381e-10, 9.016703e-10, 9.036653e-10, 
    8.844109e-10, 8.838653e-10, 8.819754e-10, 8.834544e-10, 8.807576e-10, 
    8.822691e-10, 8.831391e-10, 8.864873e-10, 8.872194e-10, 8.879026e-10, 
    8.892485e-10, 8.909772e-10, 8.940855e-10, 8.968101e-10, 8.992957e-10, 
    8.991133e-10, 8.991776e-10, 8.997343e-10, 8.983573e-10, 8.999603e-10, 
    9.002307e-10, 8.995258e-10, 9.036059e-10, 9.024403e-10, 9.03633e-10, 
    9.028737e-10, 8.840423e-10, 8.849597e-10, 8.844642e-10, 8.853966e-10, 
    8.847408e-10, 8.876606e-10, 8.885357e-10, 8.926556e-10, 8.909439e-10, 
    8.936794e-10, 8.912144e-10, 8.916409e-10, 8.937757e-10, 8.913432e-10, 
    8.966627e-10, 8.93053e-10, 8.99756e-10, 8.961561e-10, 8.999819e-10, 
    8.99285e-10, 9.004373e-10, 9.014708e-10, 9.027681e-10, 9.051655e-10, 
    9.046098e-10, 9.066119e-10, 8.863257e-10, 8.875166e-10, 8.87409e-10, 
    8.886532e-10, 8.895738e-10, 8.915655e-10, 8.948629e-10, 8.936201e-10, 
    8.958991e-10, 8.963578e-10, 8.928936e-10, 8.950228e-10, 8.883114e-10, 
    8.893817e-10, 8.887425e-10, 8.864212e-10, 8.939104e-10, 8.900352e-10, 
    8.972365e-10, 8.951052e-10, 9.013238e-10, 8.982344e-10, 9.043045e-10, 
    9.069052e-10, 9.093389e-10, 9.121969e-10, 8.881635e-10, 8.873546e-10, 
    8.888003e-10, 8.908052e-10, 8.926879e-10, 8.952357e-10, 8.954949e-10, 
    8.959734e-10, 8.972093e-10, 8.982497e-10, 8.961273e-10, 8.985102e-10, 
    8.896354e-10, 8.942503e-10, 8.870514e-10, 8.89199e-10, 8.906857e-10, 
    8.900308e-10, 8.934773e-10, 8.943038e-10, 8.976646e-10, 8.959253e-10, 
    9.062659e-10, 9.01693e-10, 9.143628e-10, 9.108266e-10, 8.870727e-10, 
    8.881594e-10, 8.919513e-10, 8.901432e-10, 8.954043e-10, 8.967143e-10, 
    8.977767e-10, 8.991393e-10, 8.992843e-10, 9.000911e-10, 8.987693e-10, 
    9.000378e-10, 8.95241e-10, 8.973844e-10, 8.915085e-10, 8.929346e-10, 
    8.922741e-10, 8.915576e-10, 8.937814e-10, 8.961615e-10, 8.962079e-10, 
    8.969722e-10, 8.991338e-10, 8.954257e-10, 9.068643e-10, 8.998097e-10, 
    8.893444e-10, 8.914429e-10, 8.917376e-10, 8.909254e-10, 8.965831e-10, 
    8.945236e-10, 9.000708e-10, 8.985707e-10, 9.010273e-10, 8.99807e-10, 
    8.996277e-10, 8.980592e-10, 8.970838e-10, 8.946189e-10, 8.926129e-10, 
    8.910426e-10, 8.914008e-10, 8.931398e-10, 8.963061e-10, 8.992995e-10, 
    8.986444e-10, 9.008405e-10, 8.950192e-10, 8.974627e-10, 8.965197e-10, 
    8.989776e-10, 8.93588e-10, 8.981911e-10, 8.924135e-10, 8.92919e-10, 
    8.944827e-10, 8.976315e-10, 8.983215e-10, 8.990663e-10, 8.986058e-10, 
    8.963857e-10, 8.960199e-10, 8.944436e-10, 8.940108e-10, 8.928085e-10, 
    8.918153e-10, 8.92724e-10, 8.93679e-10, 8.963848e-10, 8.988265e-10, 
    9.014862e-10, 9.021352e-10, 9.052527e-10, 9.027212e-10, 9.069044e-10, 
    9.033573e-10, 9.094915e-10, 8.984512e-10, 9.03244e-10, 8.945524e-10, 
    8.954874e-10, 8.971844e-10, 9.010661e-10, 8.98966e-10, 9.014198e-10, 
    8.960053e-10, 8.932024e-10, 8.924717e-10, 8.911372e-10, 8.925026e-10, 
    8.923898e-10, 8.937154e-10, 8.932892e-10, 8.964746e-10, 8.94763e-10, 
    8.996244e-10, 9.013993e-10, 9.064037e-10, 9.094726e-10, 9.125877e-10, 
    9.139648e-10, 9.143835e-10, 9.145588e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.6550256, 0.622774, 0.6290133, 0.603233, 0.6175004, 0.6006691, 0.648457, 
    0.6215008, 0.6386777, 0.6521081, 0.5540715, 0.6020899, 0.5055733, 
    0.5351748, 0.4617738, 0.5101389, 0.4523387, 0.4631328, 0.4309793, 
    0.4400891, 0.400084, 0.4268033, 0.3800653, 0.4063925, 0.4022162, 
    0.427698, 0.5923362, 0.5599834, 0.594269, 0.5896189, 0.5917048, 
    0.6172038, 0.6301585, 0.6575081, 0.6525232, 0.6324461, 0.5875314, 
    0.6026802, 0.564721, 0.5655702, 0.5241977, 0.5427238, 0.4745585, 
    0.4934337, 0.4397072, 0.4529785, 0.4403264, 0.4441469, 0.4402767, 
    0.4598083, 0.451396, 0.468743, 0.5392371, 0.5182294, 0.5816803, 
    0.6208696, 0.6472685, 0.6661547, 0.6634774, 0.6583796, 0.632329, 
    0.6080762, 0.5897633, 0.5776016, 0.5656923, 0.5301157, 0.5116103, 
    0.4707757, 0.477973, 0.4658076, 0.4543081, 0.435272, 0.4383813, 
    0.4300809, 0.4661286, 0.4420317, 0.4820914, 0.4709938, 0.5624587, 
    0.5985832, 0.6141205, 0.6278124, 0.6614203, 0.6381664, 0.6473101, 
    0.6256105, 0.6119174, 0.6186804, 0.5772702, 0.5932742, 0.5105208, 
    0.5456727, 0.4556432, 0.4764924, 0.4507034, 0.46379, 0.4414629, 
    0.4615365, 0.4270104, 0.4196484, 0.4246728, 0.4055262, 0.4626599, 
    0.4403257, 0.6188698, 0.6177653, 0.6126277, 0.6352925, 0.6366861, 
    0.6576444, 0.6389887, 0.6310825, 0.6111268, 0.5994009, 0.5883129, 
    0.5641459, 0.537527, 0.5010463, 0.4751294, 0.4583184, 0.4685982, 
    0.4595176, 0.469673, 0.4744641, 0.4223995, 0.4513173, 0.4082546, 
    0.4105863, 0.429884, 0.4103233, 0.6169903, 0.6233506, 0.6455553, 
    0.6281618, 0.6599362, 0.6421037, 0.6319017, 0.5929365, 0.5844686, 
    0.5766453, 0.5612889, 0.5417703, 0.5080957, 0.4791286, 0.4536431, 
    0.4554912, 0.4548401, 0.4492184, 0.4631958, 0.446941, 0.4442362, 
    0.4513218, 0.410899, 0.4222735, 0.4106359, 0.4180236, 0.6212815, 
    0.6105988, 0.6163652, 0.6055332, 0.6131584, 0.5794524, 0.5694536, 
    0.5234053, 0.5421519, 0.5124276, 0.5391069, 0.5343447, 0.5114642, 
    0.5376538, 0.4806842, 0.5191596, 0.4490005, 0.4859797, 0.4467233, 
    0.4537521, 0.4421409, 0.4318516, 0.4190623, 0.3959313, 0.4012322, 
    0.3822544, 0.5947661, 0.5810843, 0.5822868, 0.5680611, 0.5576086, 
    0.5351685, 0.4998415, 0.5130258, 0.4885726, 0.4838048, 0.5207915, 
    0.4981655, 0.5719807, 0.5598268, 0.5670548, 0.5936826, 0.5099744, 
    0.5524232, 0.4747117, 0.4972757, 0.433312, 0.4644867, 0.4041644, 
    0.3795677, 0.3571444, 0.3318709, 0.573658, 0.5829101, 0.5663769, 
    0.5437419, 0.5230178, 0.4959059, 0.4927972, 0.4878075, 0.4749759, 
    0.4642916, 0.4862322, 0.4616289, 0.5570162, 0.5063468, 0.5864177, 
    0.5619085, 0.5450687, 0.5524375, 0.514541, 0.5057461, 0.4703185, 
    0.4882979, 0.3855658, 0.4296898, 0.3133472, 0.3438731, 0.5861524, 
    0.5736907, 0.5309677, 0.5511639, 0.4937463, 0.4801083, 0.4691331, 
    0.4552507, 0.4537633, 0.4456316, 0.4589891, 0.4461566, 0.4958487, 
    0.4731786, 0.5357986, 0.5203699, 0.5274487, 0.5352505, 0.5113011, 
    0.4858833, 0.4853574, 0.4774517, 0.455449, 0.4935207, 0.3800358, 
    0.4485908, 0.5601932, 0.5365965, 0.5332566, 0.5423391, 0.4814689, 
    0.5034273, 0.4458294, 0.4610122, 0.4362498, 0.4484817, 0.4502935, 
    0.4662408, 0.4762828, 0.5024269, 0.5238266, 0.541019, 0.5370046, 
    0.5181788, 0.4843713, 0.4536276, 0.4602916, 0.438111, 0.4981768, 
    0.472391, 0.4821463, 0.4568787, 0.5133772, 0.4650294, 0.525948, 
    0.5205211, 0.5038605, 0.4706853, 0.4635573, 0.4559909, 0.4606543, 
    0.4835363, 0.4873279, 0.5042638, 0.5088797, 0.5217012, 0.5323993, 
    0.5226212, 0.5124203, 0.4835277, 0.4584306, 0.4317056, 0.4252734, 
    0.39517, 0.4195939, 0.3796689, 0.4134858, 0.3558739, 0.4623141, 
    0.4145064, 0.5031079, 0.4928733, 0.4752808, 0.4359206, 0.4569962, 
    0.4323924, 0.4874769, 0.5175321, 0.5253253, 0.5399678, 0.5249922, 
    0.5262048, 0.5120013, 0.5165508, 0.4825937, 0.5008799, 0.4503383, 
    0.4325851, 0.384221, 0.3559797, 0.3284368, 0.3166825, 0.3131561, 0.311689,
  0.9803688, 0.9605812, 0.9644024, 0.9486349, 0.9573536, 0.9470698, 
    0.9763314, 0.9598023, 0.9703278, 0.9785748, 0.9187353, 0.947937, 
    0.8894766, 0.9073034, 0.8283351, 0.89222, 0.8239949, 0.8289608, 
    0.8142258, 0.8183823, 0.8002425, 0.8123254, 0.7912779, 0.8030829, 
    0.8012015, 0.8127323, 0.9419871, 0.9223187, 0.9431654, 0.9403315, 
    0.9416022, 0.9571726, 0.9651051, 0.9818947, 0.9788299, 0.9665066, 
    0.9390599, 0.9482967, 0.9251902, 0.9257056, 0.9006809, 0.9118646, 
    0.8342393, 0.8430067, 0.8182077, 0.8242881, 0.8184909, 0.8202384, 
    0.8184682, 0.8274292, 0.8235616, 0.8315498, 0.9097571, 0.8970859, 
    0.9354973, 0.9594168, 0.9756016, 0.9872156, 0.9855675, 0.9824311, 
    0.9664348, 0.951592, 0.9404188, 0.9330156, 0.9257797, 0.9042513, 
    0.8931041, 0.8324897, 0.8358209, 0.8301949, 0.8248989, 0.8161827, 
    0.817602, 0.8138169, 0.8303426, 0.8192709, 0.837731, 0.83259, 0.9238204, 
    0.9457965, 0.9552878, 0.9636669, 0.9843017, 0.9700145, 0.9756273, 
    0.9623176, 0.9539395, 0.9580753, 0.9328141, 0.9425587, 0.892449, 
    0.9136485, 0.8255126, 0.8351348, 0.8232436, 0.8292636, 0.8190107, 
    0.8282249, 0.8124197, 0.809077, 0.8113573, 0.8026919, 0.8287427, 
    0.8184907, 0.9581913, 0.9575157, 0.9543735, 0.9682518, 0.9691064, 
    0.9819787, 0.9705186, 0.9656705, 0.953456, 0.9462954, 0.9395354, 
    0.9248414, 0.9087244, 0.8867589, 0.8345036, 0.826743, 0.8314827, 
    0.827295, 0.8319795, 0.8341953, 0.8103251, 0.8235256, 0.8039226, 
    0.8049753, 0.8137274, 0.8048565, 0.9570414, 0.9609336, 0.9745494, 
    0.9638804, 0.9833884, 0.9724304, 0.9661731, 0.9423535, 0.9371941, 
    0.9324344, 0.9231079, 0.9112881, 0.8909912, 0.8363569, 0.8245932, 
    0.8254426, 0.8251433, 0.8225623, 0.8289897, 0.8215182, 0.8202796, 
    0.8235274, 0.8051166, 0.8102676, 0.8049977, 0.8083401, 0.959667, 
    0.9531335, 0.9566591, 0.950039, 0.9546984, 0.9341424, 0.9280647, 
    0.900204, 0.9115189, 0.8935951, 0.9096783, 0.9068022, 0.8930171, 
    0.9088002, 0.8370789, 0.8976468, 0.8224624, 0.8395387, 0.8214185, 
    0.8246433, 0.8193204, 0.8146234, 0.8088109, 0.7983758, 0.8007582, 
    0.7922539, 0.9434683, 0.9351348, 0.935866, 0.927218, 0.9208764, 
    0.9072992, 0.8860359, 0.8939543, 0.8407431, 0.8385268, 0.8986281, 
    0.885031, 0.9295992, 0.9222221, 0.9266072, 0.942808, 0.8921204, 
    0.9177351, 0.8343102, 0.8844972, 0.8152889, 0.8295856, 0.8020785, 
    0.7910567, 0.7811152, 0.7700485, 0.9306183, 0.9362453, 0.9261952, 
    0.912481, 0.8999698, 0.8836762, 0.8427101, 0.8403873, 0.8344323, 
    0.829495, 0.8396553, 0.8282675, 0.9205194, 0.8899406, 0.9383813, 
    0.9234849, 0.9132832, 0.9177431, 0.8948655, 0.8895792, 0.8322782, 
    0.8406153, 0.7937337, 0.8136395, 0.7620388, 0.7752852, 0.9382194, 
    0.9306378, 0.9047641, 0.9169717, 0.8431524, 0.8368111, 0.8317299, 
    0.8253323, 0.8246486, 0.8209184, 0.8270517, 0.8211588, 0.883642, 
    0.8336005, 0.9076796, 0.8983746, 0.9026405, 0.9073486, 0.8929171, 
    0.8394932, 0.8392481, 0.8355796, 0.8254259, 0.8430473, 0.7912667, 
    0.8222767, 0.9224433, 0.9081627, 0.906145, 0.9116317, 0.8374423, 
    0.8881873, 0.8210089, 0.8279833, 0.8166288, 0.8222244, 0.8230554, 
    0.8303943, 0.8350377, 0.8875871, 0.9004572, 0.9108336, 0.9084079, 
    0.8970553, 0.8387905, 0.8245865, 0.827652, 0.8174785, 0.8850373, 
    0.8332365, 0.8377571, 0.8260807, 0.8941658, 0.8298376, 0.9017355, 
    0.8984653, 0.8884473, 0.8324482, 0.8291563, 0.8256727, 0.8278185, 
    0.8384025, 0.8401644, 0.8886892, 0.8914621, 0.8991761, 0.9056273, 
    0.8997306, 0.8935906, 0.8383982, 0.826795, 0.8145569, 0.81163, 0.7980353, 
    0.8090532, 0.7911032, 0.8062888, 0.780557, 0.8285846, 0.8067491, 
    0.8879954, 0.8427455, 0.8345743, 0.8164794, 0.8261348, 0.8148704, 
    0.8402336, 0.8966665, 0.9013602, 0.9101985, 0.9011594, 0.9018904, 
    0.893338, 0.8960748, 0.8379645, 0.8866584, 0.8230762, 0.814958, 
    0.7931321, 0.7806026, 0.7685559, 0.7634738, 0.7619565, 0.7613263,
  1.164514, 1.165756, 1.165537, 1.16637, 1.165932, 1.166442, 1.164789, 
    1.165799, 1.165178, 1.164638, 1.167393, 1.166402, 1.167558, 1.167566, 
    1.207629, 1.167583, 1.205616, 1.207917, 1.200938, 1.202954, 1.193841, 
    1.200002, 1.189007, 1.195325, 1.194345, 1.200203, 1.166663, 1.167312, 
    1.166614, 1.166731, 1.166679, 1.165942, 1.165496, 1.164408, 1.164621, 
    1.165412, 1.166781, 1.166386, 1.16724, 1.167226, 1.167605, 1.167513, 
    1.210309, 1.21417, 1.20287, 1.205754, 1.203006, 1.203842, 1.202995, 
    1.207212, 1.205413, 1.209097, 1.16754, 1.167606, 1.166915, 1.16582, 
    1.164838, 1.164025, 1.164145, 1.16437, 1.165417, 1.166228, 1.166727, 
    1.167002, 1.167224, 1.167589, 1.167589, 1.209522, 1.211016, 1.208481, 
    1.206039, 1.201892, 1.202579, 1.200737, 1.208548, 1.20338, 1.211863, 
    1.209567, 1.167275, 1.166499, 1.166041, 1.16558, 1.164237, 1.165197, 
    1.164836, 1.165658, 1.166111, 1.165894, 1.167009, 1.16664, 1.167585, 
    1.167486, 1.206325, 1.21071, 1.205264, 1.208055, 1.203255, 1.207579, 
    1.200049, 1.198383, 1.199522, 1.195122, 1.207817, 1.203006, 1.165887, 
    1.165924, 1.166088, 1.165307, 1.165254, 1.164402, 1.165166, 1.165462, 
    1.166135, 1.166477, 1.166762, 1.167249, 1.167552, 1.167525, 1.210427, 
    1.206896, 1.209066, 1.207151, 1.209291, 1.210289, 1.199008, 1.205396, 
    1.195759, 1.196301, 1.200693, 1.19624, 1.165949, 1.165736, 1.164907, 
    1.165568, 1.164302, 1.165045, 1.165432, 1.166648, 1.166853, 1.167021, 
    1.167293, 1.167521, 1.167573, 1.211254, 1.205896, 1.206292, 1.206153, 
    1.204943, 1.20793, 1.20445, 1.203862, 1.205397, 1.196373, 1.198979, 
    1.196312, 1.198012, 1.165807, 1.166151, 1.165969, 1.166303, 1.166072, 
    1.166963, 1.167158, 1.167606, 1.167518, 1.167592, 1.167541, 1.167571, 
    1.167588, 1.167551, 1.211574, 1.167606, 1.204896, 1.212658, 1.204403, 
    1.20592, 1.203404, 1.201132, 1.198249, 1.192855, 1.194113, 1.189546, 
    1.166601, 1.166928, 1.166902, 1.167183, 1.167347, 1.167567, 1.167515, 
    1.167595, 1.213186, 1.212214, 1.167607, 1.167499, 1.167112, 1.167315, 
    1.1672, 1.166629, 1.167583, 1.167413, 1.210341, 1.167491, 1.201457, 
    1.208202, 1.194803, 1.188884, 1.183208, 1.176438, 1.16708, 1.166888, 
    1.167212, 1.167504, 1.167606, 1.167477, 1.214041, 1.21303, 1.210395, 
    1.208161, 1.21271, 1.207599, 1.167354, 1.167563, 1.166807, 1.167284, 
    1.167492, 1.167414, 1.167599, 1.16756, 1.209426, 1.21313, 1.190355, 
    1.200649, 1.171184, 1.179706, 1.166814, 1.16708, 1.167587, 1.167429, 
    1.214233, 1.211456, 1.209178, 1.206241, 1.205922, 1.204165, 1.207038, 
    1.20428, 1.167476, 1.210022, 1.167563, 1.167607, 1.167598, 1.167566, 
    1.167588, 1.212638, 1.212531, 1.210908, 1.206283, 1.214187, 1.188999, 
    1.204807, 1.16731, 1.167558, 1.167577, 1.167516, 1.211735, 1.167544, 
    1.204208, 1.207468, 1.202108, 1.204784, 1.205175, 1.208572, 1.210666, 
    1.167536, 1.167605, 1.167527, 1.167556, 1.167606, 1.21233, 1.205893, 
    1.207315, 1.202519, 1.1675, 1.209858, 1.211874, 1.206589, 1.167596, 
    1.208317, 1.167602, 1.167607, 1.167547, 1.209503, 1.208006, 1.206399, 
    1.207392, 1.212159, 1.212933, 1.16755, 1.167577, 1.167607, 1.167581, 
    1.167606, 1.167592, 1.212157, 1.206919, 1.2011, 1.199658, 1.192673, 
    1.19837, 1.188909, 1.19697, 1.182877, 1.207744, 1.197206, 1.167542, 
    1.214057, 1.210459, 1.202035, 1.206614, 1.201252, 1.212963, 1.167605, 
    1.167603, 1.167535, 1.167604, 1.167601, 1.167591, 1.167603, 1.211966, 
    1.167524, 1.205185, 1.201295, 1.190027, 1.182905, 1.175484, 1.17215, 
    1.171129, 1.170701,
  0.5108865, 0.5006445, 0.5026337, 0.4943883, 0.4989603, 0.4935643, 
    0.5088083, 0.5002381, 0.5057072, 0.509964, 0.478443, 0.494021, 0.4623517, 
    0.4722223, 0.4475445, 0.4638847, 0.4442533, 0.4480168, 0.4367115, 
    0.4399444, 0.425548, 0.4352212, 0.4181284, 0.4278544, 0.4263292, 
    0.4355409, 0.490881, 0.4803779, 0.4915041, 0.4900041, 0.4906773, 
    0.4988654, 0.5029982, 0.5116711, 0.5100953, 0.5037264, 0.4893298, 
    0.4942108, 0.4819254, 0.4822023, 0.4685808, 0.4747145, 0.451968, 
    0.4584284, 0.4398094, 0.4444774, 0.4400282, 0.4413765, 0.4400107, 
    0.4468609, 0.4439233, 0.4499609, 0.4735645, 0.4665918, 0.487437, 
    0.5000364, 0.5084319, 0.5143995, 0.5135553, 0.5119463, 0.5036891, 
    0.4959429, 0.4900508, 0.4861151, 0.4822421, 0.4705464, 0.464378, 
    0.4506633, 0.4531427, 0.4489446, 0.4449424, 0.438238, 0.4393402, 
    0.4363913, 0.4490559, 0.4406305, 0.454556, 0.4507388, 0.4811865, 
    0.4928935, 0.4978789, 0.5022511, 0.5129063, 0.5055447, 0.508445, 
    0.5015494, 0.4971739, 0.4993375, 0.4860076, 0.4911835, 0.4640129, 
    0.4756854, 0.4454088, 0.4526337, 0.4436806, 0.448245, 0.4404297, 
    0.4474622, 0.4352951, 0.4326546, 0.4344586, 0.4275387, 0.4478526, 
    0.4400279, 0.4993979, 0.499045, 0.4974014, 0.5046316, 0.5050745, 
    0.5117141, 0.505806, 0.5032924, 0.4969207, 0.4931566, 0.4895824, 
    0.4817377, 0.4729998, 0.4608276, 0.4521646, 0.4463421, 0.4499109, 
    0.4467598, 0.4502825, 0.4519356, 0.4336433, 0.4438957, 0.4285325, 
    0.4293797, 0.4363211, 0.4292843, 0.4987972, 0.5008286, 0.5078891, 
    0.5023625, 0.5124379, 0.5067946, 0.5035531, 0.4910745, 0.4883397, 
    0.4858048, 0.480805, 0.4744002, 0.4631994, 0.4535396, 0.4447099, 
    0.4453558, 0.4451284, 0.4431598, 0.4480387, 0.4423599, 0.4414079, 
    0.4438973, 0.4294932, 0.4335983, 0.4293978, 0.4320696, 0.5001683, 
    0.4967515, 0.4985974, 0.495127, 0.4975713, 0.4867151, 0.4834672, 
    0.468317, 0.474526, 0.4646519, 0.4735216, 0.4719477, 0.4643289, 
    0.4730418, 0.4540733, 0.466902, 0.4430833, 0.4558863, 0.4422833, 
    0.444748, 0.4406691, 0.4370221, 0.4324437, 0.424022, 0.4259691, 
    0.4189478, 0.4916644, 0.487244, 0.4876336, 0.483014, 0.4796018, 
    0.4722203, 0.4604214, 0.4648523, 0.4567722, 0.4551427, 0.4674465, 
    0.4598556, 0.4842895, 0.480327, 0.4826861, 0.4913151, 0.4638297, 
    0.4779029, 0.4520208, 0.4595551, 0.4375417, 0.4484866, 0.4270416, 
    0.4179417, 0.4094219, 0.3995153, 0.4848347, 0.4878353, 0.4824653, 
    0.4750497, 0.4681881, 0.4590919, 0.4582118, 0.456511, 0.4521119, 
    0.448419, 0.4559728, 0.4474943, 0.4794075, 0.4626119, 0.4889699, 
    0.4810072, 0.4754866, 0.4779077, 0.4653594, 0.4624101, 0.4505054, 
    0.4566785, 0.420183, 0.4362517, 0.3920155, 0.4042633, 0.4888842, 
    0.4848454, 0.4708292, 0.4774899, 0.4585347, 0.4538759, 0.4500959, 
    0.4452717, 0.4447519, 0.4418992, 0.4465757, 0.442084, 0.4590726, 
    0.4514925, 0.4724287, 0.467306, 0.4696617, 0.4722474, 0.4642747, 
    0.4558536, 0.4556739, 0.4529635, 0.4453404, 0.4584579, 0.4181168, 
    0.4429389, 0.4804471, 0.4726922, 0.4715876, 0.4745877, 0.4543425, 
    0.4616299, 0.4419689, 0.4472799, 0.4385849, 0.4429012, 0.4435369, 
    0.4490948, 0.4525616, 0.461293, 0.4684573, 0.4741525, 0.4728273, 
    0.4665749, 0.4553365, 0.4447044, 0.4470291, 0.4392445, 0.4598595, 
    0.4512209, 0.4545746, 0.4458401, 0.46497, 0.4486744, 0.469163, 0.4673564, 
    0.4617757, 0.450632, 0.4481642, 0.4455302, 0.4471554, 0.4550508, 
    0.4563473, 0.4619115, 0.4634626, 0.4677497, 0.4713037, 0.4680561, 
    0.4646495, 0.4550479, 0.4463811, 0.4369701, 0.4346738, 0.4237412, 
    0.4326347, 0.4179792, 0.4304299, 0.4089315, 0.4477321, 0.4307994, 
    0.4615225, 0.4582377, 0.4522166, 0.4384679, 0.4458811, 0.4372145, 
    0.4563981, 0.4663589, 0.468956, 0.4738058, 0.4688452, 0.4692484, 
    0.4645093, 0.4660313, 0.454728, 0.4607717, 0.4435526, 0.4372831, 
    0.419682, 0.4089726, 0.3981415, 0.3933825, 0.391937, 0.3913331,
  0.05040628, 0.04850324, 0.04886981, 0.04735983, 0.048194, 0.0472103, 
    0.05001701, 0.04842852, 0.04943908, 0.05023328, 0.04451053, 0.04729315, 
    0.04172918, 0.04342415, 0.03924534, 0.04199011, 0.03870589, 0.03932309, 
    0.03748433, 0.03800546, 0.03571343, 0.03724533, 0.03456097, 0.03607566, 
    0.03583591, 0.03729654, 0.04672511, 0.04485133, 0.04683755, 0.04656712, 
    0.04668839, 0.04817662, 0.04893714, 0.05055367, 0.0502579, 0.0490718, 
    0.04644583, 0.0473276, 0.04512487, 0.04517392, 0.04279472, 0.0438577, 
    0.03997656, 0.04105711, 0.03798362, 0.0387425, 0.03801903, 0.03823752, 
    0.03801619, 0.03913299, 0.03865201, 0.03964392, 0.04365737, 0.04245295, 
    0.04610625, 0.04839146, 0.04994666, 0.05106796, 0.05090854, 0.05060541, 
    0.0490649, 0.04764261, 0.04657554, 0.04586986, 0.04518097, 0.04313387, 
    0.04207425, 0.03976016, 0.04017192, 0.03947603, 0.03881852, 0.03772992, 
    0.03790778, 0.03743291, 0.03949441, 0.03811654, 0.04040762, 0.03977266, 
    0.04499415, 0.04708876, 0.04799601, 0.0487992, 0.05078616, 0.04940891, 
    0.04994912, 0.04866982, 0.04786716, 0.04826317, 0.04585066, 0.04677968, 
    0.04201195, 0.04402721, 0.03889485, 0.0400872, 0.03861241, 0.03936068, 
    0.03808402, 0.03923182, 0.03725718, 0.03683562, 0.03712336, 0.03602596, 
    0.03929606, 0.03801898, 0.04827426, 0.04820953, 0.04790872, 0.04923946, 
    0.04932161, 0.05056176, 0.04945743, 0.04899153, 0.04782093, 0.0471364, 
    0.04649125, 0.04509166, 0.04355915, 0.04147061, 0.04000923, 0.03904781, 
    0.03963565, 0.03911638, 0.03969712, 0.03997118, 0.03699318, 0.0386475, 
    0.03618252, 0.03631626, 0.03742164, 0.03630118, 0.04816412, 0.04853711, 
    0.04984532, 0.04881976, 0.05069793, 0.04964132, 0.04903974, 0.04676, 
    0.04626803, 0.04581446, 0.04492675, 0.0438029, 0.04187335, 0.04023803, 
    0.0387805, 0.03888616, 0.03884894, 0.0385275, 0.03932669, 0.03839729, 
    0.03824261, 0.03864777, 0.03633419, 0.03698599, 0.03631911, 0.03674256, 
    0.04841569, 0.04779005, 0.04812751, 0.04749408, 0.04793976, 0.04597707, 
    0.04539828, 0.0427493, 0.04382482, 0.042121, 0.0436499, 0.04337651, 
    0.04206587, 0.04356646, 0.04032703, 0.04250615, 0.03851504, 0.04063014, 
    0.03838484, 0.03878673, 0.03812281, 0.03753423, 0.03680206, 0.0354748, 
    0.03577942, 0.03468728, 0.04686649, 0.04607169, 0.04614145, 0.04531783, 
    0.04471448, 0.04342379, 0.04140183, 0.04215524, 0.04077867, 0.04050568, 
    0.04259964, 0.04130613, 0.04554445, 0.04484236, 0.04525967, 0.04680342, 
    0.04198072, 0.04441566, 0.03998533, 0.04125536, 0.03761778, 0.03940049, 
    0.03594779, 0.03453223, 0.03323349, 0.03175559, 0.04564152, 0.04617761, 
    0.04522052, 0.04391618, 0.04272714, 0.04117716, 0.04102064, 0.04073484, 
    0.04000045, 0.03938936, 0.04064463, 0.0392371, 0.04468024, 0.0417734, 
    0.04638116, 0.04496247, 0.04399248, 0.04441651, 0.04224192, 0.0417391, 
    0.03973401, 0.04076294, 0.03487814, 0.0374105, 0.03065969, 0.0324596, 
    0.04636578, 0.04564342, 0.04318278, 0.04434318, 0.04107502, 0.04029411, 
    0.03966624, 0.03887239, 0.03878737, 0.03832241, 0.03908616, 0.03835244, 
    0.0411739, 0.03989762, 0.04345997, 0.0425755, 0.04298104, 0.04342851, 
    0.04205662, 0.04062464, 0.04059457, 0.04014208, 0.03888363, 0.04106209, 
    0.03455918, 0.03849152, 0.04486354, 0.04350572, 0.04331409, 0.04383559, 
    0.04037197, 0.04160662, 0.03833372, 0.03920184, 0.03778586, 0.03848539, 
    0.03858897, 0.03950082, 0.04007521, 0.04154947, 0.04277346, 0.04375974, 
    0.04352919, 0.04245006, 0.04053809, 0.03877959, 0.03916061, 0.03789233, 
    0.0413068, 0.03985256, 0.04041073, 0.03896549, 0.04217534, 0.03943145, 
    0.04289503, 0.04258417, 0.04163136, 0.03975498, 0.03934737, 0.03891472, 
    0.03918137, 0.0404903, 0.04070738, 0.04165441, 0.04191817, 0.04265174, 
    0.04326492, 0.04270442, 0.0421206, 0.04048982, 0.03905421, 0.03752587, 
    0.03715775, 0.03543098, 0.03683246, 0.03453799, 0.03648238, 0.03315951, 
    0.03927622, 0.03654094, 0.04158838, 0.041025, 0.04001786, 0.03776699, 
    0.03897221, 0.03756515, 0.04071591, 0.04241303, 0.04285934, 0.04369935, 
    0.04284026, 0.04290975, 0.04209666, 0.04235691, 0.04043636, 0.04146114, 
    0.03859153, 0.03757618, 0.03480067, 0.03316571, 0.03155337, 0.03085798, 
    0.03064834, 0.03056096,
  0.001354541, 0.001276427, 0.00129135, 0.001230264, 0.001263885, 
    0.001224271, 0.001338433, 0.001273393, 0.001314642, 0.001347375, 
    0.001117799, 0.00122759, 0.001011639, 0.001075901, 0.0009199581, 
    0.001021443, 0.0009004451, 0.0009227821, 0.0008567958, 0.0008753258, 
    0.0007948591, 0.0008483437, 0.0007559627, 0.0008073972, 0.000799091, 
    0.0008501522, 0.001204892, 0.001131055, 0.001209373, 0.001198604, 
    0.001203429, 0.001263181, 0.001294097, 0.001360657, 0.001348393, 
    0.001299598, 0.001193785, 0.001228972, 0.001141734, 0.001143652, 
    0.001051879, 0.001092555, 0.0009466362, 0.0009865371, 0.0008745465, 
    0.0009017648, 0.00087581, 0.000883621, 0.0008757086, 0.0009158824, 
    0.0008985042, 0.0009344674, 0.001084849, 0.001038913, 0.001180329, 
    0.001271888, 0.001335529, 0.001382072, 0.001375422, 0.001362807, 
    0.001299316, 0.001241627, 0.001198939, 0.001170992, 0.001143928, 
    0.001064799, 0.001024611, 0.0009387134, 0.0009538082, 0.0009283462, 
    0.0009045072, 0.0008655114, 0.0008718422, 0.0008549747, 0.0009290155, 
    0.0008792932, 0.0009624856, 0.0009391705, 0.001136626, 0.001219406, 
    0.001255877, 0.001288471, 0.001370323, 0.001313403, 0.001335631, 
    0.001283201, 0.001250675, 0.001266686, 0.001170235, 0.001207066, 
    0.001022265, 0.001099091, 0.0009072638, 0.0009506958, 0.0008970789, 
    0.0009241486, 0.0008781309, 0.000919467, 0.0008487618, 0.0008339214, 
    0.0008440411, 0.000805673, 0.0009217998, 0.0008758081, 0.001267136, 
    0.001264514, 0.001252352, 0.001306458, 0.001309824, 0.001360993, 
    0.001315395, 0.001296318, 0.00124881, 0.001221312, 0.001195589, 
    0.001140435, 0.001081077, 0.001001956, 0.000947834, 0.0009127964, 
    0.0009341654, 0.0009152801, 0.0009364098, 0.0009464387, 0.0008394576, 
    0.0008983421, 0.0008111089, 0.0008157627, 0.0008545758, 0.0008152373, 
    0.001262675, 0.001277803, 0.00133135, 0.001289309, 0.001366652, 
    0.001322951, 0.001298287, 0.001206282, 0.001186733, 0.001168807, 
    0.001133996, 0.001090445, 0.001017052, 0.0009562395, 0.0009031354, 
    0.00090695, 0.0009056056, 0.0008940246, 0.0009229131, 0.0008893476, 
    0.0008838032, 0.0008983517, 0.0008163874, 0.0008392046, 0.0008158618, 
    0.0008306577, 0.001272872, 0.001247565, 0.001261193, 0.001235654, 
    0.001253605, 0.001175223, 0.001152442, 0.001050152, 0.001091289, 
    0.001026373, 0.001084562, 0.001074076, 0.001024295, 0.001081358, 
    0.0009595158, 0.001040928, 0.0008935767, 0.0009707026, 0.000888901, 
    0.0009033602, 0.0008795172, 0.0008585644, 0.000832744, 0.0007866365, 
    0.0007971383, 0.0007597108, 0.001210528, 0.001178962, 0.001181721, 
    0.001149287, 0.001125725, 0.001075887, 0.0009993854, 0.001027664, 
    0.000976201, 0.0009661039, 0.001044471, 0.0009958129, 0.001158181, 
    0.001130705, 0.001147009, 0.001208012, 0.00102109, 0.001114118, 
    0.0009469574, 0.0009939192, 0.0008615282, 0.0009255964, 0.0008029634, 
    0.000754985, 0.0007112788, 0.0006626702, 0.001161997, 0.001183152, 
    0.001145476, 0.001094809, 0.00104931, 0.0009910053, 0.0009851812, 
    0.0009745777, 0.0009475123, 0.0009251917, 0.0009712387, 0.0009196589, 
    0.001124393, 0.001013298, 0.001191219, 0.001135389, 0.001097751, 
    0.001114151, 0.001030935, 0.001012011, 0.0009377578, 0.0009756184, 
    0.0007662065, 0.0008541816, 0.000627417, 0.0006856741, 0.001190608, 
    0.001162072, 0.001066667, 0.001111309, 0.0009872032, 0.0009583032, 
    0.0009352822, 0.0009064527, 0.0009033834, 0.000886662, 0.0009141852, 
    0.0008877388, 0.0009908838, 0.0009437436, 0.001077273, 0.001043556, 
    0.00105897, 0.001076068, 0.001023947, 0.0009704996, 0.0009693877, 
    0.0009527113, 0.0009068585, 0.0009867225, 0.0007559016, 0.0008927312, 
    0.001131531, 0.001079027, 0.001071687, 0.001091704, 0.0009611716, 
    0.001007045, 0.0008870677, 0.0009183791, 0.0008675007, 0.0008925109, 
    0.0008962353, 0.0009292493, 0.0009502555, 0.001004906, 0.00105107, 
    0.001088785, 0.001079928, 0.001038803, 0.0009673008, 0.0009031028, 
    0.0009168838, 0.0008712914, 0.0009958379, 0.0009420936, 0.0009626005, 
    0.0009098174, 0.001028422, 0.0009267229, 0.001055694, 0.001043884, 
    0.001007972, 0.000938524, 0.0009236647, 0.0009079818, 0.0009176366, 
    0.000965536, 0.0009735608, 0.001008836, 0.001018737, 0.001046448, 
    0.001069806, 0.001048448, 0.001026358, 0.0009655182, 0.0009130281, 
    0.0008582679, 0.0008452536, 0.0007851296, 0.0008338105, 0.0007551811, 
    0.0008215555, 0.0007088167, 0.0009210792, 0.0008236012, 0.001006362, 
    0.0009853432, 0.0009481508, 0.0008668294, 0.0009100605, 0.0008596606, 
    0.0009738768, 0.001037402, 0.001054336, 0.001086462, 0.00105361, 
    0.001056254, 0.001025455, 0.001035279, 0.0009635456, 0.001001602, 
    0.0008963273, 0.0008600518, 0.0007635675, 0.0007090232, 0.0006561142, 
    0.000633745, 0.0006270552, 0.0006242746,
  8.907525e-06, 8.124078e-06, 8.271951e-06, 7.672144e-06, 8.000459e-06, 
    7.614086e-06, 8.744089e-06, 8.094114e-06, 8.504464e-06, 8.83469e-06, 
    6.607359e-06, 7.646226e-06, 5.65255e-06, 6.224465e-06, 4.870592e-06, 
    5.738569e-06, 4.709588e-06, 4.894056e-06, 4.35666e-06, 4.505247e-06, 
    3.873724e-06, 4.289502e-06, 3.248501e-06, 3.969742e-06, 3.906031e-06, 
    4.303838e-06, 7.427363e-06, 6.730099e-06, 7.470408e-06, 7.367109e-06, 
    7.413334e-06, 7.99354e-06, 8.299265e-06, 8.96983e-06, 8.845032e-06, 
    8.354047e-06, 7.321034e-06, 7.659612e-06, 6.829529e-06, 6.847441e-06, 
    6.00846e-06, 6.37574e-06, 5.093857e-06, 5.434381e-06, 4.498962e-06, 
    4.720416e-06, 4.509155e-06, 4.57236e-06, 4.508337e-06, 4.836801e-06, 
    4.693681e-06, 4.991574e-06, 6.305588e-06, 5.892963e-06, 7.192884e-06, 
    8.079272e-06, 8.714727e-06, 9.189079e-06, 9.12081e-06, 8.99176e-06, 
    8.351239e-06, 7.7826e-06, 7.370311e-06, 7.104411e-06, 6.850019e-06, 
    6.124316e-06, 5.766466e-06, 5.027179e-06, 5.154488e-06, 4.940404e-06, 
    4.742943e-06, 4.426318e-06, 4.477173e-06, 4.342157e-06, 4.945989e-06, 
    4.5373e-06, 5.228185e-06, 5.031017e-06, 6.781911e-06, 7.567075e-06, 
    7.921853e-06, 8.243352e-06, 9.068588e-06, 8.49205e-06, 8.715753e-06, 
    8.191094e-06, 7.870926e-06, 8.028019e-06, 7.09725e-06, 7.448236e-06, 
    5.745805e-06, 6.435438e-06, 4.765627e-06, 5.128145e-06, 4.682013e-06, 
    4.905424e-06, 4.527901e-06, 4.866517e-06, 4.292815e-06, 4.175809e-06, 
    4.255463e-06, 3.956485e-06, 4.885889e-06, 4.50914e-06, 8.032443e-06, 
    8.006641e-06, 7.887331e-06, 8.42253e-06, 8.456197e-06, 8.973257e-06, 
    8.512017e-06, 8.321373e-06, 7.852698e-06, 7.585484e-06, 7.338268e-06, 
    6.81741e-06, 6.271353e-06, 5.568036e-06, 5.103966e-06, 4.811272e-06, 
    4.989044e-06, 4.831816e-06, 5.00785e-06, 5.092192e-06, 4.219316e-06, 
    4.692354e-06, 3.99834e-06, 4.034306e-06, 4.338983e-06, 4.030239e-06, 
    7.988567e-06, 8.137678e-06, 8.672527e-06, 8.251673e-06, 9.031042e-06, 
    8.587906e-06, 8.340987e-06, 7.440707e-06, 7.253782e-06, 7.083761e-06, 
    6.757435e-06, 6.356508e-06, 5.699987e-06, 5.175099e-06, 4.73167e-06, 
    4.763043e-06, 4.751977e-06, 4.657043e-06, 4.895146e-06, 4.618903e-06, 
    4.573838e-06, 4.692432e-06, 4.039143e-06, 4.217324e-06, 4.035073e-06, 
    4.150241e-06, 8.088975e-06, 7.840534e-06, 7.974012e-06, 7.724479e-06, 
    7.899597e-06, 7.14446e-06, 6.929711e-06, 5.993036e-06, 6.364197e-06, 
    5.781998e-06, 6.302982e-06, 6.207967e-06, 5.763682e-06, 6.273898e-06, 
    5.202921e-06, 5.910861e-06, 4.653386e-06, 5.298314e-06, 4.615267e-06, 
    4.733516e-06, 4.539112e-06, 4.370762e-06, 4.166578e-06, 3.811247e-06, 
    3.891111e-06, 3.609435e-06, 7.481511e-06, 7.17991e-06, 7.206111e-06, 
    6.900148e-06, 6.680661e-06, 6.224343e-06, 5.545676e-06, 5.79339e-06, 
    5.345424e-06, 5.259025e-06, 5.942383e-06, 5.514651e-06, 6.983605e-06, 
    6.726855e-06, 6.878821e-06, 7.457329e-06, 5.735463e-06, 6.573415e-06, 
    5.096568e-06, 5.49823e-06, 4.394432e-06, 4.917479e-06, 3.935685e-06, 
    3.243093e-06, 3.002659e-06, 2.738317e-06, 7.019518e-06, 7.219709e-06, 
    6.864482e-06, 6.396303e-06, 5.98552e-06, 5.472996e-06, 5.422683e-06, 
    5.3315e-06, 5.101251e-06, 4.914108e-06, 5.3029e-06, 4.868109e-06, 
    6.668325e-06, 5.667076e-06, 7.296534e-06, 6.770399e-06, 6.423182e-06, 
    6.573719e-06, 5.822281e-06, 5.655807e-06, 5.019157e-06, 5.340425e-06, 
    3.657727e-06, 4.335847e-06, 2.548768e-06, 2.863e-06, 7.290713e-06, 
    7.020222e-06, 6.141128e-06, 6.547547e-06, 5.440131e-06, 5.192618e-06, 
    4.998399e-06, 4.758948e-06, 4.733707e-06, 4.597054e-06, 4.822756e-06, 
    4.60581e-06, 5.471945e-06, 5.069477e-06, 6.236886e-06, 5.934232e-06, 
    6.071954e-06, 6.225976e-06, 5.760614e-06, 5.296577e-06, 5.287069e-06, 
    5.145198e-06, 4.762289e-06, 5.435981e-06, 3.248163e-06, 4.646484e-06, 
    6.734524e-06, 6.252771e-06, 6.186386e-06, 6.367979e-06, 5.217001e-06, 
    5.612401e-06, 4.600352e-06, 4.857491e-06, 4.442275e-06, 4.644687e-06, 
    4.675111e-06, 4.947941e-06, 5.124422e-06, 5.593734e-06, 6.001238e-06, 
    6.341385e-06, 6.260931e-06, 5.891992e-06, 5.269241e-06, 4.731402e-06, 
    4.845096e-06, 4.47274e-06, 5.514867e-06, 5.055588e-06, 5.229163e-06, 
    4.786675e-06, 5.800081e-06, 4.926866e-06, 6.042597e-06, 5.937157e-06, 
    5.620494e-06, 5.025588e-06, 4.901397e-06, 4.771542e-06, 4.851335e-06, 
    5.25418e-06, 5.322785e-06, 5.628037e-06, 5.714781e-06, 5.959989e-06, 
    6.169417e-06, 5.977823e-06, 5.781864e-06, 5.254029e-06, 4.813188e-06, 
    4.368397e-06, 4.265046e-06, 3.799839e-06, 4.174939e-06, 3.244178e-06, 
    4.079246e-06, 2.989191e-06, 4.879902e-06, 4.095161e-06, 5.606442e-06, 
    5.42408e-06, 5.10664e-06, 4.436888e-06, 4.788681e-06, 4.379511e-06, 
    5.325492e-06, 5.879555e-06, 6.030439e-06, 6.320255e-06, 6.023942e-06, 
    6.047614e-06, 5.773907e-06, 5.860737e-06, 5.237213e-06, 5.564953e-06, 
    4.675864e-06, 4.382635e-06, 3.638077e-06, 2.99032e-06, 2.702925e-06, 
    2.582652e-06, 2.546833e-06, 2.531965e-06,
  8.171996e-09, 6.972882e-09, 7.196181e-09, 6.299846e-09, 6.787351e-09, 
    6.214457e-09, 7.918669e-09, 6.927814e-09, 7.550212e-09, 8.058903e-09, 
    4.776886e-09, 6.261695e-09, 3.501305e-09, 4.253918e-09, 2.537116e-09, 
    3.612149e-09, 2.349386e-09, 2.564807e-09, 1.95272e-09, 2.117129e-09, 
    1.447282e-09, 1.879713e-09, 1.159808e-09, 1.544e-09, 1.479603e-09, 
    1.895228e-09, 5.941565e-09, 4.94749e-09, 6.004238e-09, 5.85408e-09, 
    5.92117e-09, 6.776997e-09, 7.237587e-09, 8.268988e-09, 8.074941e-09, 
    7.320782e-09, 5.787377e-09, 6.281394e-09, 5.086699e-09, 5.111871e-09, 
    3.965442e-09, 4.458814e-09, 2.803901e-09, 3.224184e-09, 2.110096e-09, 
    2.361883e-09, 2.121505e-09, 2.192643e-09, 2.120588e-09, 2.497383e-09, 
    2.33106e-09, 2.680776e-09, 4.363509e-09, 3.813254e-09, 5.602748e-09, 
    6.905515e-09, 7.873331e-09, 8.612102e-09, 8.504968e-09, 8.303183e-09, 
    7.316511e-09, 6.46299e-09, 5.858723e-09, 5.476064e-09, 5.115496e-09, 
    4.119557e-09, 3.648283e-09, 2.723466e-09, 2.877585e-09, 2.619749e-09, 
    2.387944e-09, 2.02931e-09, 2.085768e-09, 1.936884e-09, 2.626392e-09, 
    2.153099e-09, 2.967832e-09, 2.728078e-09, 5.01992e-09, 6.1455e-09, 
    6.669929e-09, 7.15288e-09, 8.423196e-09, 7.531222e-09, 7.874913e-09, 
    7.0739e-09, 6.594088e-09, 6.828622e-09, 5.46584e-09, 5.971938e-09, 
    3.621513e-09, 4.540298e-09, 2.414268e-09, 2.845507e-09, 2.317643e-09, 
    2.578253e-09, 2.142533e-09, 2.532314e-09, 1.883294e-09, 1.758042e-09, 
    1.843029e-09, 1.530529e-09, 2.55516e-09, 2.121488e-09, 6.835254e-09, 
    6.796605e-09, 6.618497e-09, 7.425058e-09, 7.476432e-09, 8.274331e-09, 
    7.561773e-09, 7.271137e-09, 6.566987e-09, 6.172483e-09, 5.812308e-09, 
    5.069684e-09, 4.317178e-09, 3.393259e-09, 2.81615e-09, 2.46748e-09, 
    2.677751e-09, 2.491535e-09, 2.700269e-09, 2.801884e-09, 1.804311e-09, 
    2.329532e-09, 1.573186e-09, 1.610133e-09, 1.933423e-09, 1.605942e-09, 
    6.769559e-09, 6.993359e-09, 7.80826e-09, 7.165474e-09, 8.364503e-09, 
    7.67811e-09, 7.300931e-09, 5.960978e-09, 5.69032e-09, 5.44659e-09, 
    4.985673e-09, 4.432637e-09, 3.562325e-09, 2.90275e-09, 2.374892e-09, 
    2.411265e-09, 2.398417e-09, 2.289005e-09, 2.566095e-09, 2.245459e-09, 
    2.194315e-09, 2.329623e-09, 1.615122e-09, 1.802185e-09, 1.610924e-09, 
    1.731022e-09, 6.920092e-09, 6.548914e-09, 6.747795e-09, 6.377032e-09, 
    6.636762e-09, 5.53333e-09, 5.22785e-09, 3.945033e-09, 4.443099e-09, 
    3.668442e-09, 4.359978e-09, 4.231712e-09, 3.644673e-09, 4.320619e-09, 
    2.93681e-09, 3.836742e-09, 2.284819e-09, 3.054391e-09, 2.241319e-09, 
    2.377029e-09, 2.155137e-09, 1.968155e-09, 1.748272e-09, 1.385431e-09, 
    1.464648e-09, 1.191778e-09, 6.020425e-09, 5.584129e-09, 5.621742e-09, 
    5.186106e-09, 4.878607e-09, 4.253754e-09, 3.36482e-09, 3.683244e-09, 
    3.112906e-09, 3.005817e-09, 3.878193e-09, 3.32546e-09, 5.304144e-09, 
    4.942962e-09, 5.156038e-09, 5.985179e-09, 3.608132e-09, 4.729951e-09, 
    2.807184e-09, 3.304676e-09, 1.994143e-09, 2.592533e-09, 1.509468e-09, 
    1.153147e-09, 8.742308e-10, 6.085719e-10, 5.355124e-09, 5.641284e-09, 
    5.135846e-09, 4.486842e-09, 3.935098e-09, 3.272803e-09, 3.209492e-09, 
    3.095581e-09, 2.812858e-09, 2.588538e-09, 3.060075e-09, 2.53419e-09, 
    4.861453e-09, 3.519962e-09, 5.751978e-09, 5.003805e-09, 4.523542e-09, 
    4.730373e-09, 3.720851e-09, 3.505486e-09, 2.713832e-09, 3.106683e-09, 
    1.237238e-09, 1.930006e-09, 4.463162e-10, 7.283277e-10, 5.743573e-09, 
    5.356124e-09, 4.142039e-09, 4.694257e-09, 3.231412e-09, 2.924185e-09, 
    2.688946e-09, 2.406508e-09, 2.377249e-09, 2.220621e-09, 2.480919e-09, 
    2.230564e-09, 3.271477e-09, 2.774417e-09, 4.270655e-09, 3.867464e-09, 
    4.049725e-09, 4.255954e-09, 3.640697e-09, 3.05224e-09, 3.040469e-09, 
    2.866262e-09, 2.410388e-09, 3.226195e-09, 1.159391e-09, 2.276925e-09, 
    4.953666e-09, 4.292082e-09, 4.202708e-09, 4.448245e-09, 2.954089e-09, 
    3.44987e-09, 2.224365e-09, 2.52169e-09, 2.046976e-09, 2.274871e-09, 
    2.309717e-09, 2.628714e-09, 2.840982e-09, 3.426022e-09, 3.955883e-09, 
    4.412079e-09, 4.303099e-09, 3.811981e-09, 3.018427e-09, 2.374582e-09, 
    2.507119e-09, 2.080829e-09, 3.325734e-09, 2.757659e-09, 2.969034e-09, 
    2.438765e-09, 3.691945e-09, 2.603667e-09, 4.010703e-09, 3.871314e-09, 
    3.460222e-09, 2.721554e-09, 2.573488e-09, 2.421145e-09, 2.514451e-09, 
    2.999841e-09, 3.08475e-09, 3.469878e-09, 3.581409e-09, 3.901394e-09, 
    4.179936e-09, 3.924929e-09, 3.668268e-09, 2.999654e-09, 2.469721e-09, 
    1.965564e-09, 1.853334e-09, 1.374232e-09, 1.757121e-09, 1.154481e-09, 
    1.656672e-09, 8.596317e-10, 2.548094e-09, 1.673252e-09, 3.442252e-09, 
    3.211247e-09, 2.819393e-09, 2.041007e-09, 2.441103e-09, 1.97775e-09, 
    3.088114e-09, 3.795682e-09, 3.994569e-09, 4.383394e-09, 3.985954e-09, 
    4.017365e-09, 3.657938e-09, 3.771055e-09, 2.978938e-09, 3.389336e-09, 
    2.310581e-09, 1.981179e-09, 1.218672e-09, 8.608514e-10, 5.76435e-10, 
    4.735225e-10, 4.447866e-10, 4.331206e-10,
  4.330856e-13, 4.283784e-13, 4.292556e-13, 4.257326e-13, 4.276493e-13, 
    4.253967e-13, 4.320918e-13, 4.282013e-13, 4.306457e-13, 4.326419e-13, 
    4.197344e-13, 4.255825e-13, 4.146965e-13, 4.176706e-13, 4.108788e-13, 
    4.151349e-13, 4.101342e-13, 4.109886e-13, 4.085595e-13, 4.092125e-13, 
    4.065496e-13, 4.082694e-13, 4.0541e-13, 4.069345e-13, 4.066782e-13, 
    4.083311e-13, 4.24323e-13, 4.204072e-13, 4.245696e-13, 4.239786e-13, 
    4.242427e-13, 4.276086e-13, 4.294182e-13, 4.33466e-13, 4.327049e-13, 
    4.297449e-13, 4.23716e-13, 4.2566e-13, 4.20956e-13, 4.210552e-13, 
    4.165313e-13, 4.184795e-13, 4.119361e-13, 4.136002e-13, 4.091845e-13, 
    4.101838e-13, 4.092298e-13, 4.095122e-13, 4.092262e-13, 4.107212e-13, 
    4.100615e-13, 4.114482e-13, 4.181033e-13, 4.159299e-13, 4.229891e-13, 
    4.281137e-13, 4.319139e-13, 4.348112e-13, 4.343912e-13, 4.336e-13, 
    4.297281e-13, 4.263742e-13, 4.239969e-13, 4.224902e-13, 4.210695e-13, 
    4.171401e-13, 4.152777e-13, 4.116174e-13, 4.12228e-13, 4.112064e-13, 
    4.102872e-13, 4.088637e-13, 4.090879e-13, 4.084966e-13, 4.112327e-13, 
    4.093552e-13, 4.125854e-13, 4.116357e-13, 4.206927e-13, 4.251254e-13, 
    4.271878e-13, 4.290855e-13, 4.340706e-13, 4.305712e-13, 4.319201e-13, 
    4.287752e-13, 4.268896e-13, 4.278115e-13, 4.224499e-13, 4.244425e-13, 
    4.151719e-13, 4.18801e-13, 4.103916e-13, 4.121009e-13, 4.100083e-13, 
    4.110419e-13, 4.093133e-13, 4.108597e-13, 4.082836e-13, 4.077858e-13, 
    4.081236e-13, 4.068809e-13, 4.109503e-13, 4.092298e-13, 4.278376e-13, 
    4.276857e-13, 4.269856e-13, 4.301544e-13, 4.303561e-13, 4.334869e-13, 
    4.306911e-13, 4.2955e-13, 4.267831e-13, 4.252316e-13, 4.238142e-13, 
    4.208889e-13, 4.179204e-13, 4.142691e-13, 4.119847e-13, 4.106026e-13, 
    4.114363e-13, 4.106981e-13, 4.115255e-13, 4.119281e-13, 4.079697e-13, 
    4.100555e-13, 4.070506e-13, 4.071976e-13, 4.084828e-13, 4.07181e-13, 
    4.275794e-13, 4.284588e-13, 4.316585e-13, 4.291349e-13, 4.338405e-13, 
    4.311478e-13, 4.29667e-13, 4.243993e-13, 4.233339e-13, 4.223741e-13, 
    4.205577e-13, 4.183762e-13, 4.149378e-13, 4.123277e-13, 4.102354e-13, 
    4.103797e-13, 4.103288e-13, 4.098947e-13, 4.109937e-13, 4.097219e-13, 
    4.095189e-13, 4.100558e-13, 4.072175e-13, 4.079613e-13, 4.072008e-13, 
    4.076784e-13, 4.28171e-13, 4.26712e-13, 4.274938e-13, 4.260362e-13, 
    4.270574e-13, 4.227157e-13, 4.215123e-13, 4.164506e-13, 4.184174e-13, 
    4.153574e-13, 4.180894e-13, 4.17583e-13, 4.152635e-13, 4.17934e-13, 
    4.124626e-13, 4.160227e-13, 4.098781e-13, 4.129281e-13, 4.097054e-13, 
    4.102439e-13, 4.093634e-13, 4.086208e-13, 4.07747e-13, 4.063034e-13, 
    4.066187e-13, 4.05532e-13, 4.246333e-13, 4.229158e-13, 4.230639e-13, 
    4.213477e-13, 4.201356e-13, 4.1767e-13, 4.141566e-13, 4.15416e-13, 
    4.131598e-13, 4.127358e-13, 4.161865e-13, 4.140009e-13, 4.218129e-13, 
    4.203893e-13, 4.212293e-13, 4.244946e-13, 4.15119e-13, 4.195493e-13, 
    4.119491e-13, 4.139186e-13, 4.087241e-13, 4.110985e-13, 4.067971e-13, 
    4.053835e-13, 4.042697e-13, 4.032074e-13, 4.220137e-13, 4.231409e-13, 
    4.211497e-13, 4.185901e-13, 4.164114e-13, 4.137925e-13, 4.13542e-13, 
    4.130912e-13, 4.119716e-13, 4.110827e-13, 4.129506e-13, 4.108672e-13, 
    4.200679e-13, 4.147703e-13, 4.235767e-13, 4.206292e-13, 4.187349e-13, 
    4.195509e-13, 4.155646e-13, 4.147131e-13, 4.115792e-13, 4.131351e-13, 
    4.057131e-13, 4.084693e-13, 4.025578e-13, 4.036865e-13, 4.235436e-13, 
    4.220177e-13, 4.172288e-13, 4.194085e-13, 4.136288e-13, 4.124126e-13, 
    4.114806e-13, 4.103608e-13, 4.102448e-13, 4.096233e-13, 4.10656e-13, 
    4.096628e-13, 4.137873e-13, 4.118193e-13, 4.177367e-13, 4.161441e-13, 
    4.168642e-13, 4.176787e-13, 4.152478e-13, 4.129196e-13, 4.12873e-13, 
    4.121832e-13, 4.103762e-13, 4.136081e-13, 4.054084e-13, 4.098467e-13, 
    4.204315e-13, 4.178213e-13, 4.174684e-13, 4.184378e-13, 4.12531e-13, 
    4.144931e-13, 4.096381e-13, 4.108176e-13, 4.089339e-13, 4.098386e-13, 
    4.099768e-13, 4.112419e-13, 4.12083e-13, 4.143987e-13, 4.164935e-13, 
    4.18295e-13, 4.178648e-13, 4.159248e-13, 4.127857e-13, 4.102342e-13, 
    4.107599e-13, 4.090683e-13, 4.140019e-13, 4.117529e-13, 4.125902e-13, 
    4.104888e-13, 4.154504e-13, 4.111426e-13, 4.167101e-13, 4.161593e-13, 
    4.14534e-13, 4.116098e-13, 4.11023e-13, 4.104189e-13, 4.107889e-13, 
    4.127122e-13, 4.130483e-13, 4.145722e-13, 4.150133e-13, 4.162782e-13, 
    4.173785e-13, 4.163712e-13, 4.153567e-13, 4.127114e-13, 4.106115e-13, 
    4.086105e-13, 4.081646e-13, 4.062588e-13, 4.077822e-13, 4.053888e-13, 
    4.073827e-13, 4.042114e-13, 4.109223e-13, 4.074487e-13, 4.144629e-13, 
    4.13549e-13, 4.119975e-13, 4.089102e-13, 4.104981e-13, 4.086589e-13, 
    4.130616e-13, 4.158604e-13, 4.166463e-13, 4.181818e-13, 4.166123e-13, 
    4.167364e-13, 4.153159e-13, 4.157631e-13, 4.126294e-13, 4.142536e-13, 
    4.099803e-13, 4.086726e-13, 4.056391e-13, 4.042163e-13, 4.030788e-13, 
    4.026668e-13, 4.025517e-13, 4.02505e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.94965e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949654e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949654e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949654e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.94965e-07, 8.949651e-07, 8.949648e-07, 8.94965e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.94965e-07, 8.949651e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.94965e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.010595e-16, 6.026879e-16, 6.023716e-16, 6.036837e-16, 6.029562e-16, 
    6.03815e-16, 6.0139e-16, 6.027522e-16, 6.018829e-16, 6.012065e-16, 
    6.062264e-16, 6.037423e-16, 6.088047e-16, 6.072232e-16, 6.111934e-16, 
    6.085583e-16, 6.117243e-16, 6.11118e-16, 6.129435e-16, 6.124208e-16, 
    6.147522e-16, 6.131848e-16, 6.159603e-16, 6.143784e-16, 6.146257e-16, 
    6.13133e-16, 6.04243e-16, 6.059171e-16, 6.041437e-16, 6.043825e-16, 
    6.042755e-16, 6.02971e-16, 6.023129e-16, 6.009354e-16, 6.011857e-16, 
    6.021975e-16, 6.044899e-16, 6.037125e-16, 6.056722e-16, 6.05628e-16, 
    6.078064e-16, 6.068246e-16, 6.104816e-16, 6.094435e-16, 6.124427e-16, 
    6.116888e-16, 6.124072e-16, 6.121894e-16, 6.1241e-16, 6.113042e-16, 
    6.117781e-16, 6.108049e-16, 6.070084e-16, 6.081251e-16, 6.04792e-16, 
    6.027836e-16, 6.014497e-16, 6.00502e-16, 6.00636e-16, 6.008914e-16, 
    6.022035e-16, 6.034366e-16, 6.043756e-16, 6.050033e-16, 6.056216e-16, 
    6.074902e-16, 6.084796e-16, 6.106913e-16, 6.102928e-16, 6.109681e-16, 
    6.116138e-16, 6.126965e-16, 6.125184e-16, 6.129951e-16, 6.109507e-16, 
    6.123095e-16, 6.10066e-16, 6.106796e-16, 6.057878e-16, 6.039224e-16, 
    6.031272e-16, 6.024323e-16, 6.00739e-16, 6.019084e-16, 6.014475e-16, 
    6.025443e-16, 6.032406e-16, 6.028963e-16, 6.050204e-16, 6.041949e-16, 
    6.085382e-16, 6.066689e-16, 6.115385e-16, 6.103746e-16, 6.118174e-16, 
    6.110814e-16, 6.123421e-16, 6.112076e-16, 6.131726e-16, 6.135999e-16, 
    6.133079e-16, 6.144301e-16, 6.111446e-16, 6.124069e-16, 6.028866e-16, 
    6.029427e-16, 6.032045e-16, 6.020536e-16, 6.019833e-16, 6.009284e-16, 
    6.018672e-16, 6.022667e-16, 6.032811e-16, 6.038804e-16, 6.044501e-16, 
    6.057019e-16, 6.070985e-16, 6.090498e-16, 6.104501e-16, 6.113882e-16, 
    6.108131e-16, 6.113208e-16, 6.107532e-16, 6.104872e-16, 6.134397e-16, 
    6.117824e-16, 6.142687e-16, 6.141313e-16, 6.130063e-16, 6.141468e-16, 
    6.029822e-16, 6.02659e-16, 6.01536e-16, 6.02415e-16, 6.008135e-16, 
    6.017099e-16, 6.022249e-16, 6.042117e-16, 6.046484e-16, 6.050526e-16, 
    6.05851e-16, 6.068749e-16, 6.086691e-16, 6.102286e-16, 6.116514e-16, 
    6.115473e-16, 6.115839e-16, 6.119014e-16, 6.111146e-16, 6.120305e-16, 
    6.12184e-16, 6.117824e-16, 6.141129e-16, 6.134475e-16, 6.141284e-16, 
    6.136952e-16, 6.027641e-16, 6.033078e-16, 6.03014e-16, 6.035664e-16, 
    6.031771e-16, 6.049068e-16, 6.05425e-16, 6.078481e-16, 6.068546e-16, 
    6.08436e-16, 6.070155e-16, 6.072671e-16, 6.084868e-16, 6.070924e-16, 
    6.101426e-16, 6.080746e-16, 6.119138e-16, 6.098505e-16, 6.120429e-16, 
    6.116452e-16, 6.123038e-16, 6.128931e-16, 6.136345e-16, 6.15001e-16, 
    6.146848e-16, 6.158272e-16, 6.041183e-16, 6.048227e-16, 6.047611e-16, 
    6.054982e-16, 6.060431e-16, 6.072238e-16, 6.091153e-16, 6.084044e-16, 
    6.097096e-16, 6.099714e-16, 6.079885e-16, 6.092059e-16, 6.052943e-16, 
    6.059266e-16, 6.055504e-16, 6.041737e-16, 6.085678e-16, 6.06314e-16, 
    6.104732e-16, 6.092545e-16, 6.12809e-16, 6.110418e-16, 6.145105e-16, 
    6.1599e-16, 6.173828e-16, 6.190068e-16, 6.052074e-16, 6.047289e-16, 
    6.055859e-16, 6.067704e-16, 6.078694e-16, 6.093289e-16, 6.094783e-16, 
    6.097514e-16, 6.104588e-16, 6.110534e-16, 6.098374e-16, 6.112024e-16, 
    6.060725e-16, 6.087634e-16, 6.045476e-16, 6.058178e-16, 6.067007e-16, 
    6.063139e-16, 6.083232e-16, 6.087963e-16, 6.107168e-16, 6.097247e-16, 
    6.156247e-16, 6.13017e-16, 6.202433e-16, 6.182272e-16, 6.045616e-16, 
    6.052059e-16, 6.074461e-16, 6.063807e-16, 6.094264e-16, 6.101751e-16, 
    6.107833e-16, 6.115604e-16, 6.116446e-16, 6.121048e-16, 6.113505e-16, 
    6.120752e-16, 6.093319e-16, 6.105583e-16, 6.071906e-16, 6.080108e-16, 
    6.076336e-16, 6.072196e-16, 6.084971e-16, 6.098565e-16, 6.098861e-16, 
    6.103213e-16, 6.115468e-16, 6.094388e-16, 6.159599e-16, 6.119347e-16, 
    6.059083e-16, 6.071474e-16, 6.07325e-16, 6.068451e-16, 6.101e-16, 
    6.089213e-16, 6.120936e-16, 6.11237e-16, 6.126406e-16, 6.119432e-16, 
    6.118405e-16, 6.109445e-16, 6.103862e-16, 6.089753e-16, 6.078262e-16, 
    6.069147e-16, 6.071268e-16, 6.081279e-16, 6.099397e-16, 6.116519e-16, 
    6.112768e-16, 6.125339e-16, 6.092057e-16, 6.106017e-16, 6.100624e-16, 
    6.11469e-16, 6.083854e-16, 6.110098e-16, 6.077135e-16, 6.08003e-16, 
    6.088979e-16, 6.10696e-16, 6.110944e-16, 6.115187e-16, 6.11257e-16, 
    6.099858e-16, 6.097776e-16, 6.088763e-16, 6.086271e-16, 6.0794e-16, 
    6.073707e-16, 6.078907e-16, 6.084365e-16, 6.099866e-16, 6.113814e-16, 
    6.129014e-16, 6.132733e-16, 6.150453e-16, 6.136022e-16, 6.159821e-16, 
    6.139577e-16, 6.174609e-16, 6.111626e-16, 6.138994e-16, 6.089388e-16, 
    6.094742e-16, 6.104411e-16, 6.126585e-16, 6.114623e-16, 6.128613e-16, 
    6.097695e-16, 6.081621e-16, 6.077467e-16, 6.0697e-16, 6.077644e-16, 
    6.076998e-16, 6.084596e-16, 6.082155e-16, 6.100381e-16, 6.090594e-16, 
    6.118378e-16, 6.128505e-16, 6.157072e-16, 6.174555e-16, 6.192339e-16, 
    6.20018e-16, 6.202567e-16, 6.203563e-16 ;

 CWDC_TO_LITR2C =
  4.568052e-16, 4.580428e-16, 4.578024e-16, 4.587996e-16, 4.582467e-16, 
    4.588994e-16, 4.570564e-16, 4.580917e-16, 4.57431e-16, 4.569169e-16, 
    4.60732e-16, 4.588441e-16, 4.626916e-16, 4.614896e-16, 4.64507e-16, 
    4.625043e-16, 4.649105e-16, 4.644497e-16, 4.658371e-16, 4.654398e-16, 
    4.672117e-16, 4.660204e-16, 4.681299e-16, 4.669275e-16, 4.671155e-16, 
    4.65981e-16, 4.592247e-16, 4.60497e-16, 4.591492e-16, 4.593307e-16, 
    4.592494e-16, 4.58258e-16, 4.577578e-16, 4.567109e-16, 4.569011e-16, 
    4.576701e-16, 4.594124e-16, 4.588215e-16, 4.603108e-16, 4.602773e-16, 
    4.619329e-16, 4.611867e-16, 4.639661e-16, 4.63177e-16, 4.654564e-16, 
    4.648834e-16, 4.654294e-16, 4.65264e-16, 4.654316e-16, 4.645912e-16, 
    4.649513e-16, 4.642117e-16, 4.613264e-16, 4.621751e-16, 4.59642e-16, 
    4.581156e-16, 4.571018e-16, 4.563815e-16, 4.564834e-16, 4.566774e-16, 
    4.576746e-16, 4.586119e-16, 4.593254e-16, 4.598025e-16, 4.602724e-16, 
    4.616926e-16, 4.624445e-16, 4.641254e-16, 4.638225e-16, 4.643358e-16, 
    4.648265e-16, 4.656493e-16, 4.65514e-16, 4.658763e-16, 4.643226e-16, 
    4.653552e-16, 4.636502e-16, 4.641165e-16, 4.603987e-16, 4.58981e-16, 
    4.583767e-16, 4.578485e-16, 4.565617e-16, 4.574504e-16, 4.571001e-16, 
    4.579336e-16, 4.584628e-16, 4.582012e-16, 4.598155e-16, 4.591881e-16, 
    4.62489e-16, 4.610684e-16, 4.647693e-16, 4.638847e-16, 4.649812e-16, 
    4.644219e-16, 4.6538e-16, 4.645177e-16, 4.660112e-16, 4.663359e-16, 
    4.66114e-16, 4.669669e-16, 4.644699e-16, 4.654293e-16, 4.581938e-16, 
    4.582365e-16, 4.584354e-16, 4.575607e-16, 4.575073e-16, 4.567056e-16, 
    4.574191e-16, 4.577227e-16, 4.584936e-16, 4.589491e-16, 4.593821e-16, 
    4.603334e-16, 4.613948e-16, 4.628778e-16, 4.639421e-16, 4.64655e-16, 
    4.64218e-16, 4.646038e-16, 4.641724e-16, 4.639702e-16, 4.662142e-16, 
    4.649546e-16, 4.668442e-16, 4.667398e-16, 4.658848e-16, 4.667516e-16, 
    4.582664e-16, 4.580209e-16, 4.571674e-16, 4.578354e-16, 4.566183e-16, 
    4.572995e-16, 4.576909e-16, 4.592009e-16, 4.595328e-16, 4.598399e-16, 
    4.604468e-16, 4.612249e-16, 4.625885e-16, 4.637737e-16, 4.648551e-16, 
    4.647759e-16, 4.648038e-16, 4.650451e-16, 4.644471e-16, 4.651432e-16, 
    4.652598e-16, 4.649546e-16, 4.667258e-16, 4.662201e-16, 4.667376e-16, 
    4.664084e-16, 4.581007e-16, 4.58514e-16, 4.582907e-16, 4.587105e-16, 
    4.584146e-16, 4.597291e-16, 4.60123e-16, 4.619646e-16, 4.612095e-16, 
    4.624114e-16, 4.613317e-16, 4.615231e-16, 4.624499e-16, 4.613902e-16, 
    4.637084e-16, 4.621367e-16, 4.650544e-16, 4.634864e-16, 4.651526e-16, 
    4.648504e-16, 4.653508e-16, 4.657987e-16, 4.663622e-16, 4.674008e-16, 
    4.671604e-16, 4.680286e-16, 4.591299e-16, 4.596653e-16, 4.596184e-16, 
    4.601787e-16, 4.605927e-16, 4.614901e-16, 4.629276e-16, 4.623873e-16, 
    4.633793e-16, 4.635783e-16, 4.620713e-16, 4.629965e-16, 4.600236e-16, 
    4.605042e-16, 4.602183e-16, 4.59172e-16, 4.625115e-16, 4.607987e-16, 
    4.639596e-16, 4.630335e-16, 4.657349e-16, 4.643917e-16, 4.67028e-16, 
    4.681524e-16, 4.692109e-16, 4.704452e-16, 4.599577e-16, 4.595939e-16, 
    4.602454e-16, 4.611454e-16, 4.619808e-16, 4.6309e-16, 4.632035e-16, 
    4.634111e-16, 4.639487e-16, 4.644006e-16, 4.634765e-16, 4.645138e-16, 
    4.606151e-16, 4.626602e-16, 4.594562e-16, 4.604215e-16, 4.610925e-16, 
    4.607985e-16, 4.623257e-16, 4.626852e-16, 4.641448e-16, 4.633908e-16, 
    4.678748e-16, 4.658929e-16, 4.71385e-16, 4.698527e-16, 4.594668e-16, 
    4.599565e-16, 4.61659e-16, 4.608493e-16, 4.631641e-16, 4.637331e-16, 
    4.641953e-16, 4.647859e-16, 4.648499e-16, 4.651997e-16, 4.646264e-16, 
    4.651771e-16, 4.630923e-16, 4.640243e-16, 4.614649e-16, 4.620882e-16, 
    4.618016e-16, 4.614869e-16, 4.624578e-16, 4.634909e-16, 4.635134e-16, 
    4.638442e-16, 4.647756e-16, 4.631734e-16, 4.681295e-16, 4.650703e-16, 
    4.604903e-16, 4.614321e-16, 4.61567e-16, 4.612022e-16, 4.63676e-16, 
    4.627802e-16, 4.651912e-16, 4.645401e-16, 4.656068e-16, 4.650768e-16, 
    4.649988e-16, 4.643178e-16, 4.638935e-16, 4.628212e-16, 4.619479e-16, 
    4.612552e-16, 4.614163e-16, 4.621772e-16, 4.635542e-16, 4.648554e-16, 
    4.645704e-16, 4.655258e-16, 4.629964e-16, 4.640573e-16, 4.636474e-16, 
    4.647164e-16, 4.623729e-16, 4.643674e-16, 4.618623e-16, 4.620823e-16, 
    4.627624e-16, 4.64129e-16, 4.644318e-16, 4.647542e-16, 4.645554e-16, 
    4.635892e-16, 4.63431e-16, 4.62746e-16, 4.625566e-16, 4.620344e-16, 
    4.616017e-16, 4.61997e-16, 4.624118e-16, 4.635898e-16, 4.646499e-16, 
    4.658051e-16, 4.660877e-16, 4.674345e-16, 4.663376e-16, 4.681464e-16, 
    4.666079e-16, 4.692703e-16, 4.644836e-16, 4.665635e-16, 4.627935e-16, 
    4.632004e-16, 4.639352e-16, 4.656204e-16, 4.647114e-16, 4.657746e-16, 
    4.634249e-16, 4.622032e-16, 4.618874e-16, 4.612973e-16, 4.619009e-16, 
    4.618519e-16, 4.624293e-16, 4.622438e-16, 4.636289e-16, 4.628851e-16, 
    4.649967e-16, 4.657663e-16, 4.679375e-16, 4.692662e-16, 4.706178e-16, 
    4.712137e-16, 4.713951e-16, 4.714708e-16 ;

 CWDC_TO_LITR3C =
  1.442543e-16, 1.446451e-16, 1.445692e-16, 1.448841e-16, 1.447095e-16, 
    1.449156e-16, 1.443336e-16, 1.446605e-16, 1.444519e-16, 1.442896e-16, 
    1.454943e-16, 1.448981e-16, 1.461131e-16, 1.457336e-16, 1.466864e-16, 
    1.46054e-16, 1.468138e-16, 1.466683e-16, 1.471064e-16, 1.46981e-16, 
    1.475405e-16, 1.471643e-16, 1.478305e-16, 1.474508e-16, 1.475102e-16, 
    1.471519e-16, 1.450183e-16, 1.454201e-16, 1.449945e-16, 1.450518e-16, 
    1.450261e-16, 1.44713e-16, 1.445551e-16, 1.442245e-16, 1.442846e-16, 
    1.445274e-16, 1.450776e-16, 1.44891e-16, 1.453613e-16, 1.453507e-16, 
    1.458736e-16, 1.456379e-16, 1.465156e-16, 1.462664e-16, 1.469862e-16, 
    1.468053e-16, 1.469777e-16, 1.469255e-16, 1.469784e-16, 1.46713e-16, 
    1.468267e-16, 1.465932e-16, 1.45682e-16, 1.4595e-16, 1.451501e-16, 
    1.446681e-16, 1.443479e-16, 1.441205e-16, 1.441526e-16, 1.442139e-16, 
    1.445288e-16, 1.448248e-16, 1.450501e-16, 1.452008e-16, 1.453492e-16, 
    1.457977e-16, 1.460351e-16, 1.465659e-16, 1.464703e-16, 1.466324e-16, 
    1.467873e-16, 1.470472e-16, 1.470044e-16, 1.471188e-16, 1.466282e-16, 
    1.469543e-16, 1.464158e-16, 1.465631e-16, 1.453891e-16, 1.449414e-16, 
    1.447505e-16, 1.445837e-16, 1.441774e-16, 1.44458e-16, 1.443474e-16, 
    1.446106e-16, 1.447777e-16, 1.446951e-16, 1.452049e-16, 1.450068e-16, 
    1.460492e-16, 1.456005e-16, 1.467692e-16, 1.464899e-16, 1.468362e-16, 
    1.466595e-16, 1.469621e-16, 1.466898e-16, 1.471614e-16, 1.47264e-16, 
    1.471939e-16, 1.474632e-16, 1.466747e-16, 1.469777e-16, 1.446928e-16, 
    1.447062e-16, 1.447691e-16, 1.444929e-16, 1.44476e-16, 1.442228e-16, 
    1.444481e-16, 1.44544e-16, 1.447875e-16, 1.449313e-16, 1.45068e-16, 
    1.453685e-16, 1.457036e-16, 1.461719e-16, 1.46508e-16, 1.467332e-16, 
    1.465951e-16, 1.46717e-16, 1.465808e-16, 1.465169e-16, 1.472255e-16, 
    1.468278e-16, 1.474245e-16, 1.473915e-16, 1.471215e-16, 1.473952e-16, 
    1.447157e-16, 1.446382e-16, 1.443687e-16, 1.445796e-16, 1.441952e-16, 
    1.444104e-16, 1.44534e-16, 1.450108e-16, 1.451156e-16, 1.452126e-16, 
    1.454042e-16, 1.4565e-16, 1.460806e-16, 1.464549e-16, 1.467963e-16, 
    1.467713e-16, 1.467801e-16, 1.468563e-16, 1.466675e-16, 1.468873e-16, 
    1.469242e-16, 1.468278e-16, 1.473871e-16, 1.472274e-16, 1.473908e-16, 
    1.472869e-16, 1.446634e-16, 1.447939e-16, 1.447234e-16, 1.448559e-16, 
    1.447625e-16, 1.451776e-16, 1.45302e-16, 1.458835e-16, 1.456451e-16, 
    1.460246e-16, 1.456837e-16, 1.457441e-16, 1.460368e-16, 1.457022e-16, 
    1.464342e-16, 1.459379e-16, 1.468593e-16, 1.463641e-16, 1.468903e-16, 
    1.467949e-16, 1.469529e-16, 1.470943e-16, 1.472723e-16, 1.476002e-16, 
    1.475243e-16, 1.477985e-16, 1.449884e-16, 1.451575e-16, 1.451427e-16, 
    1.453196e-16, 1.454503e-16, 1.457337e-16, 1.461877e-16, 1.460171e-16, 
    1.463303e-16, 1.463931e-16, 1.459173e-16, 1.462094e-16, 1.452706e-16, 
    1.454224e-16, 1.453321e-16, 1.450017e-16, 1.460563e-16, 1.455154e-16, 
    1.465136e-16, 1.462211e-16, 1.470742e-16, 1.4665e-16, 1.474825e-16, 
    1.478376e-16, 1.481719e-16, 1.485616e-16, 1.452498e-16, 1.451349e-16, 
    1.453406e-16, 1.456249e-16, 1.458887e-16, 1.462389e-16, 1.462748e-16, 
    1.463403e-16, 1.465101e-16, 1.466528e-16, 1.46361e-16, 1.466886e-16, 
    1.454574e-16, 1.461032e-16, 1.450914e-16, 1.453963e-16, 1.456082e-16, 
    1.455153e-16, 1.459976e-16, 1.461111e-16, 1.46572e-16, 1.463339e-16, 
    1.477499e-16, 1.471241e-16, 1.488584e-16, 1.483745e-16, 1.450948e-16, 
    1.452494e-16, 1.45787e-16, 1.455314e-16, 1.462623e-16, 1.46442e-16, 
    1.46588e-16, 1.467745e-16, 1.467947e-16, 1.469051e-16, 1.467241e-16, 
    1.46898e-16, 1.462397e-16, 1.46534e-16, 1.457257e-16, 1.459226e-16, 
    1.458321e-16, 1.457327e-16, 1.460393e-16, 1.463656e-16, 1.463727e-16, 
    1.464771e-16, 1.467712e-16, 1.462653e-16, 1.478304e-16, 1.468643e-16, 
    1.45418e-16, 1.457154e-16, 1.45758e-16, 1.456428e-16, 1.46424e-16, 
    1.461411e-16, 1.469025e-16, 1.466969e-16, 1.470337e-16, 1.468664e-16, 
    1.468417e-16, 1.466267e-16, 1.464927e-16, 1.461541e-16, 1.458783e-16, 
    1.456595e-16, 1.457104e-16, 1.459507e-16, 1.463855e-16, 1.467965e-16, 
    1.467065e-16, 1.470081e-16, 1.462094e-16, 1.465444e-16, 1.46415e-16, 
    1.467525e-16, 1.460125e-16, 1.466424e-16, 1.458513e-16, 1.459207e-16, 
    1.461355e-16, 1.46567e-16, 1.466627e-16, 1.467645e-16, 1.467017e-16, 
    1.463966e-16, 1.463466e-16, 1.461303e-16, 1.460705e-16, 1.459056e-16, 
    1.45769e-16, 1.458938e-16, 1.460248e-16, 1.463968e-16, 1.467315e-16, 
    1.470963e-16, 1.471856e-16, 1.476109e-16, 1.472645e-16, 1.478357e-16, 
    1.473499e-16, 1.481906e-16, 1.46679e-16, 1.473358e-16, 1.461453e-16, 
    1.462738e-16, 1.465059e-16, 1.47038e-16, 1.46751e-16, 1.470867e-16, 
    1.463447e-16, 1.459589e-16, 1.458592e-16, 1.456728e-16, 1.458635e-16, 
    1.45848e-16, 1.460303e-16, 1.459717e-16, 1.464091e-16, 1.461742e-16, 
    1.468411e-16, 1.470841e-16, 1.477697e-16, 1.481893e-16, 1.486161e-16, 
    1.488043e-16, 1.488616e-16, 1.488855e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  9.136104e-19, 9.160856e-19, 9.156048e-19, 9.175992e-19, 9.164934e-19, 
    9.177988e-19, 9.141128e-19, 9.161834e-19, 9.14862e-19, 9.138339e-19, 
    9.21464e-19, 9.176882e-19, 9.253832e-19, 9.229793e-19, 9.290139e-19, 
    9.250087e-19, 9.298209e-19, 9.288993e-19, 9.316742e-19, 9.308796e-19, 
    9.344234e-19, 9.320409e-19, 9.362597e-19, 9.338551e-19, 9.342311e-19, 
    9.319621e-19, 9.184493e-19, 9.20994e-19, 9.182984e-19, 9.186614e-19, 
    9.184987e-19, 9.165159e-19, 9.155155e-19, 9.134217e-19, 9.138021e-19, 
    9.153403e-19, 9.188247e-19, 9.17643e-19, 9.206217e-19, 9.205545e-19, 
    9.238658e-19, 9.223734e-19, 9.279321e-19, 9.263541e-19, 9.309128e-19, 
    9.297669e-19, 9.308589e-19, 9.305279e-19, 9.308632e-19, 9.291824e-19, 
    9.299027e-19, 9.284234e-19, 9.226528e-19, 9.243501e-19, 9.192839e-19, 
    9.162312e-19, 9.142035e-19, 9.127631e-19, 9.129668e-19, 9.133548e-19, 
    9.153493e-19, 9.172237e-19, 9.186509e-19, 9.19605e-19, 9.205448e-19, 
    9.233851e-19, 9.248889e-19, 9.282507e-19, 9.27645e-19, 9.286716e-19, 
    9.29653e-19, 9.312987e-19, 9.31028e-19, 9.317525e-19, 9.286451e-19, 
    9.307104e-19, 9.273003e-19, 9.28233e-19, 9.207974e-19, 9.17962e-19, 
    9.167533e-19, 9.156971e-19, 9.131233e-19, 9.149008e-19, 9.142002e-19, 
    9.158673e-19, 9.169257e-19, 9.164024e-19, 9.196311e-19, 9.183762e-19, 
    9.249781e-19, 9.221367e-19, 9.295385e-19, 9.277694e-19, 9.299625e-19, 
    9.288438e-19, 9.3076e-19, 9.290355e-19, 9.320223e-19, 9.326719e-19, 
    9.32228e-19, 9.339338e-19, 9.289398e-19, 9.308586e-19, 9.163876e-19, 
    9.164729e-19, 9.168708e-19, 9.151215e-19, 9.150146e-19, 9.134112e-19, 
    9.148382e-19, 9.154453e-19, 9.169872e-19, 9.178982e-19, 9.187641e-19, 
    9.206669e-19, 9.227897e-19, 9.257556e-19, 9.278841e-19, 9.2931e-19, 
    9.28436e-19, 9.292077e-19, 9.283449e-19, 9.279405e-19, 9.324284e-19, 
    9.299092e-19, 9.336885e-19, 9.334796e-19, 9.317696e-19, 9.335032e-19, 
    9.165329e-19, 9.160417e-19, 9.143347e-19, 9.156707e-19, 9.132366e-19, 
    9.14599e-19, 9.153818e-19, 9.184019e-19, 9.190656e-19, 9.1968e-19, 
    9.208936e-19, 9.224498e-19, 9.251771e-19, 9.275475e-19, 9.297102e-19, 
    9.295519e-19, 9.296075e-19, 9.300902e-19, 9.288942e-19, 9.302864e-19, 
    9.305197e-19, 9.299092e-19, 9.334516e-19, 9.324402e-19, 9.334752e-19, 
    9.328167e-19, 9.162015e-19, 9.170279e-19, 9.165814e-19, 9.17421e-19, 
    9.168292e-19, 9.194583e-19, 9.20246e-19, 9.239291e-19, 9.22419e-19, 
    9.248228e-19, 9.226635e-19, 9.230461e-19, 9.248999e-19, 9.227805e-19, 
    9.274168e-19, 9.242734e-19, 9.301089e-19, 9.269728e-19, 9.303052e-19, 
    9.297008e-19, 9.307017e-19, 9.315975e-19, 9.327244e-19, 9.348016e-19, 
    9.343209e-19, 9.360572e-19, 9.182598e-19, 9.193306e-19, 9.192368e-19, 
    9.203573e-19, 9.211856e-19, 9.229802e-19, 9.258553e-19, 9.247747e-19, 
    9.267587e-19, 9.271566e-19, 9.241426e-19, 9.25993e-19, 9.200472e-19, 
    9.210084e-19, 9.204366e-19, 9.18344e-19, 9.250231e-19, 9.215974e-19, 
    9.279192e-19, 9.26067e-19, 9.314697e-19, 9.287835e-19, 9.340561e-19, 
    9.363049e-19, 9.384219e-19, 9.408903e-19, 9.199153e-19, 9.191879e-19, 
    9.204906e-19, 9.222909e-19, 9.239615e-19, 9.261799e-19, 9.26407e-19, 
    9.268222e-19, 9.278973e-19, 9.288011e-19, 9.269529e-19, 9.290276e-19, 
    9.212301e-19, 9.253204e-19, 9.189124e-19, 9.208431e-19, 9.221851e-19, 
    9.215971e-19, 9.246513e-19, 9.253704e-19, 9.282896e-19, 9.267815e-19, 
    9.357495e-19, 9.317859e-19, 9.427699e-19, 9.397054e-19, 9.189336e-19, 
    9.19913e-19, 9.23318e-19, 9.216986e-19, 9.263281e-19, 9.274661e-19, 
    9.283907e-19, 9.295718e-19, 9.296997e-19, 9.303993e-19, 9.292527e-19, 
    9.303542e-19, 9.261846e-19, 9.280487e-19, 9.229297e-19, 9.241764e-19, 
    9.236032e-19, 9.229738e-19, 9.249156e-19, 9.269819e-19, 9.270269e-19, 
    9.276883e-19, 9.295511e-19, 9.26347e-19, 9.36259e-19, 9.301407e-19, 
    9.209806e-19, 9.22864e-19, 9.23134e-19, 9.224045e-19, 9.27352e-19, 
    9.255604e-19, 9.303824e-19, 9.290802e-19, 9.312137e-19, 9.301536e-19, 
    9.299976e-19, 9.286357e-19, 9.277871e-19, 9.256424e-19, 9.238958e-19, 
    9.225104e-19, 9.228327e-19, 9.243544e-19, 9.271084e-19, 9.297109e-19, 
    9.291409e-19, 9.310515e-19, 9.259927e-19, 9.281146e-19, 9.272948e-19, 
    9.294329e-19, 9.247457e-19, 9.287349e-19, 9.237246e-19, 9.241645e-19, 
    9.255248e-19, 9.282578e-19, 9.288635e-19, 9.295084e-19, 9.291107e-19, 
    9.271785e-19, 9.268621e-19, 9.25492e-19, 9.251132e-19, 9.240688e-19, 
    9.232035e-19, 9.239939e-19, 9.248236e-19, 9.271796e-19, 9.292998e-19, 
    9.316101e-19, 9.321755e-19, 9.34869e-19, 9.326753e-19, 9.362929e-19, 
    9.332158e-19, 9.385406e-19, 9.289672e-19, 9.33127e-19, 9.25587e-19, 
    9.264008e-19, 9.278704e-19, 9.312409e-19, 9.294228e-19, 9.315492e-19, 
    9.268497e-19, 9.244064e-19, 9.237749e-19, 9.225946e-19, 9.238019e-19, 
    9.237038e-19, 9.248585e-19, 9.244876e-19, 9.272578e-19, 9.257702e-19, 
    9.299935e-19, 9.315327e-19, 9.35875e-19, 9.385324e-19, 9.412355e-19, 
    9.424273e-19, 9.427901e-19, 9.429416e-19 ;

 CWDN_TO_LITR3N =
  2.885086e-19, 2.892902e-19, 2.891383e-19, 2.897682e-19, 2.89419e-19, 
    2.898312e-19, 2.886672e-19, 2.893211e-19, 2.889038e-19, 2.885791e-19, 
    2.909886e-19, 2.897963e-19, 2.922263e-19, 2.914671e-19, 2.933728e-19, 
    2.92108e-19, 2.936277e-19, 2.933366e-19, 2.942129e-19, 2.93962e-19, 
    2.950811e-19, 2.943287e-19, 2.956609e-19, 2.949016e-19, 2.950204e-19, 
    2.943038e-19, 2.900366e-19, 2.908402e-19, 2.899889e-19, 2.901036e-19, 
    2.900522e-19, 2.894261e-19, 2.891102e-19, 2.88449e-19, 2.885691e-19, 
    2.890548e-19, 2.901552e-19, 2.89782e-19, 2.907227e-19, 2.907014e-19, 
    2.917471e-19, 2.912758e-19, 2.930312e-19, 2.925329e-19, 2.939725e-19, 
    2.936106e-19, 2.939554e-19, 2.938509e-19, 2.939568e-19, 2.93426e-19, 
    2.936535e-19, 2.931863e-19, 2.913641e-19, 2.919e-19, 2.903002e-19, 
    2.893361e-19, 2.886959e-19, 2.88241e-19, 2.883053e-19, 2.884279e-19, 
    2.890576e-19, 2.896496e-19, 2.901003e-19, 2.904016e-19, 2.906984e-19, 
    2.915953e-19, 2.920702e-19, 2.931318e-19, 2.929405e-19, 2.932647e-19, 
    2.935746e-19, 2.940943e-19, 2.940088e-19, 2.942376e-19, 2.932563e-19, 
    2.939086e-19, 2.928317e-19, 2.931262e-19, 2.907781e-19, 2.898827e-19, 
    2.895011e-19, 2.891675e-19, 2.883547e-19, 2.889161e-19, 2.886948e-19, 
    2.892213e-19, 2.895555e-19, 2.893902e-19, 2.904098e-19, 2.900136e-19, 
    2.920983e-19, 2.912011e-19, 2.935385e-19, 2.929798e-19, 2.936724e-19, 
    2.933191e-19, 2.939242e-19, 2.933796e-19, 2.943229e-19, 2.94528e-19, 
    2.943878e-19, 2.949264e-19, 2.933494e-19, 2.939553e-19, 2.893855e-19, 
    2.894125e-19, 2.895381e-19, 2.889857e-19, 2.88952e-19, 2.884456e-19, 
    2.888963e-19, 2.89088e-19, 2.895749e-19, 2.898626e-19, 2.90136e-19, 
    2.907369e-19, 2.914073e-19, 2.923439e-19, 2.93016e-19, 2.934663e-19, 
    2.931903e-19, 2.93434e-19, 2.931615e-19, 2.930339e-19, 2.944511e-19, 
    2.936555e-19, 2.94849e-19, 2.94783e-19, 2.94243e-19, 2.947905e-19, 
    2.894315e-19, 2.892763e-19, 2.887373e-19, 2.891592e-19, 2.883905e-19, 
    2.888207e-19, 2.89068e-19, 2.900216e-19, 2.902312e-19, 2.904252e-19, 
    2.908085e-19, 2.912999e-19, 2.921612e-19, 2.929097e-19, 2.935927e-19, 
    2.935427e-19, 2.935603e-19, 2.937127e-19, 2.93335e-19, 2.937747e-19, 
    2.938483e-19, 2.936556e-19, 2.947742e-19, 2.944548e-19, 2.947816e-19, 
    2.945737e-19, 2.893268e-19, 2.895878e-19, 2.894467e-19, 2.897119e-19, 
    2.89525e-19, 2.903553e-19, 2.90604e-19, 2.917671e-19, 2.912902e-19, 
    2.920493e-19, 2.913674e-19, 2.914882e-19, 2.920736e-19, 2.914044e-19, 
    2.928685e-19, 2.918758e-19, 2.937186e-19, 2.927283e-19, 2.937806e-19, 
    2.935897e-19, 2.939058e-19, 2.941887e-19, 2.945446e-19, 2.952005e-19, 
    2.950487e-19, 2.95597e-19, 2.899768e-19, 2.903149e-19, 2.902853e-19, 
    2.906392e-19, 2.909007e-19, 2.914674e-19, 2.923753e-19, 2.920341e-19, 
    2.926606e-19, 2.927863e-19, 2.918345e-19, 2.924189e-19, 2.905412e-19, 
    2.908448e-19, 2.906642e-19, 2.900033e-19, 2.921125e-19, 2.910307e-19, 
    2.930271e-19, 2.924422e-19, 2.941483e-19, 2.933001e-19, 2.949651e-19, 
    2.956752e-19, 2.963438e-19, 2.971233e-19, 2.904996e-19, 2.902699e-19, 
    2.906813e-19, 2.912498e-19, 2.917773e-19, 2.924779e-19, 2.925496e-19, 
    2.926807e-19, 2.930202e-19, 2.933056e-19, 2.92722e-19, 2.933772e-19, 
    2.909148e-19, 2.922064e-19, 2.901828e-19, 2.907926e-19, 2.912163e-19, 
    2.910307e-19, 2.919951e-19, 2.922222e-19, 2.931441e-19, 2.926678e-19, 
    2.954999e-19, 2.942482e-19, 2.977168e-19, 2.967491e-19, 2.901896e-19, 
    2.904989e-19, 2.915741e-19, 2.910627e-19, 2.925247e-19, 2.92884e-19, 
    2.93176e-19, 2.93549e-19, 2.935894e-19, 2.938103e-19, 2.934482e-19, 
    2.937961e-19, 2.924794e-19, 2.93068e-19, 2.914515e-19, 2.918452e-19, 
    2.916642e-19, 2.914654e-19, 2.920786e-19, 2.927311e-19, 2.927453e-19, 
    2.929542e-19, 2.935425e-19, 2.925306e-19, 2.956607e-19, 2.937286e-19, 
    2.90836e-19, 2.914307e-19, 2.91516e-19, 2.912856e-19, 2.92848e-19, 
    2.922822e-19, 2.93805e-19, 2.933938e-19, 2.940675e-19, 2.937327e-19, 
    2.936835e-19, 2.932534e-19, 2.929854e-19, 2.923081e-19, 2.917566e-19, 
    2.913191e-19, 2.914208e-19, 2.919014e-19, 2.927711e-19, 2.935929e-19, 
    2.934129e-19, 2.940163e-19, 2.924188e-19, 2.930888e-19, 2.928299e-19, 
    2.935051e-19, 2.92025e-19, 2.932847e-19, 2.917025e-19, 2.918414e-19, 
    2.92271e-19, 2.931341e-19, 2.933253e-19, 2.93529e-19, 2.934034e-19, 
    2.927932e-19, 2.926933e-19, 2.922606e-19, 2.92141e-19, 2.918112e-19, 
    2.915379e-19, 2.917875e-19, 2.920495e-19, 2.927936e-19, 2.934631e-19, 
    2.941927e-19, 2.943712e-19, 2.952218e-19, 2.945291e-19, 2.956714e-19, 
    2.946997e-19, 2.963812e-19, 2.933581e-19, 2.946717e-19, 2.922906e-19, 
    2.925476e-19, 2.930117e-19, 2.94076e-19, 2.935019e-19, 2.941734e-19, 
    2.926894e-19, 2.919178e-19, 2.917184e-19, 2.913456e-19, 2.917269e-19, 
    2.916959e-19, 2.920606e-19, 2.919434e-19, 2.928183e-19, 2.923485e-19, 
    2.936822e-19, 2.941682e-19, 2.955395e-19, 2.963786e-19, 2.972323e-19, 
    2.976087e-19, 2.977232e-19, 2.977711e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.809094e-14, 2.821619e-14, 2.819177e-14, 2.829288e-14, 2.823673e-14, 
    2.830293e-14, 2.811618e-14, 2.822102e-14, 2.815403e-14, 2.810197e-14, 
    2.848916e-14, 2.82972e-14, 2.868852e-14, 2.856592e-14, 2.887386e-14, 
    2.866942e-14, 2.891508e-14, 2.886783e-14, 2.900978e-14, 2.896906e-14, 
    2.915084e-14, 2.902849e-14, 2.9245e-14, 2.912153e-14, 2.914084e-14, 
    2.902435e-14, 2.833592e-14, 2.846545e-14, 2.832822e-14, 2.834668e-14, 
    2.833835e-14, 2.823781e-14, 2.818722e-14, 2.808111e-14, 2.810031e-14, 
    2.817821e-14, 2.83548e-14, 2.829475e-14, 2.84459e-14, 2.844249e-14, 
    2.861096e-14, 2.853496e-14, 2.881838e-14, 2.873772e-14, 2.897073e-14, 
    2.891207e-14, 2.896793e-14, 2.895094e-14, 2.896808e-14, 2.888212e-14, 
    2.89189e-14, 2.884325e-14, 2.85495e-14, 2.863592e-14, 2.837821e-14, 
    2.822351e-14, 2.812068e-14, 2.804783e-14, 2.805808e-14, 2.807773e-14, 
    2.817861e-14, 2.827347e-14, 2.834583e-14, 2.839423e-14, 2.844193e-14, 
    2.858666e-14, 2.866315e-14, 2.883466e-14, 2.880362e-14, 2.885611e-14, 
    2.890621e-14, 2.89904e-14, 2.897652e-14, 2.901361e-14, 2.885455e-14, 
    2.896025e-14, 2.878575e-14, 2.883346e-14, 2.845536e-14, 2.831104e-14, 
    2.824991e-14, 2.819625e-14, 2.806598e-14, 2.815592e-14, 2.812044e-14, 
    2.820472e-14, 2.825834e-14, 2.823177e-14, 2.839553e-14, 2.833181e-14, 
    2.866764e-14, 2.852289e-14, 2.890039e-14, 2.880993e-14, 2.892199e-14, 
    2.886478e-14, 2.896279e-14, 2.887454e-14, 2.902737e-14, 2.90607e-14, 
    2.903787e-14, 2.91253e-14, 2.88695e-14, 2.89677e-14, 2.823118e-14, 
    2.823551e-14, 2.825562e-14, 2.816706e-14, 2.816162e-14, 2.808044e-14, 
    2.815259e-14, 2.818336e-14, 2.826137e-14, 2.830755e-14, 2.835145e-14, 
    2.844809e-14, 2.855609e-14, 2.870716e-14, 2.881577e-14, 2.888858e-14, 
    2.884388e-14, 2.888329e-14, 2.883919e-14, 2.881847e-14, 2.904815e-14, 
    2.891915e-14, 2.911265e-14, 2.910193e-14, 2.901431e-14, 2.910307e-14, 
    2.82385e-14, 2.821356e-14, 2.812718e-14, 2.819473e-14, 2.807156e-14, 
    2.81405e-14, 2.818014e-14, 2.833315e-14, 2.836671e-14, 2.839794e-14, 
    2.845954e-14, 2.853866e-14, 2.867762e-14, 2.879855e-14, 2.890901e-14, 
    2.890087e-14, 2.890372e-14, 2.892838e-14, 2.88672e-14, 2.893838e-14, 
    2.895032e-14, 2.891905e-14, 2.910043e-14, 2.904858e-14, 2.910161e-14, 
    2.90678e-14, 2.822162e-14, 2.826348e-14, 2.824081e-14, 2.82834e-14, 
    2.825336e-14, 2.838679e-14, 2.842679e-14, 2.861412e-14, 2.853712e-14, 
    2.865958e-14, 2.854949e-14, 2.8569e-14, 2.866358e-14, 2.855535e-14, 
    2.879184e-14, 2.863151e-14, 2.892932e-14, 2.876917e-14, 2.893931e-14, 
    2.890833e-14, 2.895951e-14, 2.900541e-14, 2.906308e-14, 2.91697e-14, 
    2.914494e-14, 2.92341e-14, 2.832591e-14, 2.838027e-14, 2.837543e-14, 
    2.843231e-14, 2.84744e-14, 2.856568e-14, 2.871219e-14, 2.865702e-14, 
    2.875817e-14, 2.877851e-14, 2.862471e-14, 2.871913e-14, 2.841641e-14, 
    2.846527e-14, 2.843612e-14, 2.832985e-14, 2.866957e-14, 2.849511e-14, 
    2.881727e-14, 2.872264e-14, 2.89988e-14, 2.886144e-14, 2.913134e-14, 
    2.924696e-14, 2.935561e-14, 2.948288e-14, 2.84099e-14, 2.837289e-14, 
    2.843902e-14, 2.853069e-14, 2.861561e-14, 2.872871e-14, 2.874023e-14, 
    2.87614e-14, 2.881627e-14, 2.886247e-14, 2.876809e-14, 2.887397e-14, 
    2.847667e-14, 2.868469e-14, 2.835863e-14, 2.845679e-14, 2.852492e-14, 
    2.849497e-14, 2.865038e-14, 2.868702e-14, 2.883609e-14, 2.875898e-14, 
    2.921838e-14, 2.901498e-14, 2.957967e-14, 2.942173e-14, 2.835996e-14, 
    2.840965e-14, 2.858286e-14, 2.850041e-14, 2.873617e-14, 2.879429e-14, 
    2.884145e-14, 2.890191e-14, 2.890835e-14, 2.894417e-14, 2.888543e-14, 
    2.894179e-14, 2.872868e-14, 2.882386e-14, 2.856273e-14, 2.862623e-14, 
    2.859697e-14, 2.856489e-14, 2.866378e-14, 2.87693e-14, 2.877146e-14, 
    2.880528e-14, 2.890083e-14, 2.873667e-14, 2.924467e-14, 2.893085e-14, 
    2.846387e-14, 2.855977e-14, 2.857337e-14, 2.853621e-14, 2.878839e-14, 
    2.869697e-14, 2.894329e-14, 2.887662e-14, 2.898575e-14, 2.893151e-14, 
    2.892348e-14, 2.885382e-14, 2.881043e-14, 2.870098e-14, 2.86119e-14, 
    2.85413e-14, 2.855765e-14, 2.863522e-14, 2.877567e-14, 2.890866e-14, 
    2.88795e-14, 2.897714e-14, 2.871855e-14, 2.882697e-14, 2.878503e-14, 
    2.889426e-14, 2.865546e-14, 2.885943e-14, 2.860336e-14, 2.862575e-14, 
    2.869508e-14, 2.883474e-14, 2.88655e-14, 2.889853e-14, 2.887808e-14, 
    2.877941e-14, 2.876319e-14, 2.869322e-14, 2.867391e-14, 2.862064e-14, 
    2.857651e-14, 2.86168e-14, 2.865907e-14, 2.877923e-14, 2.888759e-14, 
    2.900577e-14, 2.903468e-14, 2.917304e-14, 2.906044e-14, 2.924631e-14, 
    2.908837e-14, 2.936173e-14, 2.887109e-14, 2.908411e-14, 2.869823e-14, 
    2.87397e-14, 2.881487e-14, 2.898724e-14, 2.889404e-14, 2.900298e-14, 
    2.876254e-14, 2.863797e-14, 2.860565e-14, 2.854557e-14, 2.860698e-14, 
    2.860198e-14, 2.866078e-14, 2.864183e-14, 2.878315e-14, 2.870721e-14, 
    2.892297e-14, 2.900181e-14, 2.922449e-14, 2.936115e-14, 2.950027e-14, 
    2.956171e-14, 2.958041e-14, 2.958821e-14 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  5.938781, 5.957684, 5.954026, 5.969241, 5.960828, 5.970763, 5.942647, 
    5.958405, 5.948364, 5.940529, 5.998516, 5.969925, 6.028523, 6.010238, 
    6.058059, 6.025631, 6.064271, 6.057249, 6.078579, 6.072471, 6.09962, 
    6.0814, 6.113836, 6.095308, 6.098176, 6.080787, 5.975749, 5.99493, 
    5.974595, 5.977334, 5.976122, 5.960975, 5.953274, 5.93739, 5.940287, 
    5.951983, 5.978567, 5.969627, 5.992313, 5.991802, 6.017004, 6.005643, 
    6.049834, 6.036029, 6.072728, 6.063916, 6.0723, 6.069767, 6.072333, 
    6.059416, 6.064945, 6.053609, 6.007757, 6.020682, 5.982082, 5.9587, 
    5.943325, 5.932361, 5.93391, 5.936848, 5.95205, 5.96642, 5.977303, 
    5.984561, 5.991727, 6.01321, 6.024749, 6.052238, 6.04765, 6.055472, 
    6.063043, 6.075673, 6.073603, 6.079154, 6.055313, 6.071131, 6.043277, 
    6.052151, 5.993418, 5.97205, 5.962708, 5.95472, 5.935096, 5.948632, 
    5.943289, 5.956058, 5.964138, 5.960152, 5.984761, 5.975203, 6.025434, 
    6.003803, 6.06216, 6.048597, 6.065423, 6.056846, 6.071522, 6.058314, 
    6.081241, 6.086207, 6.082808, 6.095959, 6.057575, 6.072275, 5.960028, 
    5.960676, 5.963728, 5.950311, 5.949506, 5.937298, 5.948184, 5.9528, 
    5.964627, 5.971562, 5.978146, 5.992634, 6.008766, 6.031404, 6.049473, 
    6.060422, 6.053724, 6.059635, 6.053018, 6.049929, 6.08433, 6.064981, 
    6.094066, 6.092464, 6.079276, 6.092646, 5.961136, 5.957397, 5.944334, 
    5.954556, 5.935972, 5.94634, 5.952283, 5.975346, 5.980454, 5.985112, 
    5.994374, 6.006223, 6.026993, 6.046871, 6.063494, 6.062281, 6.062706, 
    6.066395, 6.057221, 6.067904, 6.069672, 6.06501, 6.092248, 6.084466, 
    6.09243, 6.087368, 5.958619, 5.964924, 5.961512, 5.967914, 5.963383, 
    5.983372, 5.989357, 6.017428, 6.005975, 6.024277, 6.007854, 6.010748, 
    6.024766, 6.008758, 6.044075, 6.020026, 6.066539, 6.040624, 6.068048, 
    6.063422, 6.071109, 6.077968, 6.086648, 6.102602, 6.098917, 6.11231, 
    5.974319, 5.982429, 5.981762, 5.990287, 5.996583, 6.010276, 6.032193, 
    6.023963, 6.039126, 6.042155, 6.019148, 6.033225, 5.987895, 5.995171, 
    5.990874, 5.97493, 6.025793, 5.999666, 6.049735, 6.033821, 6.076983, 
    6.056315, 6.096877, 6.11412, 6.130592, 6.149598, 5.986909, 5.981391, 
    5.991315, 6.004954, 6.017739, 6.034676, 6.036436, 6.039596, 6.049595, 
    6.056516, 6.040548, 6.058257, 5.996761, 6.028086, 5.979261, 5.993901, 
    6.004172, 5.999718, 6.023036, 6.028518, 6.052548, 6.039303, 6.109819, 
    6.079348, 6.164248, 6.140445, 5.979452, 5.986913, 6.012804, 6.000499, 
    6.035832, 6.044518, 6.053378, 6.062396, 6.063406, 6.068759, 6.059982, 
    6.068431, 6.034711, 6.05074, 6.009903, 6.01938, 6.015036, 6.010237, 
    6.025048, 6.04076, 6.041173, 6.047949, 6.062, 6.035976, 6.113611, 
    6.066559, 5.995046, 6.009305, 6.011436, 6.005898, 6.043644, 6.029949, 
    6.06864, 6.058658, 6.075037, 6.066889, 6.065687, 6.055248, 6.048732, 
    6.030561, 6.017232, 6.006711, 6.009162, 6.020725, 6.041739, 6.063463, 
    6.059072, 6.073792, 6.033265, 6.051214, 6.043174, 6.061351, 6.023727, 
    6.05578, 6.015963, 6.019313, 6.029678, 6.052262, 6.056994, 6.06191, 
    6.058893, 6.042287, 6.039891, 6.029445, 6.026523, 6.01859, 6.011989, 
    6.018001, 6.0243, 6.042326, 6.060304, 6.078053, 6.08243, 6.103, 6.086145, 
    6.113858, 6.09013, 6.131308, 6.057653, 6.089593, 6.030176, 6.036392, 
    6.049309, 6.075148, 6.061275, 6.077538, 6.039804, 6.021085, 6.016341, 
    6.007336, 6.016547, 6.015801, 6.024616, 6.021788, 6.042926, 6.031572, 
    6.065636, 6.077429, 6.110877, 6.131366, 6.152376, 6.161618, 6.164439, 
    6.165614 ;

 EFLX_LH_TOT_R =
  5.938781, 5.957684, 5.954026, 5.969241, 5.960828, 5.970763, 5.942647, 
    5.958405, 5.948364, 5.940529, 5.998516, 5.969925, 6.028523, 6.010238, 
    6.058059, 6.025631, 6.064271, 6.057249, 6.078579, 6.072471, 6.09962, 
    6.0814, 6.113836, 6.095308, 6.098176, 6.080787, 5.975749, 5.99493, 
    5.974595, 5.977334, 5.976122, 5.960975, 5.953274, 5.93739, 5.940287, 
    5.951983, 5.978567, 5.969627, 5.992313, 5.991802, 6.017004, 6.005643, 
    6.049834, 6.036029, 6.072728, 6.063916, 6.0723, 6.069767, 6.072333, 
    6.059416, 6.064945, 6.053609, 6.007757, 6.020682, 5.982082, 5.9587, 
    5.943325, 5.932361, 5.93391, 5.936848, 5.95205, 5.96642, 5.977303, 
    5.984561, 5.991727, 6.01321, 6.024749, 6.052238, 6.04765, 6.055472, 
    6.063043, 6.075673, 6.073603, 6.079154, 6.055313, 6.071131, 6.043277, 
    6.052151, 5.993418, 5.97205, 5.962708, 5.95472, 5.935096, 5.948632, 
    5.943289, 5.956058, 5.964138, 5.960152, 5.984761, 5.975203, 6.025434, 
    6.003803, 6.06216, 6.048597, 6.065423, 6.056846, 6.071522, 6.058314, 
    6.081241, 6.086207, 6.082808, 6.095959, 6.057575, 6.072275, 5.960028, 
    5.960676, 5.963728, 5.950311, 5.949506, 5.937298, 5.948184, 5.9528, 
    5.964627, 5.971562, 5.978146, 5.992634, 6.008766, 6.031404, 6.049473, 
    6.060422, 6.053724, 6.059635, 6.053018, 6.049929, 6.08433, 6.064981, 
    6.094066, 6.092464, 6.079276, 6.092646, 5.961136, 5.957397, 5.944334, 
    5.954556, 5.935972, 5.94634, 5.952283, 5.975346, 5.980454, 5.985112, 
    5.994374, 6.006223, 6.026993, 6.046871, 6.063494, 6.062281, 6.062706, 
    6.066395, 6.057221, 6.067904, 6.069672, 6.06501, 6.092248, 6.084466, 
    6.09243, 6.087368, 5.958619, 5.964924, 5.961512, 5.967914, 5.963383, 
    5.983372, 5.989357, 6.017428, 6.005975, 6.024277, 6.007854, 6.010748, 
    6.024766, 6.008758, 6.044075, 6.020026, 6.066539, 6.040624, 6.068048, 
    6.063422, 6.071109, 6.077968, 6.086648, 6.102602, 6.098917, 6.11231, 
    5.974319, 5.982429, 5.981762, 5.990287, 5.996583, 6.010276, 6.032193, 
    6.023963, 6.039126, 6.042155, 6.019148, 6.033225, 5.987895, 5.995171, 
    5.990874, 5.97493, 6.025793, 5.999666, 6.049735, 6.033821, 6.076983, 
    6.056315, 6.096877, 6.11412, 6.130592, 6.149598, 5.986909, 5.981391, 
    5.991315, 6.004954, 6.017739, 6.034676, 6.036436, 6.039596, 6.049595, 
    6.056516, 6.040548, 6.058257, 5.996761, 6.028086, 5.979261, 5.993901, 
    6.004172, 5.999718, 6.023036, 6.028518, 6.052548, 6.039303, 6.109819, 
    6.079348, 6.164248, 6.140445, 5.979452, 5.986913, 6.012804, 6.000499, 
    6.035832, 6.044518, 6.053378, 6.062396, 6.063406, 6.068759, 6.059982, 
    6.068431, 6.034711, 6.05074, 6.009903, 6.01938, 6.015036, 6.010237, 
    6.025048, 6.04076, 6.041173, 6.047949, 6.062, 6.035976, 6.113611, 
    6.066559, 5.995046, 6.009305, 6.011436, 6.005898, 6.043644, 6.029949, 
    6.06864, 6.058658, 6.075037, 6.066889, 6.065687, 6.055248, 6.048732, 
    6.030561, 6.017232, 6.006711, 6.009162, 6.020725, 6.041739, 6.063463, 
    6.059072, 6.073792, 6.033265, 6.051214, 6.043174, 6.061351, 6.023727, 
    6.05578, 6.015963, 6.019313, 6.029678, 6.052262, 6.056994, 6.06191, 
    6.058893, 6.042287, 6.039891, 6.029445, 6.026523, 6.01859, 6.011989, 
    6.018001, 6.0243, 6.042326, 6.060304, 6.078053, 6.08243, 6.103, 6.086145, 
    6.113858, 6.09013, 6.131308, 6.057653, 6.089593, 6.030176, 6.036392, 
    6.049309, 6.075148, 6.061275, 6.077538, 6.039804, 6.021085, 6.016341, 
    6.007336, 6.016547, 6.015801, 6.024616, 6.021788, 6.042926, 6.031572, 
    6.065636, 6.077429, 6.110877, 6.131366, 6.152376, 6.161618, 6.164439, 
    6.165614 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.35703e-08, 6.384985e-08, 6.379551e-08, 6.402099e-08, 6.389591e-08, 
    6.404356e-08, 6.362697e-08, 6.386096e-08, 6.371158e-08, 6.359546e-08, 
    6.445858e-08, 6.403105e-08, 6.490264e-08, 6.462999e-08, 6.531489e-08, 
    6.486022e-08, 6.540657e-08, 6.530176e-08, 6.561717e-08, 6.552681e-08, 
    6.593026e-08, 6.565888e-08, 6.613939e-08, 6.586544e-08, 6.59083e-08, 
    6.564993e-08, 6.411708e-08, 6.440536e-08, 6.410001e-08, 6.414111e-08, 
    6.412267e-08, 6.38985e-08, 6.378554e-08, 6.354892e-08, 6.359188e-08, 
    6.376565e-08, 6.41596e-08, 6.402587e-08, 6.436288e-08, 6.435527e-08, 
    6.473046e-08, 6.45613e-08, 6.519191e-08, 6.501268e-08, 6.553059e-08, 
    6.540034e-08, 6.552447e-08, 6.548683e-08, 6.552496e-08, 6.533394e-08, 
    6.541578e-08, 6.524769e-08, 6.459298e-08, 6.47854e-08, 6.421152e-08, 
    6.386645e-08, 6.363724e-08, 6.347459e-08, 6.349758e-08, 6.354141e-08, 
    6.376668e-08, 6.397845e-08, 6.413985e-08, 6.424781e-08, 6.435418e-08, 
    6.467617e-08, 6.484658e-08, 6.522815e-08, 6.515928e-08, 6.527594e-08, 
    6.538738e-08, 6.557449e-08, 6.554369e-08, 6.562612e-08, 6.527286e-08, 
    6.550764e-08, 6.512006e-08, 6.522607e-08, 6.438312e-08, 6.406194e-08, 
    6.392545e-08, 6.380596e-08, 6.351526e-08, 6.371601e-08, 6.363688e-08, 
    6.382514e-08, 6.394477e-08, 6.38856e-08, 6.425076e-08, 6.41088e-08, 
    6.485669e-08, 6.453455e-08, 6.537438e-08, 6.517342e-08, 6.542255e-08, 
    6.529542e-08, 6.551326e-08, 6.531721e-08, 6.565681e-08, 6.573075e-08, 
    6.568022e-08, 6.587433e-08, 6.530634e-08, 6.552447e-08, 6.388395e-08, 
    6.389359e-08, 6.393855e-08, 6.374094e-08, 6.372885e-08, 6.354775e-08, 
    6.370889e-08, 6.377751e-08, 6.39517e-08, 6.405474e-08, 6.415268e-08, 
    6.436803e-08, 6.460854e-08, 6.494484e-08, 6.518644e-08, 6.53484e-08, 
    6.524908e-08, 6.533676e-08, 6.523875e-08, 6.519281e-08, 6.570305e-08, 
    6.541654e-08, 6.584641e-08, 6.582263e-08, 6.562809e-08, 6.58253e-08, 
    6.390037e-08, 6.384484e-08, 6.365205e-08, 6.380292e-08, 6.352803e-08, 
    6.36819e-08, 6.377039e-08, 6.411177e-08, 6.418676e-08, 6.425632e-08, 
    6.439367e-08, 6.456996e-08, 6.48792e-08, 6.514825e-08, 6.539386e-08, 
    6.537586e-08, 6.53822e-08, 6.543707e-08, 6.530116e-08, 6.545939e-08, 
    6.548594e-08, 6.541651e-08, 6.581944e-08, 6.570433e-08, 6.582212e-08, 
    6.574717e-08, 6.386289e-08, 6.395633e-08, 6.390584e-08, 6.400078e-08, 
    6.39339e-08, 6.423132e-08, 6.432049e-08, 6.473773e-08, 6.456649e-08, 
    6.483902e-08, 6.459417e-08, 6.463756e-08, 6.484792e-08, 6.46074e-08, 
    6.513343e-08, 6.477681e-08, 6.543921e-08, 6.508311e-08, 6.546152e-08, 
    6.53928e-08, 6.550658e-08, 6.560848e-08, 6.573668e-08, 6.597322e-08, 
    6.591844e-08, 6.611626e-08, 6.409562e-08, 6.421681e-08, 6.420614e-08, 
    6.433297e-08, 6.442676e-08, 6.463005e-08, 6.49561e-08, 6.483349e-08, 
    6.505858e-08, 6.510377e-08, 6.47618e-08, 6.497177e-08, 6.429792e-08, 
    6.44068e-08, 6.434197e-08, 6.410518e-08, 6.486175e-08, 6.447348e-08, 
    6.519043e-08, 6.498011e-08, 6.559395e-08, 6.528868e-08, 6.588829e-08, 
    6.614464e-08, 6.638587e-08, 6.66678e-08, 6.428295e-08, 6.42006e-08, 
    6.434804e-08, 6.455205e-08, 6.474131e-08, 6.499293e-08, 6.501867e-08, 
    6.506582e-08, 6.518791e-08, 6.529058e-08, 6.508073e-08, 6.531631e-08, 
    6.443206e-08, 6.489545e-08, 6.416948e-08, 6.438809e-08, 6.454002e-08, 
    6.447337e-08, 6.481947e-08, 6.490105e-08, 6.523254e-08, 6.506118e-08, 
    6.608137e-08, 6.563001e-08, 6.688245e-08, 6.653246e-08, 6.417183e-08, 
    6.428267e-08, 6.466841e-08, 6.448487e-08, 6.500973e-08, 6.513893e-08, 
    6.524394e-08, 6.53782e-08, 6.539269e-08, 6.547224e-08, 6.534189e-08, 
    6.546708e-08, 6.499347e-08, 6.520511e-08, 6.462431e-08, 6.476568e-08, 
    6.470064e-08, 6.46293e-08, 6.484947e-08, 6.508403e-08, 6.508903e-08, 
    6.516425e-08, 6.537621e-08, 6.501185e-08, 6.613964e-08, 6.544317e-08, 
    6.440352e-08, 6.461701e-08, 6.464749e-08, 6.456479e-08, 6.512597e-08, 
    6.492264e-08, 6.54703e-08, 6.532228e-08, 6.55648e-08, 6.544429e-08, 
    6.542655e-08, 6.527178e-08, 6.517542e-08, 6.493197e-08, 6.473388e-08, 
    6.457679e-08, 6.461332e-08, 6.478587e-08, 6.509838e-08, 6.5394e-08, 
    6.532925e-08, 6.554637e-08, 6.497167e-08, 6.521266e-08, 6.511952e-08, 
    6.536237e-08, 6.483023e-08, 6.528341e-08, 6.471441e-08, 6.476429e-08, 
    6.49186e-08, 6.522901e-08, 6.529767e-08, 6.5371e-08, 6.532575e-08, 
    6.510631e-08, 6.507035e-08, 6.491485e-08, 6.487192e-08, 6.475343e-08, 
    6.465533e-08, 6.474496e-08, 6.483909e-08, 6.51064e-08, 6.534729e-08, 
    6.560993e-08, 6.56742e-08, 6.598109e-08, 6.573129e-08, 6.614352e-08, 
    6.579306e-08, 6.639972e-08, 6.530966e-08, 6.578274e-08, 6.492562e-08, 
    6.501796e-08, 6.518498e-08, 6.556804e-08, 6.536123e-08, 6.560308e-08, 
    6.506895e-08, 6.479183e-08, 6.472012e-08, 6.458635e-08, 6.472317e-08, 
    6.471205e-08, 6.484298e-08, 6.480091e-08, 6.511527e-08, 6.494641e-08, 
    6.542611e-08, 6.560117e-08, 6.609553e-08, 6.639859e-08, 6.670707e-08, 
    6.684326e-08, 6.688472e-08, 6.690204e-08 ;

 ERRH2O =
  -22838.9, -22872.69, -22866.07, -22893.73, -22878.32, -22896.52, -22845.69, 
    -22874.05, -22855.89, -22841.91, -22948.64, -22894.97, -23006.07, 
    -22970.56, -23060.47, -23000.49, -23072.79, -23058.71, -23101.47, 
    -23089.11, -23145.09, -23107.21, -23174.93, -23135.95, -23141.98, 
    -23105.98, -22905.66, -22941.89, -22903.53, -22908.65, -22906.35, 
    -22878.64, -22864.86, -22836.34, -22841.48, -22862.44, -22910.96, 
    -22894.33, -22936.51, -22935.55, -22983.56, -22961.74, -23044.08, 
    -23020.52, -23089.62, -23071.95, -23088.79, -23083.66, -23088.85, 
    -23063.02, -23074.03, -23051.49, -22965.8, -22990.71, -22917.47, 
    -22874.72, -22846.93, -22827.49, -22830.22, -22835.45, -22862.56, 
    -22888.47, -22908.5, -22922.03, -22935.42, -22976.53, -22998.71, 
    -23048.89, -23039.77, -23055.26, -23070.2, -23095.62, -23091.41, 
    -23102.7, -23054.85, -23086.49, -23034.59, -23048.62, -22939.08, 
    -22898.8, -22881.95, -22867.34, -22832.33, -22856.43, -22846.88, 
    -22869.67, -22884.32, -22877.06, -22922.4, -22904.62, -23000.03, 
    -22958.32, -23068.45, -23041.64, -23074.95, -23057.86, -23087.26, 
    -23060.77, -23106.92, -23117.15, -23110.15, -23137.2, -23059.32, 
    -23088.79, -22876.86, -22878.04, -22883.56, -22859.44, -22857.98, 
    -22836.21, -22855.56, -22863.88, -22885.17, -22897.9, -22910.1, 
    -22937.17, -22967.8, -23011.64, -23043.36, -23064.96, -23051.68, 
    -23063.39, -23050.3, -23044.2, -23113.31, -23074.14, -23133.28, 
    -23129.95, -23102.97, -23130.32, -22878.87, -22872.08, -22848.71, 
    -22866.97, -22833.85, -22852.31, -22863.01, -22905, -22914.36, -22923.1, 
    -22940.41, -22962.85, -23002.98, -23038.31, -23071.07, -23068.65, 
    -23069.5, -23076.91, -23058.63, -23079.94, -23083.54, -23074.13, 
    -23129.5, -23113.49, -23129.88, -23119.43, -22874.28, -22885.74, 
    -22879.54, -22891.23, -22882.99, -22919.96, -22931.18, -22984.5, 
    -22962.4, -22997.71, -22965.96, -22971.54, -22998.88, -22967.66, 
    -23036.36, -22989.59, -23077.2, -23029.74, -23080.22, -23070.93, 
    -23086.35, -23100.28, -23117.97, -23151.17, -23143.41, -23171.6, 
    -22902.98, -22918.13, -22916.79, -22932.74, -22944.6, -22970.57, 
    -23013.12, -22996.99, -23026.52, -23032.45, -22987.63, -23015.19, 
    -22928.34, -22942.07, -22933.88, -22904.17, -23000.7, -22950.53, 
    -23043.89, -23016.27, -23098.29, -23056.96, -23139.16, -23175.69, 
    -23210.78, -23252.55, -22926.46, -22916.1, -22934.64, -22960.56, 
    -22984.96, -23017.95, -23021.3, -23027.47, -23043.55, -23057.21, 
    -23029.43, -23060.65, -22945.27, -23005.12, -22912.2, -22939.7, 
    -22959.02, -22950.51, -22995.15, -23005.86, -23049.48, -23026.86, 
    -23166.59, -23103.24, -23284.68, -23232.52, -22912.49, -22926.42, 
    -22975.52, -22951.98, -23020.13, -23037.08, -23050.99, -23068.96, 
    -23070.92, -23081.68, -23064.08, -23080.98, -23018.01, -23045.84, 
    -22969.83, -22988.13, -22979.69, -22970.47, -22999.08, -23029.86, 
    -23030.51, -23040.42, -23068.71, -23020.41, -23174.97, -23077.75, 
    -22941.65, -22968.9, -22972.82, -22962.19, -23035.37, -23008.71, 
    -23081.41, -23061.45, -23094.29, -23077.89, -23075.49, -23054.7, 
    -23041.9, -23009.94, -22984, -22963.72, -22968.42, -22990.77, -23031.74, 
    -23071.1, -23062.39, -23091.78, -23015.18, -23046.84, -23034.52, 
    -23066.84, -22996.56, -23056.26, -22981.47, -22987.95, -23008.17, 
    -23049.01, -23058.16, -23068, -23061.92, -23032.79, -23028.06, -23007.68, 
    -23002.03, -22986.54, -22973.83, -22985.44, -22997.72, -23032.8, 
    -23064.81, -23100.48, -23109.32, -23152.29, -23117.23, -23175.53, 
    -23125.83, -23212.83, -23059.77, -23124.38, -23009.1, -23021.21, 
    -23043.17, -23094.74, -23066.68, -23099.54, -23027.88, -22991.54, 
    -22982.21, -22964.95, -22982.61, -22981.17, -22998.23, -22992.73, 
    -23033.96, -23011.84, -23075.43, -23099.28, -23168.62, -23212.65, 
    -23258.39, -23278.77, -23285.02, -23287.64 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -8.348114e-15, -1.586967e-14, -3.442384e-15, -1.071295e-14, -4.805658e-15, 
    -9.866948e-15, -4.221674e-15, -8.139908e-15, -5.389951e-15, 3.609534e-15, 
    -9.485775e-15, -5.411627e-15, -9.156754e-15, -1.71168e-14, -6.169292e-15, 
    -1.412968e-14, -1.54606e-14, -1.15268e-14, -1.165566e-14, -9.061214e-15, 
    -7.190861e-15, -1.268688e-14, -6.892944e-15, -3.985732e-15, 
    -6.398813e-15, -1.513341e-14, -1.137361e-14, -1.120921e-14, 
    -3.744321e-15, -7.786798e-15, -1.605037e-14, 7.1917e-15, -1.045874e-14, 
    -5.196141e-15, 8.883934e-16, -5.711458e-15, -7.467254e-15, -8.894596e-15, 
    -9.94981e-15, -1.294084e-14, -1.127619e-14, -9.664925e-15, -8.540095e-15, 
    1.116947e-15, -1.389908e-14, -6.87208e-15, -4.101396e-15, -9.769512e-15, 
    -1.62681e-14, -2.699553e-14, -7.900464e-16, -1.282021e-14, -6.096806e-15, 
    -4.419164e-15, -5.980964e-15, -5.579279e-15, -1.328882e-14, -9.32534e-16, 
    -8.985624e-15, -5.527674e-15, -5.228842e-15, -1.1977e-14, -3.357852e-15, 
    -7.740877e-15, -1.924561e-14, -7.700954e-15, -5.434426e-15, 
    -1.187856e-14, 4.843782e-15, -1.147857e-14, -1.995298e-14, -3.562995e-16, 
    3.227385e-15, -1.037076e-15, -1.720626e-16, -3.685503e-15, -1.257123e-14, 
    -1.210948e-14, -6.232559e-15, -1.021386e-14, -3.735155e-15, 
    -4.563317e-15, -2.067855e-14, -1.153012e-15, -8.390705e-15, 3.155986e-15, 
    -1.938236e-14, -1.152038e-14, 7.43574e-15, -1.909292e-14, -9.743793e-15, 
    -1.417202e-14, -1.643047e-14, -5.312555e-15, -8.47719e-15, -1.143322e-14, 
    -8.388498e-15, -1.782754e-14, -1.568844e-15, -4.827628e-15, 
    -1.085027e-14, -1.25811e-14, -2.446065e-15, -6.4768e-15, -1.607307e-14, 
    -1.816957e-15, -4.115905e-15, -8.849487e-15, -8.723576e-16, 
    -1.618428e-14, -5.903159e-15, -9.150806e-15, 4.53039e-15, -4.242274e-15, 
    -1.002012e-14, -9.63548e-15, -1.314983e-14, 8.743386e-17, -7.750347e-15, 
    -1.030234e-14, -7.858288e-15, -1.671538e-14, 1.879499e-15, -6.137e-15, 
    -4.689643e-15, -2.007377e-15, -2.813418e-15, -1.093519e-14, 
    -5.782515e-15, -1.092057e-14, -8.789512e-15, -1.328565e-14, 
    -9.264811e-16, -9.541495e-15, -1.873744e-14, -2.271684e-14, 
    -1.285887e-14, -4.016984e-15, -7.638175e-15, -4.863249e-15, 5.158376e-17, 
    2.551585e-16, -8.814216e-15, -5.251001e-15, -8.005607e-15, -1.405661e-14, 
    -2.128678e-14, -1.335069e-14, 4.769759e-15, -1.279543e-14, -7.280362e-15, 
    -3.733775e-15, -1.411091e-14, -3.539073e-15, -9.98526e-15, -2.114768e-14, 
    -7.516209e-15, -1.676181e-15, -2.391082e-15, -7.655426e-15, 
    -1.873267e-17, -6.90472e-15, -7.649008e-15, -2.445431e-15, 4.526449e-17, 
    1.142812e-16, -1.415156e-14, 5.008966e-15, -1.416807e-14, -9.551043e-15, 
    -1.288815e-14, -2.195079e-15, -1.290682e-14, -8.204673e-15, 8.615541e-17, 
    -2.414148e-15, -5.41008e-15, -9.727988e-15, -5.763864e-15, -3.934501e-15, 
    -1.299808e-14, -1.873758e-15, -9.503391e-15, -8.522214e-15, 
    -1.057797e-14, 1.210534e-15, -2.129679e-14, -5.689167e-15, -1.106546e-14, 
    -3.701911e-15, -9.408808e-15, -9.626213e-15, -1.650854e-14, 
    -9.328985e-15, -8.448236e-15, -7.809566e-15, -1.976484e-14, 1.019171e-15, 
    -2.914441e-15, -1.738273e-14, -8.672185e-15, -1.342646e-14, 
    -7.539713e-15, -1.63801e-14, -1.303487e-14, -4.981659e-15, -1.846204e-14, 
    -9.899468e-15, -8.19148e-15, -2.061223e-15, -1.436333e-14, 1.961061e-16, 
    -6.239847e-15, -3.194545e-15, -1.051708e-14, -1.309758e-14, 
    -1.657611e-14, 1.22034e-15, 3.727681e-15, -1.039776e-14, -1.013163e-14, 
    -1.283912e-14, -6.039891e-15, -6.831997e-15, -7.62411e-15, -9.176824e-15, 
    -5.886882e-15, -1.537996e-14, -5.859297e-15, -1.062457e-15, 
    -1.372585e-14, -5.767694e-15, -3.124784e-15, -3.298095e-16, 
    -8.000598e-15, 7.352073e-16, -2.0944e-14, -9.474468e-15, -5.803262e-15, 
    -2.73684e-15, -7.80647e-15, -6.795157e-15, -1.113083e-14, -5.233233e-15, 
    -4.55147e-15, 2.848085e-15, -1.70473e-14, -1.263116e-14, -8.296036e-15, 
    -4.044563e-15, -7.332795e-15, -1.043971e-14, -1.168761e-14, 
    -1.162579e-14, -7.872686e-15, -8.1056e-15, -3.9113e-15, -5.295914e-15, 
    -2.372948e-15, -1.659397e-15, -5.21969e-15, -8.453261e-15, -4.728962e-15, 
    -3.625063e-15, -1.708585e-14, -1.192769e-14, -8.205782e-15, 
    -1.150572e-14, -4.213074e-15, -1.396359e-14, -1.382551e-14, 
    -1.674421e-15, -1.170342e-14, -6.729986e-15, -1.128886e-14, -5.71551e-15, 
    -9.960265e-15, -4.220877e-15, -8.114002e-15, -2.182516e-15, 
    -1.140627e-14, -3.424737e-15, -8.598432e-15, -8.693252e-15, 
    -1.383226e-14, -9.377093e-15, -4.312672e-15, -9.712468e-15, 
    -1.425938e-14, -5.103328e-15, -1.006598e-14, -1.028555e-15, 
    -4.119142e-15, -2.214025e-15, -1.244426e-14, -1.19595e-14, -1.636929e-14, 
    -1.736289e-14, -4.166122e-15, -9.891205e-15, -1.424593e-14, 
    -1.239449e-14, -2.2548e-15, -1.099184e-14, -1.007138e-14, -1.178245e-14, 
    -1.51793e-14, -1.106158e-14, -3.53206e-15, -1.042393e-14, -8.980131e-15, 
    -1.383896e-14, -9.380093e-15, -1.084424e-14, -1.016928e-14, 
    -1.625197e-14, -1.908403e-14, 2.403012e-16, -8.829729e-15, -1.120049e-14, 
    -1.964229e-15, -1.211814e-14, -9.675679e-15, -1.53372e-14, -6.541565e-15, 
    -1.620455e-14, -1.039189e-14, -8.267922e-15, 3.822316e-16, -1.844392e-14, 
    2.082029e-15, -1.404304e-14, -1.386469e-14, -1.182944e-14, -1.540235e-14, 
    -4.038333e-15, -6.337426e-15, -8.367988e-15 ;

 ERRSOI =
  -1.463665e-10, -3.285682e-10, -2.402727e-10, -3.806203e-10, -4.156693e-10, 
    -3.035628e-10, -3.407355e-10, -4.214056e-10, -2.785323e-10, 
    -2.219673e-10, -3.583683e-10, -2.504875e-10, -4.188541e-10, 
    -3.082031e-10, -4.154015e-10, -1.793197e-10, -4.312842e-10, 
    -4.275549e-10, -4.772648e-10, -1.562107e-10, -4.83723e-10, -1.340446e-10, 
    -3.293612e-10, -2.717691e-10, -4.505432e-10, -1.988107e-10, 
    -3.567269e-10, -2.720598e-10, -7.247805e-11, -2.148665e-10, 
    -3.733183e-10, -2.474676e-10, -1.98089e-10, -4.487216e-10, -2.949428e-10, 
    -3.71151e-10, -2.711487e-10, -2.883507e-10, -3.801915e-10, -1.242798e-10, 
    -2.83018e-10, -3.67273e-10, -3.015647e-10, -4.235771e-10, -2.85014e-10, 
    -3.245127e-10, -3.597861e-10, -2.695899e-10, -3.114433e-10, 
    -3.302414e-10, -1.894569e-10, -3.436503e-10, -3.588237e-10, 
    -4.029105e-10, -3.083129e-10, -2.785931e-10, -1.041047e-10, 
    -4.920947e-10, -2.527903e-10, -1.421995e-10, -3.845356e-10, -3.44954e-10, 
    -3.100044e-10, -4.479887e-10, -4.064445e-10, -1.499516e-10, 
    -2.801204e-10, -2.243355e-10, -1.587996e-10, -3.031422e-10, 
    -2.233396e-10, -3.829675e-10, -3.370772e-10, -1.162475e-10, 
    -3.113385e-10, -3.274061e-10, -2.851581e-10, -2.771008e-10, 
    -5.153366e-10, -2.497724e-10, -3.252895e-10, -1.57017e-10, -3.03762e-10, 
    -4.915555e-10, -3.62523e-10, -3.412347e-10, -4.698499e-10, -3.749813e-10, 
    -4.928467e-10, -2.315992e-10, -2.257639e-10, -3.320692e-10, 
    -3.285422e-10, -3.735216e-10, -3.233517e-10, -3.169199e-10, -5.22987e-10, 
    -3.095116e-10, -1.117901e-10, -1.144016e-10, -3.576668e-10, 
    -4.014212e-10, -3.949618e-10, -1.372473e-10, -3.551838e-10, 
    -2.514429e-10, -2.069968e-10, -4.369355e-10, -1.168311e-10, 
    -3.939719e-10, -1.91631e-10, -2.467957e-10, -2.177587e-10, -2.918118e-10, 
    -2.178247e-10, -4.989698e-10, -9.374196e-11, -2.305645e-10, 
    -3.997654e-10, -2.95686e-10, -3.764148e-10, -2.534091e-10, -2.745322e-10, 
    -2.575442e-10, -1.663193e-10, -2.461582e-10, -2.651658e-10, 
    -1.819184e-10, -2.220848e-10, -1.900467e-10, -5.051403e-10, 
    -3.632036e-10, -2.889496e-10, -4.020503e-10, -3.887717e-10, 
    -2.760275e-10, -1.203674e-10, -1.712231e-10, -2.658708e-10, 
    -3.152734e-10, -2.216363e-10, -4.012135e-10, -4.145285e-10, 
    -2.526675e-10, -3.384065e-10, -2.399708e-10, -3.257762e-10, 
    -2.433745e-10, -3.533057e-10, -2.329415e-10, -3.50018e-10, -1.704943e-10, 
    -3.163618e-10, -2.707543e-10, -1.278956e-10, -2.323683e-10, 
    -2.371671e-10, -2.63167e-10, -3.744735e-10, -3.62785e-10, -4.282597e-10, 
    -4.544037e-10, -3.057926e-10, -1.531681e-10, -2.351515e-10, 
    -2.658689e-10, -2.544232e-10, -2.723065e-10, -2.917489e-10, 
    -5.076827e-11, -2.921544e-10, -2.357837e-10, -2.579116e-10, 
    -4.525316e-10, -3.32299e-10, -2.895421e-10, -2.548859e-10, -2.777509e-10, 
    -3.044502e-10, -1.876364e-10, -2.901947e-10, -3.450951e-10, -1.60813e-10, 
    -2.419373e-10, -2.693658e-10, -2.496031e-10, -2.809786e-10, 
    -3.178058e-10, -2.201073e-10, -2.903568e-10, -1.73104e-10, -3.427204e-10, 
    -1.630159e-10, -3.232892e-10, -2.708674e-10, -4.9013e-10, -3.034757e-10, 
    -2.872557e-10, -2.961284e-10, -4.658963e-10, -3.324355e-10, 
    -1.364723e-10, -1.797155e-10, -5.257761e-10, -2.658016e-10, 
    -1.639401e-10, -2.596249e-10, -2.896056e-10, -1.439682e-10, 
    -2.820994e-10, -2.882888e-10, -4.2596e-10, -2.677377e-10, -3.402184e-10, 
    -3.344288e-10, -4.810421e-10, -3.895747e-10, -3.270246e-10, 
    -2.650637e-10, -2.751441e-10, -2.570678e-10, -3.58209e-10, -1.751343e-10, 
    -2.913369e-10, -3.37842e-10, -4.858534e-10, -1.636431e-10, -1.187508e-10, 
    -2.91542e-10, -1.115481e-10, -1.679268e-10, -3.461383e-10, -2.172521e-10, 
    -3.131535e-10, -3.361008e-10, -4.007736e-10, -3.563579e-11, -3.48259e-10, 
    -3.010653e-10, -3.619382e-10, -1.393226e-10, -2.139709e-10, 
    -1.282455e-10, -2.410242e-10, -4.002239e-10, -2.105929e-10, 
    -1.592342e-10, -2.939113e-10, -1.318032e-10, -2.426753e-10, 
    -8.897498e-11, -3.672747e-10, -3.744833e-10, -2.940253e-10, 
    -2.631049e-10, -2.042045e-10, -2.180092e-10, -2.109981e-10, 
    -3.704768e-10, -2.824903e-10, -3.456467e-10, -2.654363e-10, 
    -4.256896e-10, -1.951895e-10, -1.237515e-10, -9.367863e-11, 
    -3.360604e-10, -3.240892e-10, -5.609841e-11, -4.193472e-10, 
    -2.845609e-10, -2.729359e-10, -5.027276e-10, -3.089464e-10, 
    -3.044654e-10, -1.687855e-10, -9.32005e-11, -2.224902e-10, -3.698706e-10, 
    -2.840219e-10, -2.24872e-10, -2.505423e-10, -3.226286e-10, -3.049315e-10, 
    -2.811213e-10, -2.839987e-10, -2.509769e-10, -1.938582e-10, 
    -3.069898e-10, -1.950099e-10, -2.502145e-10, -3.895025e-10, 
    -3.068039e-10, -3.265024e-10, -3.057234e-10, -2.418445e-10, 
    -2.397215e-10, -4.908422e-10, -3.797179e-10, -4.592836e-10, 
    -1.640084e-10, -8.857933e-11, -3.729312e-10, -3.414955e-10, 
    -4.554823e-10, -3.261105e-10, -1.560804e-10, -2.69035e-10, -1.428743e-10, 
    -3.387063e-10, -2.111248e-10, -1.411183e-10, -3.402778e-10, 
    -1.728749e-10, -4.944516e-10, -3.491294e-10, -3.028549e-10, 
    -1.996944e-10, -3.202727e-10, -4.920493e-10, -2.949051e-10, 
    -2.972657e-10, -3.262819e-10, -3.431396e-10, -1.533341e-10, 
    -9.955519e-11, -3.677172e-10, -2.107575e-10, -3.270838e-10, 
    -2.872302e-10, -2.71575e-10, -2.437415e-10, -2.663367e-10, -2.036499e-10, 
    -2.989417e-10, -4.837253e-10, -8.51638e-11, -1.295576e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.62123, -1.620132, -1.62034, -1.619464, -1.619942, -1.619374, -1.620997, 
    -1.620097, -1.620666, -1.621117, -1.617783, -1.619422, -1.615993, 
    -1.617049, -1.614362, -1.616171, -1.61399, -1.614392, -1.613124, 
    -1.613487, -1.611906, -1.612957, -1.611043, -1.612145, -1.611982, 
    -1.612995, -1.619071, -1.617995, -1.61914, -1.618986, -1.61905, -1.61994, 
    -1.620402, -1.621298, -1.621131, -1.620465, -1.618916, -1.619428, 
    -1.618091, -1.61812, -1.616651, -1.617312, -1.614829, -1.615528, 
    -1.613471, -1.613996, -1.6135, -1.613647, -1.613498, -1.614265, 
    -1.613938, -1.614604, -1.617193, -1.61644, -1.618704, -1.620097, 
    -1.620962, -1.62159, -1.621502, -1.621337, -1.620461, -1.619615, 
    -1.618974, -1.618549, -1.618125, -1.616908, -1.616214, -1.614698, 
    -1.614954, -1.614505, -1.614047, -1.613302, -1.613422, -1.613098, 
    -1.614502, -1.613577, -1.615099, -1.61469, -1.618088, -1.619286, 
    -1.61986, -1.620303, -1.621435, -1.620658, -1.620966, -1.620216, 
    -1.619748, -1.619976, -1.618537, -1.6191, -1.616173, -1.61743, -1.6141, 
    -1.6149, -1.613905, -1.614409, -1.613551, -1.614323, -1.612971, 
    -1.612684, -1.612882, -1.612094, -1.614368, -1.613508, -1.619986, 
    -1.61995, -1.619769, -1.620562, -1.620606, -1.621306, -1.620676, 
    -1.620414, -1.619715, -1.619315, -1.61893, -1.618078, -1.617143, 
    -1.615814, -1.614849, -1.614199, -1.614592, -1.614245, -1.614636, 
    -1.614816, -1.612797, -1.61394, -1.612208, -1.612301, -1.613093, 
    -1.612291, -1.619923, -1.620136, -1.620901, -1.620303, -1.621381, 
    -1.620788, -1.620452, -1.619106, -1.61879, -1.618522, -1.617972, 
    -1.617279, -1.616071, -1.615008, -1.614017, -1.614088, -1.614064, 
    -1.61385, -1.61439, -1.61376, -1.613662, -1.613931, -1.612314, -1.612777, 
    -1.612303, -1.612603, -1.620065, -1.619702, -1.619899, -1.619532, 
    -1.619797, -1.618638, -1.618289, -1.616642, -1.617297, -1.616233, 
    -1.617183, -1.617019, -1.616231, -1.617126, -1.615077, -1.616498, 
    -1.613841, -1.615294, -1.613751, -1.614021, -1.613566, -1.613167, 
    -1.612648, -1.61171, -1.611925, -1.611125, -1.619152, -1.618685, 
    -1.618712, -1.618213, -1.617846, -1.617039, -1.61576, -1.616237, 
    -1.615345, -1.615171, -1.616517, -1.615705, -1.618362, -1.617946, 
    -1.618183, -1.619123, -1.616147, -1.617679, -1.614835, -1.615662, 
    -1.613226, -1.614459, -1.612046, -1.611044, -1.610027, -1.608912, 
    -1.618415, -1.618734, -1.618149, -1.617369, -1.616607, -1.615614, 
    -1.615504, -1.615322, -1.614836, -1.61443, -1.615278, -1.614326, 
    -1.617879, -1.616007, -1.618868, -1.618023, -1.617408, -1.617662, 
    -1.616288, -1.615968, -1.614676, -1.615334, -1.611305, -1.613103, 
    -1.608009, -1.609456, -1.618848, -1.618409, -1.616903, -1.617615, 
    -1.61554, -1.615033, -1.614613, -1.614091, -1.614024, -1.613712, 
    -1.614225, -1.613727, -1.615612, -1.614773, -1.617057, -1.616511, 
    -1.616757, -1.617038, -1.616171, -1.615269, -1.615226, -1.614945, 
    -1.614178, -1.615531, -1.611115, -1.613899, -1.61793, -1.617118, 
    -1.616974, -1.617293, -1.615085, -1.61589, -1.613717, -1.614303, 
    -1.613335, -1.613819, -1.613891, -1.614504, -1.614892, -1.615857, 
    -1.616638, -1.617244, -1.617101, -1.616435, -1.615208, -1.614029, 
    -1.614292, -1.613408, -1.615691, -1.614753, -1.615121, -1.614147, 
    -1.616255, -1.614534, -1.616703, -1.616508, -1.615905, -1.614705, 
    -1.614401, -1.61412, -1.614289, -1.615172, -1.615307, -1.615914, 
    -1.616094, -1.616549, -1.616935, -1.616588, -1.616227, -1.615162, 
    -1.614216, -1.613164, -1.612897, -1.611719, -1.612711, -1.611105, 
    -1.612521, -1.610038, -1.614399, -1.612514, -1.61587, -1.615505, 
    -1.614874, -1.613355, -1.614152, -1.613208, -1.61531, -1.616424, 
    -1.616682, -1.617211, -1.61667, -1.616713, -1.616195, -1.616361, 
    -1.615126, -1.615789, -1.613899, -1.613209, -1.611218, -1.610002, 
    -1.608717, -1.60816, -1.607988, -1.607918 ;

 FCH4 =
  1.827341e-13, 1.82682e-13, 1.826929e-13, 1.826451e-13, 1.826725e-13, 
    1.826399e-13, 1.827244e-13, 1.826797e-13, 1.82709e-13, 1.827299e-13, 
    1.825304e-13, 1.826427e-13, 1.823794e-13, 1.824767e-13, 1.811538e-13, 
    1.823955e-13, 1.811598e-13, 1.811527e-13, 1.8116e-13, 1.811623e-13, 
    1.811236e-13, 1.811578e-13, 1.810734e-13, 1.811349e-13, 1.811276e-13, 
    1.811583e-13, 1.826225e-13, 1.82546e-13, 1.826266e-13, 1.826166e-13, 
    1.826211e-13, 1.826719e-13, 1.826949e-13, 1.827378e-13, 1.827305e-13, 
    1.826987e-13, 1.82612e-13, 1.82644e-13, 1.825582e-13, 1.825604e-13, 
    1.824426e-13, 1.824989e-13, 1.811404e-13, 1.8111e-13, 1.811623e-13, 
    1.811595e-13, 1.811623e-13, 1.811622e-13, 1.811623e-13, 1.811554e-13, 
    1.811602e-13, 1.811472e-13, 1.824888e-13, 1.824231e-13, 1.825989e-13, 
    1.826786e-13, 1.827226e-13, 1.827499e-13, 1.827462e-13, 1.82739e-13, 
    1.826986e-13, 1.826546e-13, 1.826169e-13, 1.825895e-13, 1.825607e-13, 
    1.824612e-13, 1.824007e-13, 1.811449e-13, 1.811358e-13, 1.811502e-13, 
    1.811589e-13, 1.811615e-13, 1.811621e-13, 1.811596e-13, 1.811499e-13, 
    1.811623e-13, 1.811297e-13, 1.811447e-13, 1.825523e-13, 1.826356e-13, 
    1.826661e-13, 1.826909e-13, 1.827433e-13, 1.827082e-13, 1.827226e-13, 
    1.82687e-13, 1.82662e-13, 1.826747e-13, 1.825887e-13, 1.826245e-13, 
    1.823969e-13, 1.825073e-13, 1.811581e-13, 1.811378e-13, 1.811605e-13, 
    1.811521e-13, 1.811623e-13, 1.81154e-13, 1.811579e-13, 1.81152e-13, 
    1.811563e-13, 1.811335e-13, 1.811531e-13, 1.811623e-13, 1.82675e-13, 
    1.82673e-13, 1.826634e-13, 1.827035e-13, 1.827058e-13, 1.82738e-13, 
    1.827095e-13, 1.826965e-13, 1.826605e-13, 1.826373e-13, 1.826138e-13, 
    1.825568e-13, 1.824837e-13, 1.82363e-13, 1.811396e-13, 1.811564e-13, 
    1.811474e-13, 1.811556e-13, 1.811462e-13, 1.811405e-13, 1.811545e-13, 
    1.811602e-13, 1.811378e-13, 1.811413e-13, 1.811595e-13, 1.811409e-13, 
    1.826715e-13, 1.826831e-13, 1.827199e-13, 1.826915e-13, 1.827412e-13, 
    1.827145e-13, 1.826978e-13, 1.826237e-13, 1.826052e-13, 1.825873e-13, 
    1.825495e-13, 1.824962e-13, 1.823884e-13, 1.811341e-13, 1.811592e-13, 
    1.811582e-13, 1.811586e-13, 1.81161e-13, 1.811526e-13, 1.811617e-13, 
    1.811621e-13, 1.811603e-13, 1.811417e-13, 1.811544e-13, 1.811413e-13, 
    1.811504e-13, 1.826794e-13, 1.826595e-13, 1.826704e-13, 1.826496e-13, 
    1.826644e-13, 1.825938e-13, 1.825699e-13, 1.824401e-13, 1.824973e-13, 
    1.824035e-13, 1.824884e-13, 1.824742e-13, 1.824001e-13, 1.824841e-13, 
    1.811318e-13, 1.824262e-13, 1.811611e-13, 1.811234e-13, 1.811617e-13, 
    1.811592e-13, 1.811623e-13, 1.811604e-13, 1.811514e-13, 1.81115e-13, 
    1.811258e-13, 1.810801e-13, 1.826276e-13, 1.825975e-13, 1.826003e-13, 
    1.825666e-13, 1.825399e-13, 1.824767e-13, 1.823586e-13, 1.824056e-13, 
    1.81119e-13, 1.81127e-13, 1.824316e-13, 1.823524e-13, 1.825761e-13, 
    1.825456e-13, 1.82564e-13, 1.826253e-13, 1.82395e-13, 1.82526e-13, 
    1.811402e-13, 1.82349e-13, 1.811609e-13, 1.811515e-13, 1.811311e-13, 
    1.810718e-13, 1.809862e-13, 1.808471e-13, 1.825802e-13, 1.826017e-13, 
    1.825624e-13, 1.825018e-13, 1.824388e-13, 1.823439e-13, 1.811113e-13, 
    1.811203e-13, 1.811399e-13, 1.811517e-13, 1.81123e-13, 1.81154e-13, 
    1.825382e-13, 1.823822e-13, 1.826096e-13, 1.82551e-13, 1.825056e-13, 
    1.82526e-13, 1.824108e-13, 1.823801e-13, 1.811455e-13, 1.811195e-13, 
    1.810894e-13, 1.811594e-13, 1.807118e-13, 1.809192e-13, 1.82609e-13, 
    1.825803e-13, 1.824639e-13, 1.825226e-13, 1.811094e-13, 1.811327e-13, 
    1.811468e-13, 1.811583e-13, 1.811591e-13, 1.811619e-13, 1.81156e-13, 
    1.811618e-13, 1.823437e-13, 1.811421e-13, 1.824786e-13, 1.824302e-13, 
    1.82453e-13, 1.82477e-13, 1.823997e-13, 1.811236e-13, 1.811245e-13, 
    1.811365e-13, 1.811581e-13, 1.811099e-13, 1.810732e-13, 1.811611e-13, 
    1.825466e-13, 1.82481e-13, 1.824709e-13, 1.824978e-13, 1.811307e-13, 
    1.823718e-13, 1.811619e-13, 1.811544e-13, 1.811618e-13, 1.811613e-13, 
    1.811607e-13, 1.811498e-13, 1.811381e-13, 1.823681e-13, 1.824415e-13, 
    1.82494e-13, 1.824822e-13, 1.82423e-13, 1.811261e-13, 1.811592e-13, 
    1.81155e-13, 1.811621e-13, 1.823524e-13, 1.811431e-13, 1.811296e-13, 
    1.811574e-13, 1.824068e-13, 1.811508e-13, 1.824483e-13, 1.824307e-13, 
    1.823733e-13, 1.81145e-13, 1.811523e-13, 1.811579e-13, 1.811547e-13, 
    1.811274e-13, 1.811211e-13, 1.823748e-13, 1.823912e-13, 1.824346e-13, 
    1.824684e-13, 1.824376e-13, 1.824035e-13, 1.811275e-13, 1.811563e-13, 
    1.811603e-13, 1.811567e-13, 1.811133e-13, 1.811519e-13, 1.81072e-13, 
    1.811449e-13, 1.809802e-13, 1.811533e-13, 1.811463e-13, 1.823706e-13, 
    1.811111e-13, 1.811394e-13, 1.811616e-13, 1.811573e-13, 1.811606e-13, 
    1.811209e-13, 1.824208e-13, 1.824463e-13, 1.824909e-13, 1.824452e-13, 
    1.824491e-13, 1.824021e-13, 1.824176e-13, 1.811289e-13, 1.823625e-13, 
    1.811606e-13, 1.811607e-13, 1.810857e-13, 1.809808e-13, 1.808244e-13, 
    1.807385e-13, 1.807103e-13, 1.806982e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  7.56001, 7.577816, 7.574367, 7.588705, 7.58077, 7.590137, 7.563644, 
    7.578502, 7.56903, 7.561646, 7.616299, 7.589347, 7.644516, 7.627287, 
    7.672421, 7.641802, 7.678262, 7.671641, 7.691704, 7.685958, 7.711526, 
    7.694357, 7.72488, 7.707453, 7.710158, 7.693782, 7.59482, 7.612925, 
    7.593735, 7.596319, 7.595171, 7.580915, 7.573676, 7.558688, 7.561418, 
    7.572448, 7.597482, 7.589054, 7.610404, 7.609922, 7.633656, 7.622955, 
    7.664663, 7.651557, 7.686199, 7.677911, 7.6858, 7.683414, 7.685831, 
    7.673681, 7.678884, 7.668213, 7.624949, 7.637122, 7.600786, 7.578797, 
    7.564286, 7.553952, 7.555412, 7.558185, 7.572511, 7.586035, 7.596277, 
    7.60311, 7.609852, 7.630118, 7.640964, 7.666936, 7.662604, 7.669977, 
    7.67709, 7.688974, 7.687025, 7.692252, 7.669816, 7.684708, 7.658376, 
    7.666841, 7.611506, 7.591336, 7.582569, 7.575023, 7.556531, 7.56929, 
    7.564255, 7.576273, 7.583886, 7.580128, 7.603297, 7.594303, 7.641606, 
    7.621233, 7.67626, 7.663497, 7.679327, 7.671256, 7.685073, 7.672637, 
    7.694212, 7.698892, 7.695689, 7.708053, 7.671944, 7.685783, 7.580014, 
    7.580626, 7.583498, 7.570873, 7.570112, 7.558604, 7.56886, 7.573214, 
    7.584342, 7.590878, 7.597075, 7.610712, 7.625909, 7.647218, 7.664322, 
    7.674621, 7.668317, 7.67388, 7.667654, 7.664744, 7.697126, 7.678921, 
    7.706274, 7.704766, 7.692369, 7.704936, 7.581059, 7.577533, 7.565235, 
    7.574859, 7.557353, 7.567128, 7.572735, 7.594452, 7.599245, 7.603633, 
    7.612346, 7.623502, 7.643064, 7.661879, 7.677511, 7.676369, 7.676769, 
    7.680244, 7.671612, 7.681664, 7.683334, 7.67894, 7.704563, 7.697242, 
    7.704733, 7.699971, 7.578683, 7.584625, 7.581411, 7.587445, 7.583179, 
    7.60201, 7.607646, 7.63407, 7.623272, 7.64051, 7.625037, 7.627767, 
    7.640997, 7.625885, 7.659152, 7.636524, 7.68038, 7.655919, 7.6818, 
    7.677443, 7.684675, 7.691134, 7.699296, 7.714312, 7.710841, 7.723435, 
    7.593471, 7.601114, 7.600475, 7.6085, 7.614429, 7.627315, 7.647953, 
    7.640201, 7.654472, 7.657326, 7.635665, 7.64893, 7.606256, 7.613117, 
    7.609057, 7.594054, 7.641941, 7.617346, 7.66457, 7.649483, 7.690208, 
    7.670774, 7.708923, 7.725163, 7.740619, 7.75851, 7.605324, 7.600125, 
    7.609464, 7.622323, 7.634346, 7.650289, 7.651939, 7.654918, 7.664431, 
    7.670945, 7.655827, 7.672583, 7.61464, 7.644093, 7.598128, 7.611924, 
    7.62158, 7.61738, 7.639323, 7.644486, 7.667224, 7.654638, 7.721124, 
    7.692451, 7.772257, 7.7499, 7.5983, 7.605321, 7.629707, 7.618114, 
    7.651372, 7.659551, 7.66799, 7.676487, 7.67743, 7.682472, 7.674207, 
    7.682158, 7.650323, 7.665513, 7.626961, 7.63589, 7.631793, 7.627275, 
    7.641219, 7.656029, 7.656399, 7.662894, 7.676178, 7.651507, 7.724727, 
    7.680459, 7.612976, 7.626424, 7.62841, 7.62319, 7.658729, 7.645839, 
    7.682357, 7.672961, 7.688372, 7.680707, 7.679578, 7.669752, 7.663624, 
    7.646419, 7.633871, 7.623954, 7.626264, 7.63716, 7.656947, 7.677491, 
    7.673364, 7.687201, 7.648956, 7.665967, 7.658295, 7.675498, 7.639982, 
    7.670314, 7.632666, 7.635821, 7.645583, 7.666966, 7.671396, 7.67603, 
    7.673182, 7.65746, 7.655199, 7.64536, 7.642616, 7.635139, 7.628924, 
    7.634588, 7.640527, 7.657488, 7.67452, 7.691218, 7.695327, 7.714719, 
    7.698856, 7.724962, 7.702651, 7.741345, 7.672052, 7.702107, 7.646046, 
    7.651898, 7.664183, 7.688502, 7.675426, 7.690746, 7.655114, 7.637508, 
    7.633023, 7.624547, 7.633217, 7.632514, 7.640811, 7.638148, 7.658052, 
    7.647361, 7.679534, 7.690639, 7.722095, 7.741367, 7.761094, 7.769778, 
    7.772428, 7.773532 ;

 FGR =
  -370.0307, -370.701, -370.571, -371.1112, -370.8119, -371.1653, -370.1671, 
    -370.7272, -370.3699, -370.0917, -372.1567, -371.1354, -373.2167, 
    -372.5682, -374.2104, -373.1152, -374.4292, -374.1802, -374.9322, 
    -374.7168, -375.6767, -375.0316, -376.1761, -375.5231, -375.6249, 
    -375.0101, -371.3419, -372.0292, -371.301, -371.399, -371.3553, 
    -370.8177, -370.546, -369.9803, -370.0832, -370.4991, -371.4431, 
    -371.1237, -371.931, -371.9128, -372.8076, -372.4049, -373.9185, -373.48, 
    -374.7258, -374.4153, -374.711, -374.6215, -374.7122, -374.2568, 
    -374.4518, -374.0515, -372.4802, -372.9382, -371.5678, -370.7393, 
    -370.1915, -369.802, -369.857, -369.9618, -370.5015, -371.01, -371.3968, 
    -371.6552, -371.9101, -372.6764, -373.0832, -374.0043, -373.841, 
    -374.1183, -374.3844, -374.8301, -374.7569, -374.9531, -374.1116, 
    -374.6705, -373.7359, -374, -371.9757, -371.21, -370.8811, -370.5959, 
    -369.8993, -370.3801, -370.1905, -370.6424, -370.9291, -370.7875, 
    -371.6623, -371.3222, -373.1073, -372.3405, -374.3534, -373.8746, 
    -374.4683, -374.1655, -374.684, -374.2173, -375.0264, -375.2022, 
    -375.082, -375.545, -374.1914, -374.7107, -370.7834, -370.8064, 
    -370.9144, -370.4398, -370.4109, -369.9773, -370.3635, -370.5277, 
    -370.9461, -371.1927, -371.4272, -371.9429, -372.5167, -373.3177, 
    -373.9056, -374.2917, -374.0551, -374.2639, -374.0304, -373.9211, 
    -375.1361, -374.4535, -375.4784, -375.4218, -374.9576, -375.4282, 
    -370.8227, -370.6898, -370.2271, -370.5892, -369.9301, -370.2985, 
    -370.5101, -371.3286, -371.5091, -371.6753, -372.0045, -372.4255, 
    -373.1616, -373.8142, -374.4, -374.3572, -374.3722, -374.5027, -374.179, 
    -374.5559, -374.6189, -374.4538, -375.4142, -375.1398, -375.4206, 
    -375.242, -370.7331, -370.9569, -370.8359, -371.0633, -370.9028, 
    -371.6146, -371.8279, -372.824, -372.417, -373.0657, -372.4832, 
    -372.5862, -373.0854, -372.515, -373.7663, -372.9167, -374.5078, 
    -373.6456, -374.561, -374.3975, -374.6686, -374.9111, -375.2169, 
    -375.7801, -375.6498, -376.1215, -371.2907, -371.5803, -371.5555, 
    -371.8591, -372.0835, -372.5688, -373.345, -373.0533, -373.5894, 
    -373.6967, -372.8827, -373.382, -371.7747, -372.0347, -371.8804, 
    -371.3132, -373.1197, -372.1945, -373.915, -373.4023, -374.8764, 
    -374.1484, -375.5779, -376.1876, -376.7646, -377.4356, -371.7392, 
    -371.5423, -371.8954, -372.3819, -372.8335, -373.4327, -373.4943, 
    -373.6063, -373.9094, -374.1539, -373.6411, -374.2152, -372.0937, 
    -373.2003, -371.4672, -371.9898, -372.3535, -372.195, -373.0202, 
    -373.2144, -374.0149, -373.5956, -376.0366, -374.9614, -377.9488, 
    -377.1132, -371.4733, -371.7388, -372.6595, -372.2225, -373.473, 
    -373.7804, -374.0429, -374.3622, -374.3971, -374.5864, -374.2762, 
    -374.5744, -373.4339, -373.9502, -372.5553, -372.8915, -372.7371, 
    -372.5672, -373.0915, -373.6488, -373.6618, -373.8524, -374.3539, 
    -373.4781, -376.1734, -374.5139, -372.0283, -372.5365, -372.6102, 
    -372.4135, -373.7495, -373.2655, -374.5819, -374.2294, -374.8073, 
    -374.52, -374.4777, -374.1091, -373.8794, -373.2874, -372.8157, 
    -372.4422, -372.5291, -372.9395, -373.6832, -374.3998, -374.2453, 
    -374.7634, -373.3824, -373.9677, -373.7337, -374.3248, -373.0453, 
    -374.1334, -372.7699, -372.8886, -373.2559, -374.0058, -374.1708, 
    -374.345, -374.2377, -373.7023, -373.617, -373.2472, -373.1445, 
    -372.8629, -372.6292, -372.8424, -373.0661, -373.7029, -374.2885, 
    -374.9144, -375.068, -375.797, -375.2021, -376.1824, -375.3468, 
    -376.7947, -374.1973, -375.3243, -373.2729, -373.4927, -373.9012, 
    -374.8135, -374.3221, -374.8974, -373.6137, -372.9531, -372.7834, 
    -372.4647, -372.7907, -372.7642, -373.0761, -372.976, -373.7241, 
    -373.3224, -374.4764, -374.8931, -376.0717, -376.7938, -377.5309, 
    -377.8557, -377.9547, -377.9961 ;

 FGR12 =
  -167.3626, -167.416, -167.4057, -167.4488, -167.425, -167.4531, -167.3735, 
    -167.418, -167.3897, -167.3676, -167.5319, -167.4507, -167.6159, 
    -167.565, -167.695, -167.6079, -167.7125, -167.6928, -167.7529, 
    -167.7357, -167.8125, -167.7609, -167.853, -167.8003, -167.8084, 
    -167.7592, -167.4673, -167.5217, -167.464, -167.4718, -167.4683, 
    -167.4253, -167.4034, -167.3587, -167.3669, -167.3999, -167.4753, 
    -167.4499, -167.5145, -167.513, -167.5839, -167.5522, -167.6719, 
    -167.6369, -167.7364, -167.7115, -167.7352, -167.728, -167.7353, 
    -167.6989, -167.7144, -167.6825, -167.5581, -167.5941, -167.4853, 
    -167.4188, -167.3754, -167.3445, -167.3489, -167.3571, -167.4001, 
    -167.4408, -167.4717, -167.4924, -167.5128, -167.5732, -167.6054, 
    -167.6786, -167.6658, -167.6877, -167.7091, -167.7447, -167.7389, 
    -167.7545, -167.6873, -167.7319, -167.6573, -167.6784, -167.5174, 
    -167.4568, -167.4301, -167.4076, -167.3522, -167.3904, -167.3753, 
    -167.4114, -167.4343, -167.423, -167.4929, -167.4658, -167.6073, 
    -167.547, -167.7066, -167.6685, -167.7158, -167.6917, -167.733, 
    -167.6958, -167.7605, -167.7745, -167.7649, -167.8022, -167.6937, 
    -167.7351, -167.4227, -167.4245, -167.4332, -167.3951, -167.3929, 
    -167.3584, -167.3892, -167.4022, -167.4357, -167.4554, -167.4741, 
    -167.5154, -167.5609, -167.624, -167.6709, -167.7017, -167.6829, 
    -167.6995, -167.6809, -167.6722, -167.7692, -167.7145, -167.7968, 
    -167.7923, -167.7549, -167.7928, -167.4258, -167.4152, -167.3783, 
    -167.4072, -167.3547, -167.3839, -167.4007, -167.4661, -167.4807, 
    -167.4939, -167.5203, -167.5538, -167.6117, -167.6636, -167.7104, 
    -167.7069, -167.7081, -167.7185, -167.6927, -167.7228, -167.7278, 
    -167.7146, -167.7917, -167.7696, -167.7922, -167.7778, -167.4187, 
    -167.4366, -167.4269, -167.445, -167.4322, -167.4889, -167.506, -167.585, 
    -167.5531, -167.6041, -167.5584, -167.5664, -167.6054, -167.5609, 
    -167.6594, -167.5922, -167.7189, -167.6497, -167.7232, -167.7101, 
    -167.7318, -167.7512, -167.7758, -167.821, -167.8106, -167.8487, 
    -167.4632, -167.4863, -167.4844, -167.5087, -167.5266, -167.5651, 
    -167.6262, -167.6033, -167.6456, -167.6541, -167.5899, -167.6291, 
    -167.5018, -167.5225, -167.5103, -167.465, -167.6083, -167.5354, 
    -167.6716, -167.6308, -167.7484, -167.6901, -167.8048, -167.8538, 
    -167.901, -167.9555, -167.499, -167.4834, -167.5116, -167.5502, 
    -167.5859, -167.6331, -167.6381, -167.6469, -167.6713, -167.6907, 
    -167.6496, -167.6956, -167.527, -167.6147, -167.4773, -167.5189, 
    -167.548, -167.5355, -167.6007, -167.616, -167.6795, -167.6461, 
    -167.8415, -167.7551, -167.9978, -167.9292, -167.4778, -167.4991, 
    -167.5721, -167.5377, -167.6364, -167.6607, -167.6819, -167.7072, 
    -167.7101, -167.7252, -167.7005, -167.7243, -167.6332, -167.6745, 
    -167.5641, -167.5905, -167.5784, -167.565, -167.6063, -167.6501, 
    -167.6514, -167.6666, -167.7059, -167.6368, -167.8522, -167.7189, 
    -167.5223, -167.5623, -167.5684, -167.5529, -167.6583, -167.62, 
    -167.7248, -167.6967, -167.7429, -167.7199, -167.7165, -167.6871, 
    -167.6688, -167.6217, -167.5845, -167.5552, -167.562, -167.5942, 
    -167.6529, -167.7102, -167.6979, -167.7394, -167.6292, -167.6758, 
    -167.657, -167.7043, -167.6026, -167.6884, -167.581, -167.5903, 
    -167.6192, -167.6787, -167.6921, -167.7059, -167.6974, -167.6544, 
    -167.6477, -167.6186, -167.6104, -167.5883, -167.5699, -167.5867, 
    -167.6042, -167.6546, -167.7014, -167.7514, -167.7638, -167.8221, 
    -167.7743, -167.853, -167.7855, -167.9029, -167.6938, -167.784, 
    -167.6206, -167.638, -167.6704, -167.7431, -167.7041, -167.7499, 
    -167.6475, -167.5952, -167.582, -167.5569, -167.5826, -167.5806, 
    -167.6051, -167.5972, -167.6562, -167.6245, -167.7164, -167.7496, 
    -167.8446, -167.9032, -167.9636, -167.9903, -167.9984, -168.0018 ;

 FGR_R =
  -370.0307, -370.701, -370.571, -371.1112, -370.8119, -371.1653, -370.1671, 
    -370.7272, -370.3699, -370.0917, -372.1567, -371.1354, -373.2167, 
    -372.5682, -374.2104, -373.1152, -374.4292, -374.1802, -374.9322, 
    -374.7168, -375.6767, -375.0316, -376.1761, -375.5231, -375.6249, 
    -375.0101, -371.3419, -372.0292, -371.301, -371.399, -371.3553, 
    -370.8177, -370.546, -369.9803, -370.0832, -370.4991, -371.4431, 
    -371.1237, -371.931, -371.9128, -372.8076, -372.4049, -373.9185, -373.48, 
    -374.7258, -374.4153, -374.711, -374.6215, -374.7122, -374.2568, 
    -374.4518, -374.0515, -372.4802, -372.9382, -371.5678, -370.7393, 
    -370.1915, -369.802, -369.857, -369.9618, -370.5015, -371.01, -371.3968, 
    -371.6552, -371.9101, -372.6764, -373.0832, -374.0043, -373.841, 
    -374.1183, -374.3844, -374.8301, -374.7569, -374.9531, -374.1116, 
    -374.6705, -373.7359, -374, -371.9757, -371.21, -370.8811, -370.5959, 
    -369.8993, -370.3801, -370.1905, -370.6424, -370.9291, -370.7875, 
    -371.6623, -371.3222, -373.1073, -372.3405, -374.3534, -373.8746, 
    -374.4683, -374.1655, -374.684, -374.2173, -375.0264, -375.2022, 
    -375.082, -375.545, -374.1914, -374.7107, -370.7834, -370.8064, 
    -370.9144, -370.4398, -370.4109, -369.9773, -370.3635, -370.5277, 
    -370.9461, -371.1927, -371.4272, -371.9429, -372.5167, -373.3177, 
    -373.9056, -374.2917, -374.0551, -374.2639, -374.0304, -373.9211, 
    -375.1361, -374.4535, -375.4784, -375.4218, -374.9576, -375.4282, 
    -370.8227, -370.6898, -370.2271, -370.5892, -369.9301, -370.2985, 
    -370.5101, -371.3286, -371.5091, -371.6753, -372.0045, -372.4255, 
    -373.1616, -373.8142, -374.4, -374.3572, -374.3722, -374.5027, -374.179, 
    -374.5559, -374.6189, -374.4538, -375.4142, -375.1398, -375.4206, 
    -375.242, -370.7331, -370.9569, -370.8359, -371.0633, -370.9028, 
    -371.6146, -371.8279, -372.824, -372.417, -373.0657, -372.4832, 
    -372.5862, -373.0854, -372.515, -373.7663, -372.9167, -374.5078, 
    -373.6456, -374.561, -374.3975, -374.6686, -374.9111, -375.2169, 
    -375.7801, -375.6498, -376.1215, -371.2907, -371.5803, -371.5555, 
    -371.8591, -372.0835, -372.5688, -373.345, -373.0533, -373.5894, 
    -373.6967, -372.8827, -373.382, -371.7747, -372.0347, -371.8804, 
    -371.3132, -373.1197, -372.1945, -373.915, -373.4023, -374.8764, 
    -374.1484, -375.5779, -376.1876, -376.7646, -377.4356, -371.7392, 
    -371.5423, -371.8954, -372.3819, -372.8335, -373.4327, -373.4943, 
    -373.6063, -373.9094, -374.1539, -373.6411, -374.2152, -372.0937, 
    -373.2003, -371.4672, -371.9898, -372.3535, -372.195, -373.0202, 
    -373.2144, -374.0149, -373.5956, -376.0366, -374.9614, -377.9488, 
    -377.1132, -371.4733, -371.7388, -372.6595, -372.2225, -373.473, 
    -373.7804, -374.0429, -374.3622, -374.3971, -374.5864, -374.2762, 
    -374.5744, -373.4339, -373.9502, -372.5553, -372.8915, -372.7371, 
    -372.5672, -373.0915, -373.6488, -373.6618, -373.8524, -374.3539, 
    -373.4781, -376.1734, -374.5139, -372.0283, -372.5365, -372.6102, 
    -372.4135, -373.7495, -373.2655, -374.5819, -374.2294, -374.8073, 
    -374.52, -374.4777, -374.1091, -373.8794, -373.2874, -372.8157, 
    -372.4422, -372.5291, -372.9395, -373.6832, -374.3998, -374.2453, 
    -374.7634, -373.3824, -373.9677, -373.7337, -374.3248, -373.0453, 
    -374.1334, -372.7699, -372.8886, -373.2559, -374.0058, -374.1708, 
    -374.345, -374.2377, -373.7023, -373.617, -373.2472, -373.1445, 
    -372.8629, -372.6292, -372.8424, -373.0661, -373.7029, -374.2885, 
    -374.9144, -375.068, -375.797, -375.2021, -376.1824, -375.3468, 
    -376.7947, -374.1973, -375.3243, -373.2729, -373.4927, -373.9012, 
    -374.8135, -374.3221, -374.8974, -373.6137, -372.9531, -372.7834, 
    -372.4647, -372.7907, -372.7642, -373.0761, -372.976, -373.7241, 
    -373.3224, -374.4764, -374.8931, -376.0717, -376.7938, -377.5309, 
    -377.8557, -377.9547, -377.9961 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  77.91566, 77.96246, 77.95338, 77.99108, 77.9702, 77.99487, 77.92519, 
    77.96429, 77.93935, 77.91993, 78.06425, 77.99277, 78.13919, 78.09333, 
    78.20826, 78.132, 78.22375, 78.20614, 78.25935, 78.24411, 78.312, 
    78.26639, 78.34733, 78.30115, 78.30834, 78.26487, 78.00724, 78.05532, 
    78.00437, 78.01123, 78.00817, 77.9706, 77.95163, 77.91215, 77.91933, 
    77.94836, 78.01432, 77.99196, 78.04848, 78.0472, 78.11027, 78.08179, 
    78.18761, 78.15786, 78.24475, 78.22277, 78.24371, 78.23737, 78.24378, 
    78.21156, 78.22536, 78.19703, 78.0871, 78.1195, 78.02305, 77.96513, 
    77.92689, 77.8997, 77.90354, 77.91085, 77.94853, 77.98402, 78.01108, 
    78.02917, 78.04702, 78.10095, 78.12975, 78.19367, 78.18213, 78.20174, 
    78.22059, 78.25213, 78.24695, 78.26083, 78.20128, 78.24083, 78.17599, 
    78.19338, 78.05158, 77.99801, 77.97501, 77.95512, 77.90649, 77.94006, 
    77.92682, 77.95837, 77.97839, 77.9685, 78.02967, 78.00586, 78.13145, 
    78.07723, 78.21839, 78.1845, 78.22652, 78.20509, 78.24179, 78.20877, 
    78.26601, 78.27845, 78.26994, 78.3027, 78.20693, 78.24368, 77.96821, 
    77.96982, 77.97736, 77.94422, 77.94221, 77.91193, 77.9389, 77.95036, 
    77.97957, 77.9968, 78.01321, 78.04931, 78.08968, 78.14635, 78.1867, 
    78.21403, 78.19729, 78.21207, 78.19553, 78.1878, 78.27377, 78.22547, 
    78.29799, 78.29399, 78.26115, 78.29444, 77.97095, 77.96168, 77.92938, 
    77.95466, 77.90865, 77.93436, 77.94913, 78.00629, 78.01894, 78.03058, 
    78.05363, 78.08324, 78.1353, 78.18023, 78.22169, 78.21867, 78.21973, 
    78.22897, 78.20605, 78.23273, 78.23717, 78.2255, 78.29345, 78.27404, 
    78.29391, 78.28127, 77.9647, 77.98032, 77.97188, 77.98774, 77.97654, 
    78.02632, 78.04125, 78.11141, 78.08264, 78.12852, 78.08733, 78.0946, 
    78.12988, 78.08957, 78.17812, 78.11796, 78.22932, 78.16956, 78.23309, 
    78.22152, 78.24071, 78.25786, 78.2795, 78.31933, 78.31011, 78.34348, 
    78.00365, 78.02393, 78.02219, 78.04345, 78.05915, 78.09338, 78.14828, 
    78.12766, 78.16561, 78.17321, 78.11559, 78.1509, 78.03754, 78.05573, 
    78.04494, 78.00523, 78.13233, 78.06693, 78.18736, 78.15235, 78.25541, 
    78.20387, 78.30503, 78.34813, 78.38895, 78.43636, 78.03505, 78.02127, 
    78.04599, 78.08015, 78.1121, 78.1545, 78.15887, 78.16681, 78.18697, 
    78.20428, 78.16926, 78.20862, 78.05984, 78.13804, 78.01601, 78.05258, 
    78.07816, 78.06697, 78.12531, 78.13905, 78.19443, 78.16605, 78.33744, 
    78.26141, 78.47263, 78.41357, 78.01644, 78.03503, 78.09978, 78.06892, 
    78.15736, 78.17913, 78.19642, 78.21901, 78.22149, 78.23488, 78.21293, 
    78.23404, 78.15459, 78.18985, 78.09243, 78.1162, 78.10529, 78.09327, 
    78.13036, 78.16981, 78.17074, 78.18292, 78.21837, 78.15772, 78.34709, 
    78.22971, 78.05528, 78.09107, 78.09631, 78.0824, 78.17695, 78.14265, 
    78.23457, 78.20963, 78.25052, 78.23019, 78.2272, 78.2011, 78.18484, 
    78.14421, 78.11084, 78.08443, 78.09058, 78.11959, 78.17224, 78.22167, 
    78.21073, 78.24741, 78.15094, 78.19109, 78.17582, 78.21637, 78.12708, 
    78.20277, 78.1076, 78.116, 78.14198, 78.19378, 78.20547, 78.2178, 
    78.21021, 78.17359, 78.16756, 78.14137, 78.13409, 78.11418, 78.09766, 
    78.11273, 78.12855, 78.17365, 78.21379, 78.25809, 78.26897, 78.3205, 
    78.27842, 78.34772, 78.28862, 78.39103, 78.20732, 78.28706, 78.14319, 
    78.15876, 78.18637, 78.25094, 78.21618, 78.25687, 78.16734, 78.12054, 
    78.10857, 78.08601, 78.10908, 78.10721, 78.12927, 78.12218, 78.17515, 
    78.14669, 78.2271, 78.25658, 78.33994, 78.391, 78.44311, 78.46606, 
    78.47306, 78.47598 ;

 FIRA_R =
  77.91566, 77.96246, 77.95338, 77.99108, 77.9702, 77.99487, 77.92519, 
    77.96429, 77.93935, 77.91993, 78.06425, 77.99277, 78.13919, 78.09333, 
    78.20826, 78.132, 78.22375, 78.20614, 78.25935, 78.24411, 78.312, 
    78.26639, 78.34733, 78.30115, 78.30834, 78.26487, 78.00724, 78.05532, 
    78.00437, 78.01123, 78.00817, 77.9706, 77.95163, 77.91215, 77.91933, 
    77.94836, 78.01432, 77.99196, 78.04848, 78.0472, 78.11027, 78.08179, 
    78.18761, 78.15786, 78.24475, 78.22277, 78.24371, 78.23737, 78.24378, 
    78.21156, 78.22536, 78.19703, 78.0871, 78.1195, 78.02305, 77.96513, 
    77.92689, 77.8997, 77.90354, 77.91085, 77.94853, 77.98402, 78.01108, 
    78.02917, 78.04702, 78.10095, 78.12975, 78.19367, 78.18213, 78.20174, 
    78.22059, 78.25213, 78.24695, 78.26083, 78.20128, 78.24083, 78.17599, 
    78.19338, 78.05158, 77.99801, 77.97501, 77.95512, 77.90649, 77.94006, 
    77.92682, 77.95837, 77.97839, 77.9685, 78.02967, 78.00586, 78.13145, 
    78.07723, 78.21839, 78.1845, 78.22652, 78.20509, 78.24179, 78.20877, 
    78.26601, 78.27845, 78.26994, 78.3027, 78.20693, 78.24368, 77.96821, 
    77.96982, 77.97736, 77.94422, 77.94221, 77.91193, 77.9389, 77.95036, 
    77.97957, 77.9968, 78.01321, 78.04931, 78.08968, 78.14635, 78.1867, 
    78.21403, 78.19729, 78.21207, 78.19553, 78.1878, 78.27377, 78.22547, 
    78.29799, 78.29399, 78.26115, 78.29444, 77.97095, 77.96168, 77.92938, 
    77.95466, 77.90865, 77.93436, 77.94913, 78.00629, 78.01894, 78.03058, 
    78.05363, 78.08324, 78.1353, 78.18023, 78.22169, 78.21867, 78.21973, 
    78.22897, 78.20605, 78.23273, 78.23717, 78.2255, 78.29345, 78.27404, 
    78.29391, 78.28127, 77.9647, 77.98032, 77.97188, 77.98774, 77.97654, 
    78.02632, 78.04125, 78.11141, 78.08264, 78.12852, 78.08733, 78.0946, 
    78.12988, 78.08957, 78.17812, 78.11796, 78.22932, 78.16956, 78.23309, 
    78.22152, 78.24071, 78.25786, 78.2795, 78.31933, 78.31011, 78.34348, 
    78.00365, 78.02393, 78.02219, 78.04345, 78.05915, 78.09338, 78.14828, 
    78.12766, 78.16561, 78.17321, 78.11559, 78.1509, 78.03754, 78.05573, 
    78.04494, 78.00523, 78.13233, 78.06693, 78.18736, 78.15235, 78.25541, 
    78.20387, 78.30503, 78.34813, 78.38895, 78.43636, 78.03505, 78.02127, 
    78.04599, 78.08015, 78.1121, 78.1545, 78.15887, 78.16681, 78.18697, 
    78.20428, 78.16926, 78.20862, 78.05984, 78.13804, 78.01601, 78.05258, 
    78.07816, 78.06697, 78.12531, 78.13905, 78.19443, 78.16605, 78.33744, 
    78.26141, 78.47263, 78.41357, 78.01644, 78.03503, 78.09978, 78.06892, 
    78.15736, 78.17913, 78.19642, 78.21901, 78.22149, 78.23488, 78.21293, 
    78.23404, 78.15459, 78.18985, 78.09243, 78.1162, 78.10529, 78.09327, 
    78.13036, 78.16981, 78.17074, 78.18292, 78.21837, 78.15772, 78.34709, 
    78.22971, 78.05528, 78.09107, 78.09631, 78.0824, 78.17695, 78.14265, 
    78.23457, 78.20963, 78.25052, 78.23019, 78.2272, 78.2011, 78.18484, 
    78.14421, 78.11084, 78.08443, 78.09058, 78.11959, 78.17224, 78.22167, 
    78.21073, 78.24741, 78.15094, 78.19109, 78.17582, 78.21637, 78.12708, 
    78.20277, 78.1076, 78.116, 78.14198, 78.19378, 78.20547, 78.2178, 
    78.21021, 78.17359, 78.16756, 78.14137, 78.13409, 78.11418, 78.09766, 
    78.11273, 78.12855, 78.17365, 78.21379, 78.25809, 78.26897, 78.3205, 
    78.27842, 78.34772, 78.28862, 78.39103, 78.20732, 78.28706, 78.14319, 
    78.15876, 78.18637, 78.25094, 78.21618, 78.25687, 78.16734, 78.12054, 
    78.10857, 78.08601, 78.10908, 78.10721, 78.12927, 78.12218, 78.17515, 
    78.14669, 78.2271, 78.25658, 78.33994, 78.391, 78.44311, 78.46606, 
    78.47306, 78.47598 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  266.8766, 266.9234, 266.9143, 266.952, 266.9312, 266.9558, 266.8861, 
    266.9252, 266.9003, 266.8809, 267.0252, 266.9537, 267.1001, 267.0543, 
    267.1692, 267.093, 267.1847, 267.1671, 267.2203, 267.205, 267.2729, 
    267.2273, 267.3083, 267.2621, 267.2693, 267.2258, 266.9682, 267.0163, 
    266.9653, 266.9722, 266.9691, 266.9315, 266.9126, 266.8731, 266.8803, 
    266.9093, 266.9753, 266.9529, 267.0094, 267.0081, 267.0712, 267.0427, 
    267.1486, 267.1188, 267.2057, 267.1837, 267.2047, 267.1983, 267.2047, 
    267.1725, 267.1863, 267.158, 267.048, 267.0804, 266.984, 266.9261, 
    266.8878, 266.8606, 266.8645, 266.8718, 266.9095, 266.945, 266.972, 
    266.9901, 267.008, 267.0619, 267.0907, 267.1546, 267.1431, 267.1627, 
    267.1815, 267.2131, 267.2079, 267.2218, 267.1622, 267.2018, 267.1369, 
    267.1543, 267.0125, 266.959, 266.9359, 266.916, 266.8674, 266.901, 
    266.8878, 266.9193, 266.9393, 266.9294, 266.9906, 266.9668, 267.0924, 
    267.0382, 267.1793, 267.1454, 267.1875, 267.166, 267.2027, 267.1697, 
    267.227, 267.2394, 267.2309, 267.2636, 267.1679, 267.2046, 266.9291, 
    266.9308, 266.9383, 266.9052, 266.9031, 266.8729, 266.8998, 266.9113, 
    266.9405, 266.9577, 266.9742, 267.0103, 267.0506, 267.1073, 267.1476, 
    267.175, 267.1582, 267.173, 267.1565, 267.1487, 267.2347, 267.1864, 
    267.2589, 267.2549, 267.2221, 267.2554, 266.9319, 266.9226, 266.8903, 
    266.9156, 266.8696, 266.8953, 266.9101, 266.9672, 266.9799, 266.9915, 
    267.0146, 267.0442, 267.0963, 267.1412, 267.1826, 267.1796, 267.1807, 
    267.1899, 267.167, 267.1937, 267.1981, 267.1864, 267.2544, 267.235, 
    267.2549, 267.2422, 266.9256, 266.9413, 266.9328, 266.9487, 266.9375, 
    266.9873, 267.0022, 267.0724, 267.0436, 267.0894, 267.0482, 267.0555, 
    267.0908, 267.0505, 267.1391, 267.0789, 267.1902, 267.1305, 267.194, 
    267.1825, 267.2017, 267.2188, 267.2404, 267.2803, 267.2711, 267.3044, 
    266.9646, 266.9849, 266.9831, 267.0044, 267.0201, 267.0543, 267.1092, 
    267.0886, 267.1266, 267.1342, 267.0765, 267.1118, 266.9985, 267.0167, 
    267.0059, 266.9662, 267.0933, 267.0279, 267.1483, 267.1133, 267.2163, 
    267.1648, 267.266, 267.3091, 267.3499, 267.3973, 266.996, 266.9822, 
    267.0069, 267.0411, 267.073, 267.1154, 267.1198, 267.1277, 267.1479, 
    267.1652, 267.1302, 267.1696, 267.0208, 267.099, 266.977, 267.0135, 
    267.0391, 267.0279, 267.0862, 267.1, 267.1554, 267.127, 267.2984, 
    267.2224, 267.4336, 267.3745, 266.9774, 266.996, 267.0607, 267.0298, 
    267.1183, 267.1401, 267.1573, 267.18, 267.1824, 267.1958, 267.1739, 
    267.195, 267.1155, 267.1508, 267.0534, 267.0771, 267.0662, 267.0542, 
    267.0913, 267.1307, 267.1317, 267.1439, 267.1793, 267.1187, 267.308, 
    267.1906, 267.0162, 267.052, 267.0573, 267.0433, 267.1379, 267.1036, 
    267.1955, 267.1706, 267.2115, 267.1911, 267.1881, 267.162, 267.1458, 
    267.1052, 267.0718, 267.0453, 267.0515, 267.0805, 267.1332, 267.1826, 
    267.1717, 267.2083, 267.1119, 267.152, 267.1367, 267.1773, 267.088, 
    267.1637, 267.0685, 267.0769, 267.1029, 267.1547, 267.1664, 267.1787, 
    267.1711, 267.1345, 267.1285, 267.1023, 267.095, 267.0751, 267.0586, 
    267.0737, 267.0895, 267.1346, 267.1747, 267.219, 267.2299, 267.2814, 
    267.2393, 267.3087, 267.2495, 267.352, 267.1682, 267.248, 267.1041, 
    267.1197, 267.1473, 267.2119, 267.1771, 267.2178, 267.1283, 267.0815, 
    267.0695, 267.0469, 267.07, 267.0681, 267.0902, 267.0831, 267.1361, 
    267.1076, 267.188, 267.2175, 267.3009, 267.3519, 267.4041, 267.427, 
    267.434, 267.4369 ;

 FIRE_R =
  266.8766, 266.9234, 266.9143, 266.952, 266.9312, 266.9558, 266.8861, 
    266.9252, 266.9003, 266.8809, 267.0252, 266.9537, 267.1001, 267.0543, 
    267.1692, 267.093, 267.1847, 267.1671, 267.2203, 267.205, 267.2729, 
    267.2273, 267.3083, 267.2621, 267.2693, 267.2258, 266.9682, 267.0163, 
    266.9653, 266.9722, 266.9691, 266.9315, 266.9126, 266.8731, 266.8803, 
    266.9093, 266.9753, 266.9529, 267.0094, 267.0081, 267.0712, 267.0427, 
    267.1486, 267.1188, 267.2057, 267.1837, 267.2047, 267.1983, 267.2047, 
    267.1725, 267.1863, 267.158, 267.048, 267.0804, 266.984, 266.9261, 
    266.8878, 266.8606, 266.8645, 266.8718, 266.9095, 266.945, 266.972, 
    266.9901, 267.008, 267.0619, 267.0907, 267.1546, 267.1431, 267.1627, 
    267.1815, 267.2131, 267.2079, 267.2218, 267.1622, 267.2018, 267.1369, 
    267.1543, 267.0125, 266.959, 266.9359, 266.916, 266.8674, 266.901, 
    266.8878, 266.9193, 266.9393, 266.9294, 266.9906, 266.9668, 267.0924, 
    267.0382, 267.1793, 267.1454, 267.1875, 267.166, 267.2027, 267.1697, 
    267.227, 267.2394, 267.2309, 267.2636, 267.1679, 267.2046, 266.9291, 
    266.9308, 266.9383, 266.9052, 266.9031, 266.8729, 266.8998, 266.9113, 
    266.9405, 266.9577, 266.9742, 267.0103, 267.0506, 267.1073, 267.1476, 
    267.175, 267.1582, 267.173, 267.1565, 267.1487, 267.2347, 267.1864, 
    267.2589, 267.2549, 267.2221, 267.2554, 266.9319, 266.9226, 266.8903, 
    266.9156, 266.8696, 266.8953, 266.9101, 266.9672, 266.9799, 266.9915, 
    267.0146, 267.0442, 267.0963, 267.1412, 267.1826, 267.1796, 267.1807, 
    267.1899, 267.167, 267.1937, 267.1981, 267.1864, 267.2544, 267.235, 
    267.2549, 267.2422, 266.9256, 266.9413, 266.9328, 266.9487, 266.9375, 
    266.9873, 267.0022, 267.0724, 267.0436, 267.0894, 267.0482, 267.0555, 
    267.0908, 267.0505, 267.1391, 267.0789, 267.1902, 267.1305, 267.194, 
    267.1825, 267.2017, 267.2188, 267.2404, 267.2803, 267.2711, 267.3044, 
    266.9646, 266.9849, 266.9831, 267.0044, 267.0201, 267.0543, 267.1092, 
    267.0886, 267.1266, 267.1342, 267.0765, 267.1118, 266.9985, 267.0167, 
    267.0059, 266.9662, 267.0933, 267.0279, 267.1483, 267.1133, 267.2163, 
    267.1648, 267.266, 267.3091, 267.3499, 267.3973, 266.996, 266.9822, 
    267.0069, 267.0411, 267.073, 267.1154, 267.1198, 267.1277, 267.1479, 
    267.1652, 267.1302, 267.1696, 267.0208, 267.099, 266.977, 267.0135, 
    267.0391, 267.0279, 267.0862, 267.1, 267.1554, 267.127, 267.2984, 
    267.2224, 267.4336, 267.3745, 266.9774, 266.996, 267.0607, 267.0298, 
    267.1183, 267.1401, 267.1573, 267.18, 267.1824, 267.1958, 267.1739, 
    267.195, 267.1155, 267.1508, 267.0534, 267.0771, 267.0662, 267.0542, 
    267.0913, 267.1307, 267.1317, 267.1439, 267.1793, 267.1187, 267.308, 
    267.1906, 267.0162, 267.052, 267.0573, 267.0433, 267.1379, 267.1036, 
    267.1955, 267.1706, 267.2115, 267.1911, 267.1881, 267.162, 267.1458, 
    267.1052, 267.0718, 267.0453, 267.0515, 267.0805, 267.1332, 267.1826, 
    267.1717, 267.2083, 267.1119, 267.152, 267.1367, 267.1773, 267.088, 
    267.1637, 267.0685, 267.0769, 267.1029, 267.1547, 267.1664, 267.1787, 
    267.1711, 267.1345, 267.1285, 267.1023, 267.095, 267.0751, 267.0586, 
    267.0737, 267.0895, 267.1346, 267.1747, 267.219, 267.2299, 267.2814, 
    267.2393, 267.3087, 267.2495, 267.352, 267.1682, 267.248, 267.1041, 
    267.1197, 267.1473, 267.2119, 267.1771, 267.2178, 267.1283, 267.0815, 
    267.0695, 267.0469, 267.07, 267.0681, 267.0902, 267.0831, 267.1361, 
    267.1076, 267.188, 267.2175, 267.3009, 267.3519, 267.4041, 267.427, 
    267.434, 267.4369 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  286.2084, 286.813, 286.6957, 287.183, 286.913, 287.2318, 286.3314, 
    286.8367, 286.5143, 286.2634, 288.1261, 287.2048, 289.0811, 288.4968, 
    289.9763, 288.9897, 290.1733, 289.949, 290.6263, 290.4323, 291.2972, 
    290.7159, 291.747, 291.1588, 291.2505, 290.6966, 287.3911, 288.011, 
    287.3541, 287.4426, 287.4031, 286.9183, 286.6732, 286.1629, 286.2557, 
    286.6308, 287.4824, 287.1942, 287.9223, 287.9059, 288.7125, 288.3496, 
    289.7132, 289.3182, 290.4404, 290.1607, 290.4272, 290.3465, 290.4282, 
    290.018, 290.1937, 289.833, 288.4174, 288.8301, 287.5948, 286.8476, 
    286.3534, 286.002, 286.0517, 286.1462, 286.633, 287.0917, 287.4405, 
    287.6736, 287.9035, 288.5943, 288.9608, 289.7905, 289.6434, 289.8932, 
    290.1329, 290.5345, 290.4684, 290.6452, 289.8871, 290.3907, 289.5487, 
    289.7866, 287.9628, 287.2721, 286.9755, 286.7181, 286.0898, 286.5235, 
    286.3525, 286.7601, 287.0188, 286.891, 287.68, 287.3733, 288.9826, 
    288.2916, 290.1049, 289.6736, 290.2084, 289.9356, 290.4028, 289.9824, 
    290.7112, 290.8697, 290.7614, 291.1784, 289.959, 290.4269, 286.8872, 
    286.9081, 287.0054, 286.5774, 286.5514, 286.1602, 286.5085, 286.6567, 
    287.034, 287.2565, 287.468, 287.9331, 288.4504, 289.1721, 289.7015, 
    290.0493, 289.8363, 290.0244, 289.814, 289.7155, 290.8101, 290.1951, 
    291.1184, 291.0674, 290.6493, 291.0732, 286.9227, 286.8028, 286.3855, 
    286.7121, 286.1176, 286.45, 286.6408, 287.379, 287.5418, 287.6917, 
    287.9887, 288.3682, 289.0314, 289.6193, 290.147, 290.1083, 290.1219, 
    290.2395, 289.9478, 290.2874, 290.3441, 290.1954, 291.0606, 290.8134, 
    291.0663, 290.9055, 286.8419, 287.0438, 286.9346, 287.1398, 286.995, 
    287.637, 287.8295, 288.7273, 288.3605, 288.945, 288.4202, 288.513, 
    288.9629, 288.4487, 289.5762, 288.8108, 290.2441, 289.4676, 290.292, 
    290.1447, 290.3889, 290.6074, 290.8828, 291.3903, 291.2729, 291.6978, 
    287.3449, 287.6061, 287.5837, 287.8575, 288.0599, 288.4973, 289.1966, 
    288.9338, 289.4167, 289.5135, 288.7801, 289.2299, 287.7814, 288.016, 
    287.8767, 287.3651, 288.9937, 288.16, 289.71, 289.2482, 290.5762, 
    289.9203, 291.2081, 291.7575, 292.2773, 292.8818, 287.7493, 287.5717, 
    287.8903, 288.3289, 288.7358, 289.2756, 289.3311, 289.432, 289.705, 
    289.9252, 289.4634, 289.9805, 288.0692, 289.0663, 287.5041, 287.9754, 
    288.3033, 288.1604, 288.904, 289.0789, 289.8001, 289.4223, 291.6214, 
    290.6528, 293.3441, 292.5913, 287.5096, 287.749, 288.579, 288.1852, 
    289.3119, 289.5888, 289.8252, 290.1129, 290.1443, 290.3149, 290.0354, 
    290.304, 289.2768, 289.7417, 288.4851, 288.7881, 288.6489, 288.4958, 
    288.9682, 289.4704, 289.482, 289.6536, 290.1056, 289.3165, 291.7448, 
    290.2498, 288.0101, 288.4682, 288.5346, 288.3573, 289.561, 289.125, 
    290.3109, 289.9933, 290.5139, 290.2551, 290.217, 289.8849, 289.6779, 
    289.1448, 288.7198, 288.3832, 288.4615, 288.8313, 289.5013, 290.1468, 
    290.0076, 290.4743, 289.2303, 289.7575, 289.5468, 290.0792, 288.9267, 
    289.9069, 288.6784, 288.7854, 289.1163, 289.7919, 289.9404, 290.0974, 
    290.0007, 289.5185, 289.4417, 289.1085, 289.016, 288.7622, 288.5517, 
    288.7438, 288.9454, 289.5191, 290.0465, 290.6104, 290.7487, 291.4057, 
    290.8697, 291.753, 291.0002, 292.3045, 289.9644, 290.9798, 289.1317, 
    289.3297, 289.6977, 290.5196, 290.0767, 290.5951, 289.4387, 288.8436, 
    288.6906, 288.4035, 288.6972, 288.6733, 288.9544, 288.8641, 289.5381, 
    289.1762, 290.2158, 290.5912, 291.653, 292.3036, 292.9675, 293.2602, 
    293.3494, 293.3866 ;

 FSH_G =
  299.3114, 299.9171, 299.7995, 300.2876, 300.0172, 300.3365, 299.4346, 
    299.9407, 299.6179, 299.3665, 301.2322, 300.3095, 302.1889, 301.6035, 
    303.0854, 302.0973, 303.2828, 303.0581, 303.7366, 303.5423, 304.4085, 
    303.8263, 304.8591, 304.2699, 304.3618, 303.807, 300.496, 301.117, 
    300.459, 300.5476, 300.5081, 300.0225, 299.7769, 299.2658, 299.3588, 
    299.7346, 300.5875, 300.2989, 301.0282, 301.0117, 301.8196, 301.4561, 
    302.8219, 302.4264, 303.5504, 303.2702, 303.5371, 303.4563, 303.5381, 
    303.1272, 303.3032, 302.942, 301.5241, 301.9374, 300.7001, 299.9517, 
    299.4567, 299.1047, 299.1545, 299.2491, 299.7367, 300.1961, 300.5456, 
    300.7791, 301.0093, 301.7012, 302.0684, 302.8994, 302.752, 303.0022, 
    303.2423, 303.6445, 303.5785, 303.7555, 302.9962, 303.5005, 302.6573, 
    302.8955, 301.0687, 300.3769, 300.0797, 299.822, 299.1927, 299.6271, 
    299.4557, 299.8641, 300.1231, 299.9951, 300.7855, 300.4782, 302.0901, 
    301.398, 303.2143, 302.7823, 303.318, 303.0448, 303.5127, 303.0916, 
    303.8216, 303.9803, 303.8718, 304.2896, 303.0681, 303.5368, 299.9914, 
    300.0122, 300.1098, 299.681, 299.655, 299.2631, 299.6121, 299.7604, 
    300.1384, 300.3613, 300.5731, 301.039, 301.5571, 302.28, 302.8103, 
    303.1586, 302.9452, 303.1336, 302.9229, 302.8243, 303.9207, 303.3047, 
    304.2295, 304.1784, 303.7596, 304.1842, 300.0269, 299.9068, 299.4888, 
    299.8159, 299.2205, 299.5533, 299.7445, 300.484, 300.647, 300.7972, 
    301.0946, 301.4747, 302.1391, 302.7279, 303.2564, 303.2177, 303.2314, 
    303.3491, 303.057, 303.3971, 303.4539, 303.305, 304.1716, 303.924, 
    304.1773, 304.0162, 299.946, 300.1482, 300.0389, 300.2443, 300.0993, 
    300.7424, 300.9352, 301.8344, 301.4671, 302.0526, 301.5269, 301.6198, 
    302.0704, 301.5555, 302.6848, 301.9181, 303.3537, 302.5759, 303.4017, 
    303.2542, 303.4988, 303.7176, 303.9935, 304.5018, 304.3842, 304.8098, 
    300.4498, 300.7114, 300.689, 300.9633, 301.166, 301.6041, 302.3046, 
    302.0414, 302.5251, 302.6219, 301.8874, 302.3379, 300.887, 301.1219, 
    300.9825, 300.4701, 302.1013, 301.2662, 302.8188, 302.3562, 303.6863, 
    303.0294, 304.3193, 304.8696, 305.3902, 305.9958, 300.8549, 300.677, 
    300.9961, 301.4354, 301.843, 302.3837, 302.4393, 302.5404, 302.8137, 
    303.0343, 302.5718, 303.0897, 301.1752, 302.174, 300.6092, 301.0813, 
    301.4098, 301.2667, 302.0114, 302.1867, 302.909, 302.5306, 304.7333, 
    303.7631, 306.4588, 305.7047, 300.6147, 300.8546, 301.6859, 301.2915, 
    302.42, 302.6974, 302.9342, 303.2223, 303.2538, 303.4246, 303.1447, 
    303.4138, 302.3848, 302.8505, 301.5919, 301.8954, 301.756, 301.6026, 
    302.0758, 302.5788, 302.5904, 302.7623, 303.2149, 302.4247, 304.8569, 
    303.3594, 301.1161, 301.575, 301.6414, 301.4639, 302.6696, 302.2328, 
    303.4206, 303.1025, 303.6239, 303.3647, 303.3265, 302.9939, 302.7866, 
    302.2527, 301.8269, 301.4898, 301.5683, 301.9386, 302.6097, 303.2563, 
    303.1168, 303.5843, 302.3383, 302.8663, 302.6553, 303.1885, 302.0342, 
    303.016, 301.7856, 301.8927, 302.2242, 302.9008, 303.0496, 303.2068, 
    303.11, 302.627, 302.55, 302.2163, 302.1236, 301.8694, 301.6586, 301.851, 
    302.0529, 302.6275, 303.1558, 303.7206, 303.8592, 304.5172, 303.9803, 
    304.865, 304.1109, 305.4174, 303.0736, 304.0906, 302.2395, 302.4378, 
    302.8064, 303.6296, 303.1861, 303.7053, 302.5471, 301.9509, 301.7978, 
    301.5101, 301.8043, 301.7804, 302.0619, 301.9715, 302.6466, 302.2841, 
    303.3253, 303.7014, 304.7649, 305.4166, 306.0816, 306.3748, 306.4641, 
    306.5014 ;

 FSH_NODYNLNDUSE =
  286.2084, 286.813, 286.6957, 287.183, 286.913, 287.2318, 286.3314, 
    286.8367, 286.5143, 286.2634, 288.1261, 287.2048, 289.0811, 288.4968, 
    289.9763, 288.9897, 290.1733, 289.949, 290.6263, 290.4323, 291.2972, 
    290.7159, 291.747, 291.1588, 291.2505, 290.6966, 287.3911, 288.011, 
    287.3541, 287.4426, 287.4031, 286.9183, 286.6732, 286.1629, 286.2557, 
    286.6308, 287.4824, 287.1942, 287.9223, 287.9059, 288.7125, 288.3496, 
    289.7132, 289.3182, 290.4404, 290.1607, 290.4272, 290.3465, 290.4282, 
    290.018, 290.1937, 289.833, 288.4174, 288.8301, 287.5948, 286.8476, 
    286.3534, 286.002, 286.0517, 286.1462, 286.633, 287.0917, 287.4405, 
    287.6736, 287.9035, 288.5943, 288.9608, 289.7905, 289.6434, 289.8932, 
    290.1329, 290.5345, 290.4684, 290.6452, 289.8871, 290.3907, 289.5487, 
    289.7866, 287.9628, 287.2721, 286.9755, 286.7181, 286.0898, 286.5235, 
    286.3525, 286.7601, 287.0188, 286.891, 287.68, 287.3733, 288.9826, 
    288.2916, 290.1049, 289.6736, 290.2084, 289.9356, 290.4028, 289.9824, 
    290.7112, 290.8697, 290.7614, 291.1784, 289.959, 290.4269, 286.8872, 
    286.9081, 287.0054, 286.5774, 286.5514, 286.1602, 286.5085, 286.6567, 
    287.034, 287.2565, 287.468, 287.9331, 288.4504, 289.1721, 289.7015, 
    290.0493, 289.8363, 290.0244, 289.814, 289.7155, 290.8101, 290.1951, 
    291.1184, 291.0674, 290.6493, 291.0732, 286.9227, 286.8028, 286.3855, 
    286.7121, 286.1176, 286.45, 286.6408, 287.379, 287.5418, 287.6917, 
    287.9887, 288.3682, 289.0314, 289.6193, 290.147, 290.1083, 290.1219, 
    290.2395, 289.9478, 290.2874, 290.3441, 290.1954, 291.0606, 290.8134, 
    291.0663, 290.9055, 286.8419, 287.0438, 286.9346, 287.1398, 286.995, 
    287.637, 287.8295, 288.7273, 288.3605, 288.945, 288.4202, 288.513, 
    288.9629, 288.4487, 289.5762, 288.8108, 290.2441, 289.4676, 290.292, 
    290.1447, 290.3889, 290.6074, 290.8828, 291.3903, 291.2729, 291.6978, 
    287.3449, 287.6061, 287.5837, 287.8575, 288.0599, 288.4973, 289.1966, 
    288.9338, 289.4167, 289.5135, 288.7801, 289.2299, 287.7814, 288.016, 
    287.8767, 287.3651, 288.9937, 288.16, 289.71, 289.2482, 290.5762, 
    289.9203, 291.2081, 291.7575, 292.2773, 292.8818, 287.7493, 287.5717, 
    287.8903, 288.3289, 288.7358, 289.2756, 289.3311, 289.432, 289.705, 
    289.9252, 289.4634, 289.9805, 288.0692, 289.0663, 287.5041, 287.9754, 
    288.3033, 288.1604, 288.904, 289.0789, 289.8001, 289.4223, 291.6214, 
    290.6528, 293.3441, 292.5913, 287.5096, 287.749, 288.579, 288.1852, 
    289.3119, 289.5888, 289.8252, 290.1129, 290.1443, 290.3149, 290.0354, 
    290.304, 289.2768, 289.7417, 288.4851, 288.7881, 288.6489, 288.4958, 
    288.9682, 289.4704, 289.482, 289.6536, 290.1056, 289.3165, 291.7448, 
    290.2498, 288.0101, 288.4682, 288.5346, 288.3573, 289.561, 289.125, 
    290.3109, 289.9933, 290.5139, 290.2551, 290.217, 289.8849, 289.6779, 
    289.1448, 288.7198, 288.3832, 288.4615, 288.8313, 289.5013, 290.1468, 
    290.0076, 290.4743, 289.2303, 289.7575, 289.5468, 290.0792, 288.9267, 
    289.9069, 288.6784, 288.7854, 289.1163, 289.7919, 289.9404, 290.0974, 
    290.0007, 289.5185, 289.4417, 289.1085, 289.016, 288.7622, 288.5517, 
    288.7438, 288.9454, 289.5191, 290.0465, 290.6104, 290.7487, 291.4057, 
    290.8697, 291.753, 291.0002, 292.3045, 289.9644, 290.9798, 289.1317, 
    289.3297, 289.6977, 290.5196, 290.0767, 290.5951, 289.4387, 288.8436, 
    288.6906, 288.4035, 288.6972, 288.6733, 288.9544, 288.8641, 289.5381, 
    289.1762, 290.2158, 290.5912, 291.653, 292.3036, 292.9675, 293.2602, 
    293.3494, 293.3866 ;

 FSH_R =
  286.2084, 286.813, 286.6957, 287.183, 286.913, 287.2318, 286.3314, 
    286.8367, 286.5143, 286.2634, 288.1261, 287.2048, 289.0811, 288.4968, 
    289.9763, 288.9897, 290.1733, 289.949, 290.6263, 290.4323, 291.2972, 
    290.7159, 291.747, 291.1588, 291.2505, 290.6966, 287.3911, 288.011, 
    287.3541, 287.4426, 287.4031, 286.9183, 286.6732, 286.1629, 286.2557, 
    286.6308, 287.4824, 287.1942, 287.9223, 287.9059, 288.7125, 288.3496, 
    289.7132, 289.3182, 290.4404, 290.1607, 290.4272, 290.3465, 290.4282, 
    290.018, 290.1937, 289.833, 288.4174, 288.8301, 287.5948, 286.8476, 
    286.3534, 286.002, 286.0517, 286.1462, 286.633, 287.0917, 287.4405, 
    287.6736, 287.9035, 288.5943, 288.9608, 289.7905, 289.6434, 289.8932, 
    290.1329, 290.5345, 290.4684, 290.6452, 289.8871, 290.3907, 289.5487, 
    289.7866, 287.9628, 287.2721, 286.9755, 286.7181, 286.0898, 286.5235, 
    286.3525, 286.7601, 287.0188, 286.891, 287.68, 287.3733, 288.9826, 
    288.2916, 290.1049, 289.6736, 290.2084, 289.9356, 290.4028, 289.9824, 
    290.7112, 290.8697, 290.7614, 291.1784, 289.959, 290.4269, 286.8872, 
    286.9081, 287.0054, 286.5774, 286.5514, 286.1602, 286.5085, 286.6567, 
    287.034, 287.2565, 287.468, 287.9331, 288.4504, 289.1721, 289.7015, 
    290.0493, 289.8363, 290.0244, 289.814, 289.7155, 290.8101, 290.1951, 
    291.1184, 291.0674, 290.6493, 291.0732, 286.9227, 286.8028, 286.3855, 
    286.7121, 286.1176, 286.45, 286.6408, 287.379, 287.5418, 287.6917, 
    287.9887, 288.3682, 289.0314, 289.6193, 290.147, 290.1083, 290.1219, 
    290.2395, 289.9478, 290.2874, 290.3441, 290.1954, 291.0606, 290.8134, 
    291.0663, 290.9055, 286.8419, 287.0438, 286.9346, 287.1398, 286.995, 
    287.637, 287.8295, 288.7273, 288.3605, 288.945, 288.4202, 288.513, 
    288.9629, 288.4487, 289.5762, 288.8108, 290.2441, 289.4676, 290.292, 
    290.1447, 290.3889, 290.6074, 290.8828, 291.3903, 291.2729, 291.6978, 
    287.3449, 287.6061, 287.5837, 287.8575, 288.0599, 288.4973, 289.1966, 
    288.9338, 289.4167, 289.5135, 288.7801, 289.2299, 287.7814, 288.016, 
    287.8767, 287.3651, 288.9937, 288.16, 289.71, 289.2482, 290.5762, 
    289.9203, 291.2081, 291.7575, 292.2773, 292.8818, 287.7493, 287.5717, 
    287.8903, 288.3289, 288.7358, 289.2756, 289.3311, 289.432, 289.705, 
    289.9252, 289.4634, 289.9805, 288.0692, 289.0663, 287.5041, 287.9754, 
    288.3033, 288.1604, 288.904, 289.0789, 289.8001, 289.4223, 291.6214, 
    290.6528, 293.3441, 292.5913, 287.5096, 287.749, 288.579, 288.1852, 
    289.3119, 289.5888, 289.8252, 290.1129, 290.1443, 290.3149, 290.0354, 
    290.304, 289.2768, 289.7417, 288.4851, 288.7881, 288.6489, 288.4958, 
    288.9682, 289.4704, 289.482, 289.6536, 290.1056, 289.3165, 291.7448, 
    290.2498, 288.0101, 288.4682, 288.5346, 288.3573, 289.561, 289.125, 
    290.3109, 289.9933, 290.5139, 290.2551, 290.217, 289.8849, 289.6779, 
    289.1448, 288.7198, 288.3832, 288.4615, 288.8313, 289.5013, 290.1468, 
    290.0076, 290.4743, 289.2303, 289.7575, 289.5468, 290.0792, 288.9267, 
    289.9069, 288.6784, 288.7854, 289.1163, 289.7919, 289.9404, 290.0974, 
    290.0007, 289.5185, 289.4417, 289.1085, 289.016, 288.7622, 288.5517, 
    288.7438, 288.9454, 289.5191, 290.0465, 290.6104, 290.7487, 291.4057, 
    290.8697, 291.753, 291.0002, 292.3045, 289.9644, 290.9798, 289.1317, 
    289.3297, 289.6977, 290.5196, 290.0767, 290.5951, 289.4387, 288.8436, 
    288.6906, 288.4035, 288.6972, 288.6733, 288.9544, 288.8641, 289.5381, 
    289.1762, 290.2158, 290.5912, 291.653, 292.3036, 292.9675, 293.2602, 
    293.3494, 293.3866 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.10301, -13.10401, -13.10382, -13.10462, -13.10418, -13.1047, -13.10322, 
    -13.10404, -13.10352, -13.10311, -13.10614, -13.10465, -13.10773, 
    -13.10679, -13.10917, -13.10757, -13.10949, -13.10914, -13.11026, 
    -13.10994, -13.11133, -13.1104, -13.11209, -13.11112, -13.11126, 
    -13.11037, -13.10497, -13.10595, -13.10491, -13.10505, -13.10499, 
    -13.10418, -13.10377, -13.10295, -13.1031, -13.10371, -13.10511, 
    -13.10465, -13.10586, -13.10583, -13.10714, -13.10656, -13.10875, 
    -13.10814, -13.10995, -13.10949, -13.10993, -13.10979, -13.10993, 
    -13.10925, -13.10954, -13.10895, -13.10666, -13.10733, -13.1053, 
    -13.10404, -13.10326, -13.10268, -13.10276, -13.10291, -13.10371, 
    -13.10448, -13.10506, -13.10544, -13.10583, -13.10692, -13.10753, 
    -13.10887, -13.10864, -13.10904, -13.10944, -13.1101, -13.10999, 
    -13.11028, -13.10904, -13.10986, -13.10852, -13.10888, -13.10586, 
    -13.10478, -13.10426, -13.10386, -13.10282, -13.10353, -13.10325, 
    -13.10393, -13.10436, -13.10415, -13.10546, -13.10495, -13.10757, 
    -13.10645, -13.1094, -13.10869, -13.10957, -13.10912, -13.10988, 
    -13.1092, -13.11039, -13.11064, -13.11047, -13.11116, -13.10916, 
    -13.10992, -13.10414, -13.10418, -13.10434, -13.10362, -13.10358, 
    -13.10294, -13.10352, -13.10375, -13.10439, -13.10475, -13.1051, 
    -13.10587, -13.10671, -13.10789, -13.10874, -13.10931, -13.10896, 
    -13.10927, -13.10892, -13.10876, -13.11055, -13.10954, -13.11106, 
    -13.11098, -13.11028, -13.11099, -13.1042, -13.10401, -13.10331, 
    -13.10386, -13.10287, -13.10341, -13.10372, -13.10494, -13.10523, 
    -13.10547, -13.10597, -13.10659, -13.10766, -13.10859, -13.10947, 
    -13.10941, -13.10943, -13.10962, -13.10914, -13.1097, -13.10978, 
    -13.10955, -13.11097, -13.11056, -13.11098, -13.11072, -13.10407, 
    -13.1044, -13.10422, -13.10455, -13.10431, -13.10536, -13.10568, 
    -13.10715, -13.10657, -13.10752, -13.10667, -13.10682, -13.10752, 
    -13.10672, -13.10854, -13.10728, -13.10962, -13.10835, -13.1097, 
    -13.10947, -13.10987, -13.11022, -13.11068, -13.1115, -13.11131, 
    -13.11202, -13.1049, -13.10532, -13.1053, -13.10575, -13.10608, -13.1068, 
    -13.10793, -13.10751, -13.1083, -13.10845, -13.10726, -13.10798, 
    -13.10561, -13.10599, -13.10578, -13.10492, -13.10759, -13.10623, 
    -13.10875, -13.10802, -13.11017, -13.10908, -13.11121, -13.11209, 
    -13.11298, -13.11397, -13.10557, -13.10528, -13.10581, -13.10651, 
    -13.10718, -13.10806, -13.10816, -13.10832, -13.10875, -13.10911, 
    -13.10836, -13.1092, -13.10605, -13.10772, -13.10516, -13.10592, 
    -13.10647, -13.10625, -13.10747, -13.10775, -13.10889, -13.10831, 
    -13.11186, -13.11028, -13.11476, -13.11349, -13.10517, -13.10557, 
    -13.10692, -13.10629, -13.10813, -13.10858, -13.10894, -13.1094, 
    -13.10946, -13.10974, -13.10929, -13.10972, -13.10806, -13.1088, 
    -13.10678, -13.10727, -13.10705, -13.1068, -13.10757, -13.10837, 
    -13.10841, -13.10865, -13.10933, -13.10814, -13.11203, -13.10957, 
    -13.106, -13.10673, -13.10686, -13.10657, -13.10853, -13.10782, 
    -13.10973, -13.10922, -13.11007, -13.10964, -13.10958, -13.10904, 
    -13.1087, -13.10785, -13.10716, -13.10662, -13.10674, -13.10734, 
    -13.10842, -13.10946, -13.10923, -13.11001, -13.10799, -13.10882, 
    -13.1085, -13.10935, -13.1075, -13.10902, -13.1071, -13.10727, -13.10781, 
    -13.10886, -13.10913, -13.10938, -13.10923, -13.10845, -13.10833, 
    -13.1078, -13.10764, -13.10723, -13.10689, -13.1072, -13.10752, 
    -13.10846, -13.10929, -13.11022, -13.11046, -13.1115, -13.11062, 
    -13.11204, -13.11079, -13.11298, -13.10913, -13.1108, -13.10784, 
    -13.10816, -13.10871, -13.11005, -13.10935, -13.11018, -13.10833, 
    -13.10735, -13.10712, -13.10665, -13.10713, -13.10709, -13.10755, 
    -13.1074, -13.10849, -13.10791, -13.10957, -13.11018, -13.11194, 
    -13.11301, -13.11413, -13.11462, -13.11478, -13.11484 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531 ;

 FSRND =
  0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505 ;

 FSRVD =
  0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.809094e-14, 2.821619e-14, 2.819177e-14, 2.829288e-14, 2.823673e-14, 
    2.830293e-14, 2.811618e-14, 2.822102e-14, 2.815403e-14, 2.810197e-14, 
    2.848916e-14, 2.82972e-14, 2.868852e-14, 2.856592e-14, 2.887386e-14, 
    2.866942e-14, 2.891508e-14, 2.886783e-14, 2.900978e-14, 2.896906e-14, 
    2.915084e-14, 2.902849e-14, 2.9245e-14, 2.912153e-14, 2.914084e-14, 
    2.902435e-14, 2.833592e-14, 2.846545e-14, 2.832822e-14, 2.834668e-14, 
    2.833835e-14, 2.823781e-14, 2.818722e-14, 2.808111e-14, 2.810031e-14, 
    2.817821e-14, 2.83548e-14, 2.829475e-14, 2.84459e-14, 2.844249e-14, 
    2.861096e-14, 2.853496e-14, 2.881838e-14, 2.873772e-14, 2.897073e-14, 
    2.891207e-14, 2.896793e-14, 2.895094e-14, 2.896808e-14, 2.888212e-14, 
    2.89189e-14, 2.884325e-14, 2.85495e-14, 2.863592e-14, 2.837821e-14, 
    2.822351e-14, 2.812068e-14, 2.804783e-14, 2.805808e-14, 2.807773e-14, 
    2.817861e-14, 2.827347e-14, 2.834583e-14, 2.839423e-14, 2.844193e-14, 
    2.858666e-14, 2.866315e-14, 2.883466e-14, 2.880362e-14, 2.885611e-14, 
    2.890621e-14, 2.89904e-14, 2.897652e-14, 2.901361e-14, 2.885455e-14, 
    2.896025e-14, 2.878575e-14, 2.883346e-14, 2.845536e-14, 2.831104e-14, 
    2.824991e-14, 2.819625e-14, 2.806598e-14, 2.815592e-14, 2.812044e-14, 
    2.820472e-14, 2.825834e-14, 2.823177e-14, 2.839553e-14, 2.833181e-14, 
    2.866764e-14, 2.852289e-14, 2.890039e-14, 2.880993e-14, 2.892199e-14, 
    2.886478e-14, 2.896279e-14, 2.887454e-14, 2.902737e-14, 2.90607e-14, 
    2.903787e-14, 2.91253e-14, 2.88695e-14, 2.89677e-14, 2.823118e-14, 
    2.823551e-14, 2.825562e-14, 2.816706e-14, 2.816162e-14, 2.808044e-14, 
    2.815259e-14, 2.818336e-14, 2.826137e-14, 2.830755e-14, 2.835145e-14, 
    2.844809e-14, 2.855609e-14, 2.870716e-14, 2.881577e-14, 2.888858e-14, 
    2.884388e-14, 2.888329e-14, 2.883919e-14, 2.881847e-14, 2.904815e-14, 
    2.891915e-14, 2.911265e-14, 2.910193e-14, 2.901431e-14, 2.910307e-14, 
    2.82385e-14, 2.821356e-14, 2.812718e-14, 2.819473e-14, 2.807156e-14, 
    2.81405e-14, 2.818014e-14, 2.833315e-14, 2.836671e-14, 2.839794e-14, 
    2.845954e-14, 2.853866e-14, 2.867762e-14, 2.879855e-14, 2.890901e-14, 
    2.890087e-14, 2.890372e-14, 2.892838e-14, 2.88672e-14, 2.893838e-14, 
    2.895032e-14, 2.891905e-14, 2.910043e-14, 2.904858e-14, 2.910161e-14, 
    2.90678e-14, 2.822162e-14, 2.826348e-14, 2.824081e-14, 2.82834e-14, 
    2.825336e-14, 2.838679e-14, 2.842679e-14, 2.861412e-14, 2.853712e-14, 
    2.865958e-14, 2.854949e-14, 2.8569e-14, 2.866358e-14, 2.855535e-14, 
    2.879184e-14, 2.863151e-14, 2.892932e-14, 2.876917e-14, 2.893931e-14, 
    2.890833e-14, 2.895951e-14, 2.900541e-14, 2.906308e-14, 2.91697e-14, 
    2.914494e-14, 2.92341e-14, 2.832591e-14, 2.838027e-14, 2.837543e-14, 
    2.843231e-14, 2.84744e-14, 2.856568e-14, 2.871219e-14, 2.865702e-14, 
    2.875817e-14, 2.877851e-14, 2.862471e-14, 2.871913e-14, 2.841641e-14, 
    2.846527e-14, 2.843612e-14, 2.832985e-14, 2.866957e-14, 2.849511e-14, 
    2.881727e-14, 2.872264e-14, 2.89988e-14, 2.886144e-14, 2.913134e-14, 
    2.924696e-14, 2.935561e-14, 2.948288e-14, 2.84099e-14, 2.837289e-14, 
    2.843902e-14, 2.853069e-14, 2.861561e-14, 2.872871e-14, 2.874023e-14, 
    2.87614e-14, 2.881627e-14, 2.886247e-14, 2.876809e-14, 2.887397e-14, 
    2.847667e-14, 2.868469e-14, 2.835863e-14, 2.845679e-14, 2.852492e-14, 
    2.849497e-14, 2.865038e-14, 2.868702e-14, 2.883609e-14, 2.875898e-14, 
    2.921838e-14, 2.901498e-14, 2.957967e-14, 2.942173e-14, 2.835996e-14, 
    2.840965e-14, 2.858286e-14, 2.850041e-14, 2.873617e-14, 2.879429e-14, 
    2.884145e-14, 2.890191e-14, 2.890835e-14, 2.894417e-14, 2.888543e-14, 
    2.894179e-14, 2.872868e-14, 2.882386e-14, 2.856273e-14, 2.862623e-14, 
    2.859697e-14, 2.856489e-14, 2.866378e-14, 2.87693e-14, 2.877146e-14, 
    2.880528e-14, 2.890083e-14, 2.873667e-14, 2.924467e-14, 2.893085e-14, 
    2.846387e-14, 2.855977e-14, 2.857337e-14, 2.853621e-14, 2.878839e-14, 
    2.869697e-14, 2.894329e-14, 2.887662e-14, 2.898575e-14, 2.893151e-14, 
    2.892348e-14, 2.885382e-14, 2.881043e-14, 2.870098e-14, 2.86119e-14, 
    2.85413e-14, 2.855765e-14, 2.863522e-14, 2.877567e-14, 2.890866e-14, 
    2.88795e-14, 2.897714e-14, 2.871855e-14, 2.882697e-14, 2.878503e-14, 
    2.889426e-14, 2.865546e-14, 2.885943e-14, 2.860336e-14, 2.862575e-14, 
    2.869508e-14, 2.883474e-14, 2.88655e-14, 2.889853e-14, 2.887808e-14, 
    2.877941e-14, 2.876319e-14, 2.869322e-14, 2.867391e-14, 2.862064e-14, 
    2.857651e-14, 2.86168e-14, 2.865907e-14, 2.877923e-14, 2.888759e-14, 
    2.900577e-14, 2.903468e-14, 2.917304e-14, 2.906044e-14, 2.924631e-14, 
    2.908837e-14, 2.936173e-14, 2.887109e-14, 2.908411e-14, 2.869823e-14, 
    2.87397e-14, 2.881487e-14, 2.898724e-14, 2.889404e-14, 2.900298e-14, 
    2.876254e-14, 2.863797e-14, 2.860565e-14, 2.854557e-14, 2.860698e-14, 
    2.860198e-14, 2.866078e-14, 2.864183e-14, 2.878315e-14, 2.870721e-14, 
    2.892297e-14, 2.900181e-14, 2.922449e-14, 2.936115e-14, 2.950027e-14, 
    2.956171e-14, 2.958041e-14, 2.958821e-14 ;

 F_DENIT_vr =
  1.604022e-12, 1.611174e-12, 1.609779e-12, 1.615553e-12, 1.612347e-12, 
    1.616127e-12, 1.605463e-12, 1.61145e-12, 1.607624e-12, 1.604651e-12, 
    1.62676e-12, 1.615799e-12, 1.638144e-12, 1.631144e-12, 1.648727e-12, 
    1.637053e-12, 1.651081e-12, 1.648383e-12, 1.656488e-12, 1.654163e-12, 
    1.664543e-12, 1.657557e-12, 1.66992e-12, 1.66287e-12, 1.663972e-12, 
    1.65732e-12, 1.618011e-12, 1.625407e-12, 1.617571e-12, 1.618625e-12, 
    1.618149e-12, 1.612408e-12, 1.609519e-12, 1.60346e-12, 1.604557e-12, 
    1.609005e-12, 1.619089e-12, 1.615659e-12, 1.62429e-12, 1.624096e-12, 
    1.633715e-12, 1.629376e-12, 1.645559e-12, 1.640953e-12, 1.654258e-12, 
    1.650909e-12, 1.654099e-12, 1.653129e-12, 1.654107e-12, 1.649199e-12, 
    1.651299e-12, 1.64698e-12, 1.630206e-12, 1.63514e-12, 1.620425e-12, 
    1.611591e-12, 1.60572e-12, 1.60156e-12, 1.602145e-12, 1.603267e-12, 
    1.609028e-12, 1.614444e-12, 1.618576e-12, 1.62134e-12, 1.624064e-12, 
    1.632328e-12, 1.636695e-12, 1.646489e-12, 1.644717e-12, 1.647713e-12, 
    1.650574e-12, 1.655382e-12, 1.654589e-12, 1.656707e-12, 1.647625e-12, 
    1.65366e-12, 1.643696e-12, 1.64642e-12, 1.624831e-12, 1.616589e-12, 
    1.613099e-12, 1.610035e-12, 1.602597e-12, 1.607732e-12, 1.605706e-12, 
    1.610519e-12, 1.61358e-12, 1.612063e-12, 1.621414e-12, 1.617775e-12, 
    1.636952e-12, 1.628687e-12, 1.650242e-12, 1.645077e-12, 1.651476e-12, 
    1.648209e-12, 1.653805e-12, 1.648766e-12, 1.657493e-12, 1.659396e-12, 
    1.658093e-12, 1.663085e-12, 1.648478e-12, 1.654086e-12, 1.612029e-12, 
    1.612277e-12, 1.613425e-12, 1.608368e-12, 1.608058e-12, 1.603422e-12, 
    1.607542e-12, 1.609299e-12, 1.613753e-12, 1.61639e-12, 1.618897e-12, 
    1.624415e-12, 1.630582e-12, 1.639209e-12, 1.64541e-12, 1.649568e-12, 
    1.647015e-12, 1.649266e-12, 1.646747e-12, 1.645565e-12, 1.658679e-12, 
    1.651314e-12, 1.662363e-12, 1.661751e-12, 1.656747e-12, 1.661815e-12, 
    1.612447e-12, 1.611023e-12, 1.606091e-12, 1.609948e-12, 1.602915e-12, 
    1.606852e-12, 1.609115e-12, 1.617852e-12, 1.619768e-12, 1.621552e-12, 
    1.625069e-12, 1.629587e-12, 1.637522e-12, 1.644427e-12, 1.650734e-12, 
    1.65027e-12, 1.650432e-12, 1.651841e-12, 1.648347e-12, 1.652411e-12, 
    1.653093e-12, 1.651308e-12, 1.661665e-12, 1.658704e-12, 1.661732e-12, 
    1.659801e-12, 1.611484e-12, 1.613874e-12, 1.612579e-12, 1.615011e-12, 
    1.613296e-12, 1.620915e-12, 1.623199e-12, 1.633896e-12, 1.629499e-12, 
    1.636492e-12, 1.630205e-12, 1.631319e-12, 1.63672e-12, 1.63054e-12, 
    1.644044e-12, 1.634889e-12, 1.651894e-12, 1.642749e-12, 1.652465e-12, 
    1.650695e-12, 1.653618e-12, 1.656239e-12, 1.659532e-12, 1.66562e-12, 
    1.664206e-12, 1.669297e-12, 1.617439e-12, 1.620543e-12, 1.620267e-12, 
    1.623515e-12, 1.625918e-12, 1.63113e-12, 1.639496e-12, 1.636345e-12, 
    1.642121e-12, 1.643283e-12, 1.634501e-12, 1.639892e-12, 1.622606e-12, 
    1.625397e-12, 1.623732e-12, 1.617663e-12, 1.637062e-12, 1.6271e-12, 
    1.645496e-12, 1.640092e-12, 1.655862e-12, 1.648018e-12, 1.663429e-12, 
    1.670032e-12, 1.676236e-12, 1.683503e-12, 1.622235e-12, 1.620122e-12, 
    1.623898e-12, 1.629132e-12, 1.633981e-12, 1.640439e-12, 1.641097e-12, 
    1.642306e-12, 1.645439e-12, 1.648077e-12, 1.642688e-12, 1.648734e-12, 
    1.626047e-12, 1.637925e-12, 1.619307e-12, 1.624912e-12, 1.628802e-12, 
    1.627092e-12, 1.635967e-12, 1.638058e-12, 1.646571e-12, 1.642168e-12, 
    1.6684e-12, 1.656785e-12, 1.68903e-12, 1.680011e-12, 1.619383e-12, 
    1.62222e-12, 1.632111e-12, 1.627403e-12, 1.640865e-12, 1.644184e-12, 
    1.646877e-12, 1.650329e-12, 1.650697e-12, 1.652742e-12, 1.649388e-12, 
    1.652606e-12, 1.640438e-12, 1.645872e-12, 1.630961e-12, 1.634587e-12, 
    1.632917e-12, 1.631085e-12, 1.636731e-12, 1.642757e-12, 1.64288e-12, 
    1.644811e-12, 1.650267e-12, 1.640893e-12, 1.669901e-12, 1.651981e-12, 
    1.625316e-12, 1.630792e-12, 1.631569e-12, 1.629447e-12, 1.643847e-12, 
    1.638627e-12, 1.652692e-12, 1.648885e-12, 1.655116e-12, 1.652019e-12, 
    1.651561e-12, 1.647583e-12, 1.645105e-12, 1.638856e-12, 1.633769e-12, 
    1.629738e-12, 1.630672e-12, 1.635101e-12, 1.643121e-12, 1.650714e-12, 
    1.649049e-12, 1.654625e-12, 1.639859e-12, 1.64605e-12, 1.643655e-12, 
    1.649892e-12, 1.636257e-12, 1.647903e-12, 1.633282e-12, 1.63456e-12, 
    1.638519e-12, 1.646493e-12, 1.64825e-12, 1.650136e-12, 1.648968e-12, 
    1.643334e-12, 1.642408e-12, 1.638412e-12, 1.63731e-12, 1.634268e-12, 
    1.631748e-12, 1.634049e-12, 1.636462e-12, 1.643324e-12, 1.649511e-12, 
    1.656259e-12, 1.65791e-12, 1.665811e-12, 1.659381e-12, 1.669995e-12, 
    1.660976e-12, 1.676585e-12, 1.648569e-12, 1.660732e-12, 1.638698e-12, 
    1.641067e-12, 1.645359e-12, 1.655201e-12, 1.64988e-12, 1.6561e-12, 
    1.64237e-12, 1.635258e-12, 1.633412e-12, 1.629982e-12, 1.633488e-12, 
    1.633203e-12, 1.63656e-12, 1.635478e-12, 1.643548e-12, 1.639211e-12, 
    1.651531e-12, 1.656033e-12, 1.668749e-12, 1.676552e-12, 1.684496e-12, 
    1.688004e-12, 1.689072e-12, 1.689517e-12,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  7.629381e-16, 7.636697e-16, 7.635265e-16, 7.641119e-16, 7.637866e-16, 
    7.641681e-16, 7.630832e-16, 7.636945e-16, 7.633038e-16, 7.629979e-16, 
    7.652265e-16, 7.641324e-16, 7.663338e-16, 7.656526e-16, 7.673468e-16, 
    7.662276e-16, 7.675691e-16, 7.673117e-16, 7.680758e-16, 7.678569e-16, 
    7.688236e-16, 7.681742e-16, 7.693141e-16, 7.686674e-16, 7.687688e-16, 
    7.681497e-16, 7.643578e-16, 7.650968e-16, 7.643127e-16, 7.644188e-16, 
    7.6437e-16, 7.637909e-16, 7.634979e-16, 7.628748e-16, 7.629871e-16, 
    7.634434e-16, 7.644615e-16, 7.641158e-16, 7.649769e-16, 7.649577e-16, 
    7.659011e-16, 7.654773e-16, 7.670419e-16, 7.665984e-16, 7.678652e-16, 
    7.675488e-16, 7.678494e-16, 7.677571e-16, 7.678487e-16, 7.673853e-16, 
    7.67583e-16, 7.671729e-16, 7.655651e-16, 7.660453e-16, 7.645975e-16, 
    7.637092e-16, 7.631077e-16, 7.626787e-16, 7.627381e-16, 7.628544e-16, 
    7.634448e-16, 7.63993e-16, 7.64408e-16, 7.646832e-16, 7.64953e-16, 
    7.657675e-16, 7.6619e-16, 7.671301e-16, 7.669596e-16, 7.672457e-16, 
    7.675165e-16, 7.679688e-16, 7.67894e-16, 7.68092e-16, 7.672338e-16, 
    7.678058e-16, 7.668569e-16, 7.671181e-16, 7.650376e-16, 7.642118e-16, 
    7.638611e-16, 7.635481e-16, 7.627845e-16, 7.633127e-16, 7.631044e-16, 
    7.635947e-16, 7.639051e-16, 7.637505e-16, 7.6469e-16, 7.643257e-16, 
    7.662139e-16, 7.654085e-16, 7.674858e-16, 7.66993e-16, 7.676008e-16, 
    7.672911e-16, 7.678198e-16, 7.67343e-16, 7.681641e-16, 7.683421e-16, 
    7.682192e-16, 7.686823e-16, 7.673125e-16, 7.678432e-16, 7.637503e-16, 
    7.637756e-16, 7.638911e-16, 7.63377e-16, 7.633448e-16, 7.628678e-16, 
    7.632902e-16, 7.634701e-16, 7.63921e-16, 7.641863e-16, 7.644371e-16, 
    7.649865e-16, 7.655933e-16, 7.664293e-16, 7.670243e-16, 7.674194e-16, 
    7.671763e-16, 7.673897e-16, 7.671499e-16, 7.670359e-16, 7.682739e-16, 
    7.675826e-16, 7.686141e-16, 7.685575e-16, 7.680917e-16, 7.68562e-16, 
    7.637918e-16, 7.636463e-16, 7.631429e-16, 7.635359e-16, 7.628144e-16, 
    7.632196e-16, 7.634508e-16, 7.643334e-16, 7.645237e-16, 7.647019e-16, 
    7.6505e-16, 7.65494e-16, 7.66266e-16, 7.669294e-16, 7.675293e-16, 
    7.674844e-16, 7.674996e-16, 7.676322e-16, 7.673009e-16, 7.67685e-16, 
    7.677489e-16, 7.675802e-16, 7.68548e-16, 7.682732e-16, 7.685537e-16, 
    7.683737e-16, 7.636924e-16, 7.639339e-16, 7.638022e-16, 7.640483e-16, 
    7.63874e-16, 7.646399e-16, 7.648666e-16, 7.659163e-16, 7.654855e-16, 
    7.66167e-16, 7.655535e-16, 7.656628e-16, 7.661888e-16, 7.655846e-16, 
    7.668917e-16, 7.660089e-16, 7.676367e-16, 7.667663e-16, 7.676895e-16, 
    7.675213e-16, 7.677964e-16, 7.680429e-16, 7.683488e-16, 7.689122e-16, 
    7.687807e-16, 7.692474e-16, 7.642923e-16, 7.646026e-16, 7.645741e-16, 
    7.648965e-16, 7.651339e-16, 7.656456e-16, 7.664562e-16, 7.661512e-16, 
    7.667069e-16, 7.668189e-16, 7.659706e-16, 7.664922e-16, 7.648024e-16, 
    7.650788e-16, 7.649129e-16, 7.643072e-16, 7.662171e-16, 7.652447e-16, 
    7.670263e-16, 7.665063e-16, 7.68006e-16, 7.672662e-16, 7.687087e-16, 
    7.693154e-16, 7.698743e-16, 7.705235e-16, 7.647701e-16, 7.645584e-16, 
    7.649333e-16, 7.654506e-16, 7.659222e-16, 7.665461e-16, 7.666084e-16, 
    7.667242e-16, 7.670239e-16, 7.672757e-16, 7.667604e-16, 7.673366e-16, 
    7.651439e-16, 7.663e-16, 7.644706e-16, 7.650291e-16, 7.654105e-16, 
    7.652422e-16, 7.661075e-16, 7.663089e-16, 7.671265e-16, 7.667038e-16, 
    7.691653e-16, 7.680911e-16, 7.710082e-16, 7.702118e-16, 7.644841e-16, 
    7.647661e-16, 7.657401e-16, 7.652785e-16, 7.665851e-16, 7.669047e-16, 
    7.671608e-16, 7.674896e-16, 7.675228e-16, 7.677164e-16, 7.673977e-16, 
    7.677023e-16, 7.665403e-16, 7.670621e-16, 7.656213e-16, 7.659741e-16, 
    7.65811e-16, 7.656315e-16, 7.661797e-16, 7.667613e-16, 7.667714e-16, 
    7.669564e-16, 7.674791e-16, 7.665782e-16, 7.693022e-16, 7.676389e-16, 
    7.650724e-16, 7.656112e-16, 7.656853e-16, 7.654776e-16, 7.66871e-16, 
    7.663689e-16, 7.677115e-16, 7.673503e-16, 7.679379e-16, 7.676466e-16, 
    7.676022e-16, 7.672248e-16, 7.669873e-16, 7.66387e-16, 7.658936e-16, 
    7.654998e-16, 7.6559e-16, 7.660221e-16, 7.667945e-16, 7.675184e-16, 
    7.673601e-16, 7.678851e-16, 7.664778e-16, 7.670729e-16, 7.668425e-16, 
    7.67437e-16, 7.661407e-16, 7.672623e-16, 7.65851e-16, 7.659745e-16, 
    7.66357e-16, 7.67124e-16, 7.672889e-16, 7.674685e-16, 7.673561e-16, 
    7.668188e-16, 7.667287e-16, 7.663431e-16, 7.662364e-16, 7.659413e-16, 
    7.656949e-16, 7.659193e-16, 7.661526e-16, 7.668132e-16, 7.674034e-16, 
    7.680384e-16, 7.681921e-16, 7.68925e-16, 7.683299e-16, 7.693083e-16, 
    7.684795e-16, 7.699021e-16, 7.673228e-16, 7.684656e-16, 7.663741e-16, 
    7.66601e-16, 7.670142e-16, 7.679462e-16, 7.674423e-16, 7.680295e-16, 
    7.667246e-16, 7.660388e-16, 7.658578e-16, 7.655231e-16, 7.658641e-16, 
    7.658364e-16, 7.661614e-16, 7.660558e-16, 7.668331e-16, 7.664158e-16, 
    7.675927e-16, 7.680167e-16, 7.691917e-16, 7.698981e-16, 7.706046e-16, 
    7.709129e-16, 7.710062e-16, 7.710446e-16 ;

 F_N2O_NIT =
  2.408274e-14, 2.429058e-14, 2.42501e-14, 2.441827e-14, 2.43249e-14, 
    2.443513e-14, 2.412479e-14, 2.429884e-14, 2.418765e-14, 2.410139e-14, 
    2.474633e-14, 2.442577e-14, 2.508157e-14, 2.487545e-14, 2.539489e-14, 
    2.504943e-14, 2.546484e-14, 2.538487e-14, 2.562591e-14, 2.555673e-14, 
    2.586632e-14, 2.565786e-14, 2.602755e-14, 2.581645e-14, 2.584942e-14, 
    2.565099e-14, 2.449012e-14, 2.470632e-14, 2.447733e-14, 2.45081e-14, 
    2.449429e-14, 2.432682e-14, 2.424266e-14, 2.406686e-14, 2.409872e-14, 
    2.422786e-14, 2.452192e-14, 2.442188e-14, 2.467437e-14, 2.466866e-14, 
    2.49513e-14, 2.482365e-14, 2.530119e-14, 2.516498e-14, 2.555961e-14, 
    2.546007e-14, 2.555493e-14, 2.552614e-14, 2.55553e-14, 2.540939e-14, 
    2.547184e-14, 2.534364e-14, 2.484756e-14, 2.499285e-14, 2.456082e-14, 
    2.430293e-14, 2.41324e-14, 2.401177e-14, 2.40288e-14, 2.406129e-14, 
    2.422861e-14, 2.438647e-14, 2.450712e-14, 2.4588e-14, 2.466783e-14, 
    2.491029e-14, 2.50391e-14, 2.532878e-14, 2.527637e-14, 2.536518e-14, 
    2.545017e-14, 2.55932e-14, 2.556963e-14, 2.563274e-14, 2.536282e-14, 
    2.554204e-14, 2.524652e-14, 2.532717e-14, 2.46896e-14, 2.444886e-14, 
    2.434692e-14, 2.425786e-14, 2.40419e-14, 2.419093e-14, 2.413212e-14, 
    2.427213e-14, 2.436132e-14, 2.431718e-14, 2.459021e-14, 2.448388e-14, 
    2.504674e-14, 2.480349e-14, 2.544025e-14, 2.528711e-14, 2.547702e-14, 
    2.538002e-14, 2.554634e-14, 2.539662e-14, 2.565625e-14, 2.571296e-14, 
    2.567419e-14, 2.582326e-14, 2.538832e-14, 2.55549e-14, 2.431596e-14, 
    2.432316e-14, 2.435669e-14, 2.420946e-14, 2.420047e-14, 2.406598e-14, 
    2.418562e-14, 2.423667e-14, 2.436649e-14, 2.444344e-14, 2.451672e-14, 
    2.467823e-14, 2.485925e-14, 2.511352e-14, 2.529702e-14, 2.542041e-14, 
    2.534471e-14, 2.541153e-14, 2.533683e-14, 2.530186e-14, 2.56917e-14, 
    2.547242e-14, 2.580179e-14, 2.578351e-14, 2.563422e-14, 2.578556e-14, 
    2.43282e-14, 2.428681e-14, 2.414338e-14, 2.425558e-14, 2.405135e-14, 
    2.416556e-14, 2.423136e-14, 2.44861e-14, 2.454224e-14, 2.459437e-14, 
    2.469749e-14, 2.483016e-14, 2.506378e-14, 2.526796e-14, 2.545511e-14, 
    2.544137e-14, 2.54462e-14, 2.54881e-14, 2.538438e-14, 2.550514e-14, 
    2.552544e-14, 2.547238e-14, 2.578105e-14, 2.569267e-14, 2.578311e-14, 
    2.572554e-14, 2.430026e-14, 2.436994e-14, 2.433227e-14, 2.440313e-14, 
    2.435319e-14, 2.457563e-14, 2.464252e-14, 2.495677e-14, 2.482754e-14, 
    2.503336e-14, 2.48484e-14, 2.488113e-14, 2.504009e-14, 2.485837e-14, 
    2.525668e-14, 2.498629e-14, 2.548972e-14, 2.521843e-14, 2.550677e-14, 
    2.545428e-14, 2.554121e-14, 2.56192e-14, 2.571748e-14, 2.589936e-14, 
    2.585718e-14, 2.600965e-14, 2.447402e-14, 2.456476e-14, 2.455676e-14, 
    2.465189e-14, 2.472236e-14, 2.487547e-14, 2.512206e-14, 2.502918e-14, 
    2.519981e-14, 2.523414e-14, 2.497495e-14, 2.513393e-14, 2.462556e-14, 
    2.470733e-14, 2.465862e-14, 2.448113e-14, 2.505055e-14, 2.475748e-14, 
    2.530003e-14, 2.514023e-14, 2.560807e-14, 2.537485e-14, 2.583397e-14, 
    2.603156e-14, 2.621821e-14, 2.643723e-14, 2.461435e-14, 2.455261e-14, 
    2.466321e-14, 2.481666e-14, 2.495947e-14, 2.514999e-14, 2.516952e-14, 
    2.520531e-14, 2.529813e-14, 2.537632e-14, 2.521663e-14, 2.539593e-14, 
    2.472632e-14, 2.507607e-14, 2.452925e-14, 2.469326e-14, 2.480757e-14, 
    2.475738e-14, 2.501854e-14, 2.508029e-14, 2.533207e-14, 2.520175e-14, 
    2.598272e-14, 2.563568e-14, 2.660461e-14, 2.633196e-14, 2.453105e-14, 
    2.461413e-14, 2.49044e-14, 2.476607e-14, 2.516273e-14, 2.526087e-14, 
    2.534078e-14, 2.544314e-14, 2.54542e-14, 2.551496e-14, 2.541543e-14, 
    2.551102e-14, 2.515037e-14, 2.53112e-14, 2.48711e-14, 2.497785e-14, 
    2.492871e-14, 2.487486e-14, 2.504123e-14, 2.521911e-14, 2.522291e-14, 
    2.528008e-14, 2.544159e-14, 2.516429e-14, 2.602769e-14, 2.549271e-14, 
    2.470488e-14, 2.486562e-14, 2.488862e-14, 2.482626e-14, 2.525101e-14, 
    2.509668e-14, 2.551348e-14, 2.540048e-14, 2.558575e-14, 2.54936e-14, 
    2.548005e-14, 2.536197e-14, 2.52886e-14, 2.510372e-14, 2.495381e-14, 
    2.483527e-14, 2.48628e-14, 2.499311e-14, 2.523e-14, 2.545517e-14, 
    2.540576e-14, 2.557161e-14, 2.51338e-14, 2.531691e-14, 2.524606e-14, 
    2.543101e-14, 2.50267e-14, 2.537085e-14, 2.493912e-14, 2.497682e-14, 
    2.509361e-14, 2.53294e-14, 2.53817e-14, 2.543763e-14, 2.540311e-14, 
    2.523605e-14, 2.520873e-14, 2.509075e-14, 2.505823e-14, 2.496858e-14, 
    2.489449e-14, 2.496218e-14, 2.503336e-14, 2.52361e-14, 2.541952e-14, 
    2.562028e-14, 2.566953e-14, 2.590539e-14, 2.571331e-14, 2.603068e-14, 
    2.576074e-14, 2.622892e-14, 2.539085e-14, 2.575286e-14, 2.509893e-14, 
    2.516896e-14, 2.529588e-14, 2.558823e-14, 2.543017e-14, 2.561506e-14, 
    2.520766e-14, 2.499762e-14, 2.494341e-14, 2.484246e-14, 2.494572e-14, 
    2.493731e-14, 2.503631e-14, 2.500447e-14, 2.524284e-14, 2.511465e-14, 
    2.547968e-14, 2.561357e-14, 2.599363e-14, 2.622805e-14, 2.646779e-14, 
    2.657398e-14, 2.660635e-14, 2.661989e-14 ;

 F_NIT =
  4.01379e-11, 4.04843e-11, 4.041683e-11, 4.069712e-11, 4.05415e-11, 
    4.072521e-11, 4.020798e-11, 4.049806e-11, 4.031275e-11, 4.016898e-11, 
    4.124388e-11, 4.070961e-11, 4.180262e-11, 4.145908e-11, 4.232481e-11, 
    4.174906e-11, 4.244139e-11, 4.230813e-11, 4.270985e-11, 4.259455e-11, 
    4.311054e-11, 4.27631e-11, 4.337926e-11, 4.302742e-11, 4.308236e-11, 
    4.275164e-11, 4.081686e-11, 4.11772e-11, 4.079555e-11, 4.084683e-11, 
    4.082381e-11, 4.05447e-11, 4.040443e-11, 4.011144e-11, 4.016454e-11, 
    4.037977e-11, 4.086986e-11, 4.070314e-11, 4.112395e-11, 4.111443e-11, 
    4.158549e-11, 4.137275e-11, 4.216865e-11, 4.194164e-11, 4.259935e-11, 
    4.243344e-11, 4.259155e-11, 4.254357e-11, 4.259216e-11, 4.234898e-11, 
    4.245307e-11, 4.223941e-11, 4.141261e-11, 4.165474e-11, 4.093471e-11, 
    4.050488e-11, 4.022066e-11, 4.001962e-11, 4.0048e-11, 4.010215e-11, 
    4.038102e-11, 4.064411e-11, 4.084521e-11, 4.098e-11, 4.111304e-11, 
    4.151715e-11, 4.173184e-11, 4.221463e-11, 4.212728e-11, 4.22753e-11, 
    4.241695e-11, 4.265533e-11, 4.261604e-11, 4.272124e-11, 4.227136e-11, 
    4.257008e-11, 4.207753e-11, 4.221195e-11, 4.114933e-11, 4.07481e-11, 
    4.05782e-11, 4.042976e-11, 4.006983e-11, 4.031821e-11, 4.02202e-11, 
    4.045355e-11, 4.06022e-11, 4.052864e-11, 4.098369e-11, 4.080646e-11, 
    4.174457e-11, 4.133914e-11, 4.240042e-11, 4.214519e-11, 4.24617e-11, 
    4.230004e-11, 4.257723e-11, 4.232771e-11, 4.276041e-11, 4.285494e-11, 
    4.279032e-11, 4.303877e-11, 4.231387e-11, 4.259151e-11, 4.05266e-11, 
    4.05386e-11, 4.059448e-11, 4.03491e-11, 4.033411e-11, 4.010996e-11, 
    4.030937e-11, 4.039444e-11, 4.061081e-11, 4.073908e-11, 4.08612e-11, 
    4.113038e-11, 4.143208e-11, 4.185587e-11, 4.21617e-11, 4.236735e-11, 
    4.224118e-11, 4.235256e-11, 4.222805e-11, 4.216976e-11, 4.28195e-11, 
    4.245403e-11, 4.300298e-11, 4.297251e-11, 4.272371e-11, 4.297593e-11, 
    4.054701e-11, 4.047801e-11, 4.023897e-11, 4.042598e-11, 4.008558e-11, 
    4.027594e-11, 4.038559e-11, 4.081016e-11, 4.090374e-11, 4.099062e-11, 
    4.116248e-11, 4.138359e-11, 4.177297e-11, 4.211327e-11, 4.242518e-11, 
    4.240228e-11, 4.241034e-11, 4.248016e-11, 4.23073e-11, 4.250857e-11, 
    4.25424e-11, 4.245397e-11, 4.296841e-11, 4.282111e-11, 4.297184e-11, 
    4.287589e-11, 4.050043e-11, 4.061657e-11, 4.055378e-11, 4.067188e-11, 
    4.058865e-11, 4.095938e-11, 4.107087e-11, 4.159462e-11, 4.137924e-11, 
    4.172227e-11, 4.141401e-11, 4.146854e-11, 4.173349e-11, 4.143062e-11, 
    4.209447e-11, 4.164381e-11, 4.248287e-11, 4.203071e-11, 4.251128e-11, 
    4.242379e-11, 4.256868e-11, 4.269867e-11, 4.286247e-11, 4.31656e-11, 
    4.309529e-11, 4.334942e-11, 4.079003e-11, 4.094126e-11, 4.092793e-11, 
    4.108647e-11, 4.120394e-11, 4.145912e-11, 4.18701e-11, 4.171529e-11, 
    4.199969e-11, 4.205691e-11, 4.162491e-11, 4.188988e-11, 4.10426e-11, 
    4.117888e-11, 4.10977e-11, 4.080189e-11, 4.175092e-11, 4.126246e-11, 
    4.216672e-11, 4.190038e-11, 4.268011e-11, 4.229141e-11, 4.305662e-11, 
    4.338594e-11, 4.369702e-11, 4.406205e-11, 4.102392e-11, 4.092101e-11, 
    4.110534e-11, 4.13611e-11, 4.159911e-11, 4.191665e-11, 4.19492e-11, 
    4.200885e-11, 4.216355e-11, 4.229386e-11, 4.202771e-11, 4.232655e-11, 
    4.121053e-11, 4.179345e-11, 4.088209e-11, 4.115544e-11, 4.134594e-11, 
    4.126231e-11, 4.169757e-11, 4.180049e-11, 4.222012e-11, 4.200292e-11, 
    4.330453e-11, 4.272613e-11, 4.434102e-11, 4.388661e-11, 4.088508e-11, 
    4.102354e-11, 4.150734e-11, 4.127678e-11, 4.193788e-11, 4.210144e-11, 
    4.223463e-11, 4.240524e-11, 4.242366e-11, 4.252493e-11, 4.235904e-11, 
    4.251836e-11, 4.191728e-11, 4.218534e-11, 4.145184e-11, 4.162975e-11, 
    4.154785e-11, 4.14581e-11, 4.173538e-11, 4.203185e-11, 4.203818e-11, 
    4.213347e-11, 4.240265e-11, 4.194049e-11, 4.337948e-11, 4.248784e-11, 
    4.11748e-11, 4.144271e-11, 4.148103e-11, 4.137709e-11, 4.208502e-11, 
    4.182779e-11, 4.252246e-11, 4.233413e-11, 4.264292e-11, 4.248933e-11, 
    4.246675e-11, 4.226995e-11, 4.214766e-11, 4.183954e-11, 4.158968e-11, 
    4.139211e-11, 4.1438e-11, 4.165518e-11, 4.205001e-11, 4.242529e-11, 
    4.234293e-11, 4.261936e-11, 4.188967e-11, 4.219486e-11, 4.207676e-11, 
    4.238502e-11, 4.171117e-11, 4.228475e-11, 4.156521e-11, 4.162803e-11, 
    4.182268e-11, 4.221566e-11, 4.230284e-11, 4.239606e-11, 4.233851e-11, 
    4.206008e-11, 4.201455e-11, 4.181792e-11, 4.176371e-11, 4.161431e-11, 
    4.149082e-11, 4.160363e-11, 4.172227e-11, 4.206016e-11, 4.236586e-11, 
    4.270047e-11, 4.278256e-11, 4.317565e-11, 4.285552e-11, 4.338446e-11, 
    4.293457e-11, 4.371487e-11, 4.231808e-11, 4.292144e-11, 4.183155e-11, 
    4.194826e-11, 4.21598e-11, 4.264705e-11, 4.238362e-11, 4.269177e-11, 
    4.201276e-11, 4.16627e-11, 4.157235e-11, 4.14041e-11, 4.15762e-11, 
    4.156218e-11, 4.172718e-11, 4.167412e-11, 4.207139e-11, 4.185775e-11, 
    4.246613e-11, 4.268928e-11, 4.332271e-11, 4.371341e-11, 4.411298e-11, 
    4.428997e-11, 4.434392e-11, 4.436648e-11 ;

 F_NIT_vr =
  2.343868e-10, 2.354246e-10, 2.352223e-10, 2.360599e-10, 2.355949e-10, 
    2.361431e-10, 2.345959e-10, 2.354642e-10, 2.349095e-10, 2.344781e-10, 
    2.376854e-10, 2.360954e-10, 2.393391e-10, 2.383229e-10, 2.408758e-10, 
    2.391803e-10, 2.412178e-10, 2.408263e-10, 2.420039e-10, 2.41666e-10, 
    2.431732e-10, 2.42159e-10, 2.43955e-10, 2.429305e-10, 2.430904e-10, 
    2.421244e-10, 2.364169e-10, 2.374891e-10, 2.36353e-10, 2.365058e-10, 
    2.364369e-10, 2.356035e-10, 2.351838e-10, 2.343053e-10, 2.344643e-10, 
    2.351094e-10, 2.365728e-10, 2.360754e-10, 2.373282e-10, 2.373e-10, 
    2.386962e-10, 2.380663e-10, 2.40416e-10, 2.397474e-10, 2.416798e-10, 
    2.411931e-10, 2.416565e-10, 2.415155e-10, 2.416576e-10, 2.409445e-10, 
    2.412495e-10, 2.406221e-10, 2.381871e-10, 2.389034e-10, 2.367671e-10, 
    2.354842e-10, 2.34633e-10, 2.340295e-10, 2.341143e-10, 2.34277e-10, 
    2.351127e-10, 2.35899e-10, 2.364988e-10, 2.368998e-10, 2.372952e-10, 
    2.384938e-10, 2.391284e-10, 2.405507e-10, 2.402937e-10, 2.407286e-10, 
    2.411444e-10, 2.418427e-10, 2.417276e-10, 2.420351e-10, 2.407158e-10, 
    2.415923e-10, 2.401454e-10, 2.405408e-10, 2.374052e-10, 2.362105e-10, 
    2.357032e-10, 2.35259e-10, 2.341797e-10, 2.349248e-10, 2.346307e-10, 
    2.353293e-10, 2.357736e-10, 2.355534e-10, 2.369105e-10, 2.363823e-10, 
    2.391657e-10, 2.379659e-10, 2.410962e-10, 2.403459e-10, 2.412754e-10, 
    2.408009e-10, 2.416135e-10, 2.408817e-10, 2.421493e-10, 2.424256e-10, 
    2.422363e-10, 2.429618e-10, 2.408397e-10, 2.416541e-10, 2.355486e-10, 
    2.355846e-10, 2.357513e-10, 2.350169e-10, 2.34972e-10, 2.342995e-10, 
    2.348972e-10, 2.35152e-10, 2.357987e-10, 2.361812e-10, 2.36545e-10, 
    2.37346e-10, 2.382409e-10, 2.394935e-10, 2.403942e-10, 2.409982e-10, 
    2.406275e-10, 2.409543e-10, 2.405884e-10, 2.404167e-10, 2.423214e-10, 
    2.412514e-10, 2.428567e-10, 2.427679e-10, 2.420406e-10, 2.427772e-10, 
    2.356092e-10, 2.354026e-10, 2.346867e-10, 2.352465e-10, 2.342258e-10, 
    2.347969e-10, 2.35125e-10, 2.36393e-10, 2.366715e-10, 2.369303e-10, 
    2.37441e-10, 2.380967e-10, 2.392485e-10, 2.402512e-10, 2.411677e-10, 
    2.411001e-10, 2.411236e-10, 2.413281e-10, 2.408207e-10, 2.414109e-10, 
    2.415098e-10, 2.412506e-10, 2.427553e-10, 2.423251e-10, 2.42765e-10, 
    2.424845e-10, 2.354694e-10, 2.358161e-10, 2.356282e-10, 2.35981e-10, 
    2.35732e-10, 2.368375e-10, 2.371689e-10, 2.387218e-10, 2.380838e-10, 
    2.390989e-10, 2.381864e-10, 2.38348e-10, 2.391312e-10, 2.38235e-10, 
    2.401953e-10, 2.388654e-10, 2.413358e-10, 2.400067e-10, 2.414186e-10, 
    2.411617e-10, 2.415862e-10, 2.419669e-10, 2.424453e-10, 2.433296e-10, 
    2.431242e-10, 2.438642e-10, 2.363335e-10, 2.367837e-10, 2.367439e-10, 
    2.372153e-10, 2.37564e-10, 2.383208e-10, 2.395353e-10, 2.39078e-10, 
    2.399167e-10, 2.400853e-10, 2.388101e-10, 2.395926e-10, 2.370829e-10, 
    2.374876e-10, 2.372463e-10, 2.363653e-10, 2.391813e-10, 2.377348e-10, 
    2.404063e-10, 2.396216e-10, 2.419119e-10, 2.407721e-10, 2.430113e-10, 
    2.439701e-10, 2.448727e-10, 2.459283e-10, 2.370295e-10, 2.367228e-10, 
    2.372709e-10, 2.380302e-10, 2.387345e-10, 2.396723e-10, 2.39768e-10, 
    2.399434e-10, 2.403984e-10, 2.407815e-10, 2.399984e-10, 2.408768e-10, 
    2.375813e-10, 2.393068e-10, 2.366039e-10, 2.374171e-10, 2.37982e-10, 
    2.37734e-10, 2.390226e-10, 2.393263e-10, 2.40562e-10, 2.39923e-10, 
    2.437327e-10, 2.420455e-10, 2.467324e-10, 2.454208e-10, 2.366156e-10, 
    2.370274e-10, 2.384627e-10, 2.377795e-10, 2.397342e-10, 2.402161e-10, 
    2.406072e-10, 2.411083e-10, 2.411619e-10, 2.414589e-10, 2.409718e-10, 
    2.414392e-10, 2.396717e-10, 2.40461e-10, 2.382959e-10, 2.388221e-10, 
    2.385797e-10, 2.383137e-10, 2.391335e-10, 2.40008e-10, 2.400264e-10, 
    2.403064e-10, 2.410971e-10, 2.397377e-10, 2.439497e-10, 2.413462e-10, 
    2.374767e-10, 2.38271e-10, 2.383843e-10, 2.380764e-10, 2.401671e-10, 
    2.39409e-10, 2.414517e-10, 2.408988e-10, 2.418039e-10, 2.413539e-10, 
    2.412872e-10, 2.407096e-10, 2.403495e-10, 2.394418e-10, 2.387031e-10, 
    2.381182e-10, 2.382537e-10, 2.388964e-10, 2.400608e-10, 2.411638e-10, 
    2.409218e-10, 2.417321e-10, 2.395874e-10, 2.404861e-10, 2.401382e-10, 
    2.410443e-10, 2.390648e-10, 2.407546e-10, 2.38633e-10, 2.388185e-10, 
    2.393932e-10, 2.405507e-10, 2.408064e-10, 2.410802e-10, 2.409107e-10, 
    2.400922e-10, 2.399578e-10, 2.393777e-10, 2.392173e-10, 2.387759e-10, 
    2.3841e-10, 2.387439e-10, 2.39094e-10, 2.400906e-10, 2.40989e-10, 
    2.419693e-10, 2.422093e-10, 2.433559e-10, 2.42422e-10, 2.43963e-10, 
    2.426523e-10, 2.449215e-10, 2.408518e-10, 2.426188e-10, 2.394194e-10, 
    2.397633e-10, 2.40386e-10, 2.418155e-10, 2.41043e-10, 2.419461e-10, 
    2.399524e-10, 2.38919e-10, 2.386516e-10, 2.381534e-10, 2.386625e-10, 
    2.386211e-10, 2.391086e-10, 2.389514e-10, 2.40123e-10, 2.394934e-10, 
    2.412823e-10, 2.419361e-10, 2.437838e-10, 2.449176e-10, 2.460731e-10, 
    2.465832e-10, 2.467385e-10, 2.468032e-10,
  1.334709e-10, 1.344787e-10, 1.342825e-10, 1.350969e-10, 1.34645e-10, 
    1.351785e-10, 1.33675e-10, 1.345187e-10, 1.339799e-10, 1.335616e-10, 
    1.366825e-10, 1.351333e-10, 1.382986e-10, 1.373056e-10, 1.39805e-10, 
    1.381438e-10, 1.401408e-10, 1.39757e-10, 1.409134e-10, 1.405817e-10, 
    1.420644e-10, 1.410665e-10, 1.428353e-10, 1.418259e-10, 1.419836e-10, 
    1.410336e-10, 1.354446e-10, 1.364892e-10, 1.353828e-10, 1.355315e-10, 
    1.354648e-10, 1.346543e-10, 1.342465e-10, 1.33394e-10, 1.335487e-10, 
    1.341748e-10, 1.355984e-10, 1.351146e-10, 1.363353e-10, 1.363077e-10, 
    1.376712e-10, 1.370558e-10, 1.39355e-10, 1.387002e-10, 1.405956e-10, 
    1.40118e-10, 1.405731e-10, 1.404351e-10, 1.405749e-10, 1.398748e-10, 
    1.401746e-10, 1.395591e-10, 1.37171e-10, 1.378713e-10, 1.357865e-10, 
    1.345385e-10, 1.33712e-10, 1.331266e-10, 1.332093e-10, 1.33367e-10, 
    1.341785e-10, 1.349432e-10, 1.35527e-10, 1.35918e-10, 1.363037e-10, 
    1.374735e-10, 1.380942e-10, 1.394875e-10, 1.392357e-10, 1.396624e-10, 
    1.400705e-10, 1.407566e-10, 1.406436e-10, 1.409462e-10, 1.396512e-10, 
    1.405114e-10, 1.390924e-10, 1.3948e-10, 1.364085e-10, 1.352451e-10, 
    1.347516e-10, 1.343202e-10, 1.332729e-10, 1.339958e-10, 1.337107e-10, 
    1.343895e-10, 1.348214e-10, 1.346077e-10, 1.359287e-10, 1.354146e-10, 
    1.38131e-10, 1.369585e-10, 1.400229e-10, 1.392874e-10, 1.401994e-10, 
    1.397338e-10, 1.405319e-10, 1.398135e-10, 1.410589e-10, 1.413306e-10, 
    1.411449e-10, 1.418587e-10, 1.397737e-10, 1.405731e-10, 1.346018e-10, 
    1.346366e-10, 1.34799e-10, 1.340857e-10, 1.340421e-10, 1.333898e-10, 
    1.339702e-10, 1.342176e-10, 1.348465e-10, 1.35219e-10, 1.355734e-10, 
    1.36354e-10, 1.372275e-10, 1.384526e-10, 1.39335e-10, 1.399277e-10, 
    1.395642e-10, 1.398851e-10, 1.395264e-10, 1.393583e-10, 1.412287e-10, 
    1.401774e-10, 1.417559e-10, 1.416684e-10, 1.409534e-10, 1.416783e-10, 
    1.346611e-10, 1.344606e-10, 1.337653e-10, 1.343093e-10, 1.333188e-10, 
    1.338729e-10, 1.341919e-10, 1.354253e-10, 1.356969e-10, 1.359488e-10, 
    1.36447e-10, 1.370873e-10, 1.382131e-10, 1.391954e-10, 1.400943e-10, 
    1.400284e-10, 1.400516e-10, 1.402526e-10, 1.397548e-10, 1.403344e-10, 
    1.404318e-10, 1.401773e-10, 1.416567e-10, 1.412335e-10, 1.416666e-10, 
    1.413909e-10, 1.345258e-10, 1.348632e-10, 1.346808e-10, 1.350239e-10, 
    1.347821e-10, 1.358582e-10, 1.361814e-10, 1.376976e-10, 1.370747e-10, 
    1.380666e-10, 1.371753e-10, 1.373331e-10, 1.38099e-10, 1.372235e-10, 
    1.391412e-10, 1.378399e-10, 1.402605e-10, 1.389572e-10, 1.403423e-10, 
    1.400904e-10, 1.405075e-10, 1.408814e-10, 1.413524e-10, 1.422227e-10, 
    1.42021e-10, 1.4275e-10, 1.353669e-10, 1.358057e-10, 1.357671e-10, 
    1.362268e-10, 1.365671e-10, 1.373058e-10, 1.384937e-10, 1.380465e-10, 
    1.388678e-10, 1.390329e-10, 1.377854e-10, 1.385508e-10, 1.360996e-10, 
    1.364946e-10, 1.362594e-10, 1.354015e-10, 1.381495e-10, 1.367367e-10, 
    1.393496e-10, 1.385813e-10, 1.408281e-10, 1.39709e-10, 1.4191e-10, 
    1.428546e-10, 1.437457e-10, 1.447894e-10, 1.360454e-10, 1.35747e-10, 
    1.362815e-10, 1.370221e-10, 1.377107e-10, 1.386281e-10, 1.387221e-10, 
    1.388942e-10, 1.393404e-10, 1.39716e-10, 1.389486e-10, 1.398103e-10, 
    1.365862e-10, 1.382724e-10, 1.356342e-10, 1.364267e-10, 1.369784e-10, 
    1.367363e-10, 1.379955e-10, 1.382929e-10, 1.395036e-10, 1.388773e-10, 
    1.426212e-10, 1.409604e-10, 1.455859e-10, 1.44288e-10, 1.356428e-10, 
    1.360444e-10, 1.374453e-10, 1.367781e-10, 1.386894e-10, 1.391613e-10, 
    1.395454e-10, 1.400369e-10, 1.4009e-10, 1.403815e-10, 1.399039e-10, 
    1.403627e-10, 1.3863e-10, 1.394033e-10, 1.372849e-10, 1.377995e-10, 
    1.375627e-10, 1.373031e-10, 1.381048e-10, 1.389607e-10, 1.38979e-10, 
    1.392539e-10, 1.400294e-10, 1.386972e-10, 1.42836e-10, 1.402747e-10, 
    1.364828e-10, 1.372583e-10, 1.373693e-10, 1.370686e-10, 1.39114e-10, 
    1.383716e-10, 1.403744e-10, 1.398321e-10, 1.407211e-10, 1.402791e-10, 
    1.402141e-10, 1.396472e-10, 1.392947e-10, 1.384056e-10, 1.376836e-10, 
    1.371122e-10, 1.37245e-10, 1.37873e-10, 1.390131e-10, 1.400948e-10, 
    1.398576e-10, 1.406535e-10, 1.385505e-10, 1.394309e-10, 1.390904e-10, 
    1.399789e-10, 1.380347e-10, 1.396896e-10, 1.376128e-10, 1.377944e-10, 
    1.383569e-10, 1.394906e-10, 1.39742e-10, 1.400105e-10, 1.398448e-10, 
    1.390421e-10, 1.389108e-10, 1.383432e-10, 1.381866e-10, 1.377549e-10, 
    1.373978e-10, 1.37724e-10, 1.380669e-10, 1.390425e-10, 1.399237e-10, 
    1.408867e-10, 1.411228e-10, 1.422516e-10, 1.413324e-10, 1.428503e-10, 
    1.415594e-10, 1.437967e-10, 1.397857e-10, 1.415215e-10, 1.383825e-10, 
    1.387195e-10, 1.393296e-10, 1.407329e-10, 1.399747e-10, 1.408616e-10, 
    1.389056e-10, 1.378947e-10, 1.376336e-10, 1.371469e-10, 1.376447e-10, 
    1.376042e-10, 1.380812e-10, 1.379278e-10, 1.390749e-10, 1.384583e-10, 
    1.402125e-10, 1.408546e-10, 1.426735e-10, 1.437927e-10, 1.449351e-10, 
    1.454404e-10, 1.455943e-10, 1.456587e-10,
  1.248463e-10, 1.259499e-10, 1.25735e-10, 1.266275e-10, 1.261321e-10, 
    1.267169e-10, 1.250697e-10, 1.259938e-10, 1.254035e-10, 1.249455e-10, 
    1.28367e-10, 1.266674e-10, 1.301426e-10, 1.290513e-10, 1.318002e-10, 
    1.299725e-10, 1.3217e-10, 1.317473e-10, 1.330212e-10, 1.326557e-10, 
    1.342906e-10, 1.3319e-10, 1.351414e-10, 1.340274e-10, 1.342014e-10, 
    1.331538e-10, 1.270087e-10, 1.281548e-10, 1.269409e-10, 1.27104e-10, 
    1.270308e-10, 1.261423e-10, 1.256955e-10, 1.247621e-10, 1.249314e-10, 
    1.256171e-10, 1.271774e-10, 1.266469e-10, 1.279859e-10, 1.279555e-10, 
    1.29453e-10, 1.287769e-10, 1.313048e-10, 1.305843e-10, 1.32671e-10, 
    1.321449e-10, 1.326463e-10, 1.324942e-10, 1.326482e-10, 1.31877e-10, 
    1.322072e-10, 1.315294e-10, 1.289035e-10, 1.296729e-10, 1.273837e-10, 
    1.260154e-10, 1.251102e-10, 1.244694e-10, 1.245599e-10, 1.247325e-10, 
    1.256211e-10, 1.26459e-10, 1.27099e-10, 1.27528e-10, 1.279512e-10, 
    1.292358e-10, 1.299179e-10, 1.314507e-10, 1.311736e-10, 1.316432e-10, 
    1.320926e-10, 1.328485e-10, 1.32724e-10, 1.330574e-10, 1.316308e-10, 
    1.325782e-10, 1.310158e-10, 1.314424e-10, 1.280662e-10, 1.267899e-10, 
    1.262489e-10, 1.257763e-10, 1.246295e-10, 1.25421e-10, 1.251087e-10, 
    1.258522e-10, 1.263255e-10, 1.260913e-10, 1.275397e-10, 1.269758e-10, 
    1.299584e-10, 1.286701e-10, 1.320402e-10, 1.312304e-10, 1.322346e-10, 
    1.317218e-10, 1.326009e-10, 1.318096e-10, 1.331816e-10, 1.334811e-10, 
    1.332764e-10, 1.340636e-10, 1.317658e-10, 1.326462e-10, 1.260848e-10, 
    1.261229e-10, 1.263009e-10, 1.255194e-10, 1.254717e-10, 1.247575e-10, 
    1.253929e-10, 1.256639e-10, 1.26353e-10, 1.267613e-10, 1.2715e-10, 
    1.280063e-10, 1.289656e-10, 1.303119e-10, 1.312828e-10, 1.319353e-10, 
    1.315351e-10, 1.318884e-10, 1.314935e-10, 1.313085e-10, 1.333689e-10, 
    1.322103e-10, 1.339502e-10, 1.338537e-10, 1.330653e-10, 1.338646e-10, 
    1.261498e-10, 1.259301e-10, 1.251686e-10, 1.257644e-10, 1.246798e-10, 
    1.252864e-10, 1.256357e-10, 1.269875e-10, 1.272854e-10, 1.275618e-10, 
    1.281085e-10, 1.288115e-10, 1.300487e-10, 1.311291e-10, 1.321188e-10, 
    1.320462e-10, 1.320717e-10, 1.322932e-10, 1.317449e-10, 1.323833e-10, 
    1.324905e-10, 1.322102e-10, 1.338408e-10, 1.333741e-10, 1.338517e-10, 
    1.335477e-10, 1.260015e-10, 1.263713e-10, 1.261714e-10, 1.265474e-10, 
    1.262824e-10, 1.274623e-10, 1.27817e-10, 1.294821e-10, 1.287977e-10, 
    1.298876e-10, 1.289082e-10, 1.290815e-10, 1.299232e-10, 1.289611e-10, 
    1.310695e-10, 1.296384e-10, 1.323018e-10, 1.308671e-10, 1.323919e-10, 
    1.321145e-10, 1.32574e-10, 1.32986e-10, 1.335052e-10, 1.344652e-10, 
    1.342427e-10, 1.350472e-10, 1.269235e-10, 1.274047e-10, 1.273624e-10, 
    1.278667e-10, 1.282403e-10, 1.290516e-10, 1.303572e-10, 1.298655e-10, 
    1.307687e-10, 1.309503e-10, 1.295785e-10, 1.3042e-10, 1.277272e-10, 
    1.281607e-10, 1.279026e-10, 1.269614e-10, 1.299787e-10, 1.284265e-10, 
    1.312989e-10, 1.304535e-10, 1.329272e-10, 1.316945e-10, 1.341202e-10, 
    1.351627e-10, 1.36147e-10, 1.373009e-10, 1.276677e-10, 1.273404e-10, 
    1.279268e-10, 1.287399e-10, 1.294964e-10, 1.30505e-10, 1.306084e-10, 
    1.307977e-10, 1.312888e-10, 1.317022e-10, 1.308576e-10, 1.31806e-10, 
    1.282612e-10, 1.301139e-10, 1.272167e-10, 1.280862e-10, 1.28692e-10, 
    1.284261e-10, 1.298094e-10, 1.301364e-10, 1.314684e-10, 1.307791e-10, 
    1.349051e-10, 1.330731e-10, 1.381822e-10, 1.367464e-10, 1.272261e-10, 
    1.276666e-10, 1.292048e-10, 1.28472e-10, 1.305725e-10, 1.310917e-10, 
    1.315144e-10, 1.320555e-10, 1.32114e-10, 1.324352e-10, 1.319091e-10, 
    1.324144e-10, 1.305071e-10, 1.31358e-10, 1.290286e-10, 1.29594e-10, 
    1.293338e-10, 1.290486e-10, 1.299296e-10, 1.308709e-10, 1.308911e-10, 
    1.311935e-10, 1.320473e-10, 1.30581e-10, 1.351422e-10, 1.323176e-10, 
    1.281477e-10, 1.289994e-10, 1.291213e-10, 1.287909e-10, 1.310396e-10, 
    1.302229e-10, 1.324273e-10, 1.3183e-10, 1.328093e-10, 1.323223e-10, 
    1.322507e-10, 1.316265e-10, 1.312385e-10, 1.302603e-10, 1.294667e-10, 
    1.288388e-10, 1.289847e-10, 1.296748e-10, 1.309286e-10, 1.321193e-10, 
    1.318581e-10, 1.327348e-10, 1.304197e-10, 1.313883e-10, 1.310136e-10, 
    1.319917e-10, 1.298525e-10, 1.316731e-10, 1.293888e-10, 1.295884e-10, 
    1.302067e-10, 1.314541e-10, 1.317308e-10, 1.320265e-10, 1.31844e-10, 
    1.309605e-10, 1.30816e-10, 1.301917e-10, 1.300195e-10, 1.29545e-10, 
    1.291526e-10, 1.295111e-10, 1.298879e-10, 1.309609e-10, 1.319309e-10, 
    1.329919e-10, 1.332521e-10, 1.344971e-10, 1.334832e-10, 1.35158e-10, 
    1.337335e-10, 1.362034e-10, 1.31779e-10, 1.336917e-10, 1.302349e-10, 
    1.306055e-10, 1.312769e-10, 1.328223e-10, 1.319871e-10, 1.329641e-10, 
    1.308103e-10, 1.296986e-10, 1.294117e-10, 1.28877e-10, 1.294239e-10, 
    1.293794e-10, 1.299036e-10, 1.29735e-10, 1.309965e-10, 1.303183e-10, 
    1.322489e-10, 1.329564e-10, 1.349628e-10, 1.361989e-10, 1.37462e-10, 
    1.380211e-10, 1.381915e-10, 1.382627e-10,
  1.280644e-10, 1.292798e-10, 1.29043e-10, 1.300265e-10, 1.294805e-10, 
    1.301251e-10, 1.283103e-10, 1.293281e-10, 1.286779e-10, 1.281736e-10, 
    1.319452e-10, 1.300704e-10, 1.339061e-10, 1.327005e-10, 1.35739e-10, 
    1.337182e-10, 1.361482e-10, 1.356805e-10, 1.370906e-10, 1.366859e-10, 
    1.384971e-10, 1.372775e-10, 1.394404e-10, 1.382053e-10, 1.383982e-10, 
    1.372374e-10, 1.304467e-10, 1.317111e-10, 1.303719e-10, 1.305518e-10, 
    1.304711e-10, 1.294918e-10, 1.289996e-10, 1.279717e-10, 1.28158e-10, 
    1.289131e-10, 1.306328e-10, 1.300478e-10, 1.315245e-10, 1.31491e-10, 
    1.331442e-10, 1.323976e-10, 1.35191e-10, 1.343942e-10, 1.367028e-10, 
    1.361204e-10, 1.366754e-10, 1.36507e-10, 1.366776e-10, 1.35824e-10, 
    1.361894e-10, 1.354394e-10, 1.325373e-10, 1.333871e-10, 1.308603e-10, 
    1.293521e-10, 1.283549e-10, 1.276496e-10, 1.277492e-10, 1.279391e-10, 
    1.289175e-10, 1.298407e-10, 1.305463e-10, 1.310193e-10, 1.314862e-10, 
    1.329043e-10, 1.336578e-10, 1.353524e-10, 1.350458e-10, 1.355653e-10, 
    1.360626e-10, 1.368993e-10, 1.367614e-10, 1.371307e-10, 1.355516e-10, 
    1.366001e-10, 1.348713e-10, 1.353431e-10, 1.316134e-10, 1.302055e-10, 
    1.296093e-10, 1.290885e-10, 1.278258e-10, 1.286972e-10, 1.283533e-10, 
    1.291721e-10, 1.296936e-10, 1.294356e-10, 1.310323e-10, 1.304104e-10, 
    1.337025e-10, 1.322797e-10, 1.360045e-10, 1.351087e-10, 1.362196e-10, 
    1.356522e-10, 1.366252e-10, 1.357494e-10, 1.372682e-10, 1.376e-10, 
    1.373732e-10, 1.382453e-10, 1.357009e-10, 1.366754e-10, 1.294283e-10, 
    1.294704e-10, 1.296665e-10, 1.288056e-10, 1.28753e-10, 1.279666e-10, 
    1.286662e-10, 1.289647e-10, 1.297239e-10, 1.30174e-10, 1.306025e-10, 
    1.315471e-10, 1.326059e-10, 1.340932e-10, 1.351667e-10, 1.358885e-10, 
    1.354457e-10, 1.358366e-10, 1.353996e-10, 1.35195e-10, 1.374756e-10, 
    1.361928e-10, 1.381197e-10, 1.380128e-10, 1.371395e-10, 1.380248e-10, 
    1.295e-10, 1.292579e-10, 1.284192e-10, 1.290753e-10, 1.278811e-10, 
    1.285489e-10, 1.289337e-10, 1.304234e-10, 1.307518e-10, 1.310567e-10, 
    1.316598e-10, 1.324358e-10, 1.338023e-10, 1.349967e-10, 1.360915e-10, 
    1.360111e-10, 1.360394e-10, 1.362845e-10, 1.356778e-10, 1.363843e-10, 
    1.36503e-10, 1.361927e-10, 1.379984e-10, 1.374814e-10, 1.380105e-10, 
    1.376737e-10, 1.293366e-10, 1.297441e-10, 1.295238e-10, 1.299382e-10, 
    1.296462e-10, 1.30947e-10, 1.313383e-10, 1.331763e-10, 1.324205e-10, 
    1.336244e-10, 1.325425e-10, 1.327339e-10, 1.336637e-10, 1.326009e-10, 
    1.349307e-10, 1.333491e-10, 1.362941e-10, 1.34707e-10, 1.363938e-10, 
    1.360868e-10, 1.365953e-10, 1.370516e-10, 1.376266e-10, 1.386906e-10, 
    1.384439e-10, 1.39336e-10, 1.303528e-10, 1.308835e-10, 1.308367e-10, 
    1.313931e-10, 1.318053e-10, 1.327008e-10, 1.341432e-10, 1.335999e-10, 
    1.345981e-10, 1.347989e-10, 1.332827e-10, 1.342127e-10, 1.312392e-10, 
    1.317175e-10, 1.314326e-10, 1.303946e-10, 1.33725e-10, 1.320108e-10, 
    1.351844e-10, 1.342497e-10, 1.369865e-10, 1.356221e-10, 1.383082e-10, 
    1.394641e-10, 1.405562e-10, 1.418376e-10, 1.311735e-10, 1.308124e-10, 
    1.314593e-10, 1.323568e-10, 1.331921e-10, 1.343066e-10, 1.344208e-10, 
    1.346302e-10, 1.351732e-10, 1.356306e-10, 1.346965e-10, 1.357454e-10, 
    1.318285e-10, 1.338743e-10, 1.30676e-10, 1.316352e-10, 1.323038e-10, 
    1.320103e-10, 1.335379e-10, 1.338991e-10, 1.353719e-10, 1.346096e-10, 
    1.391784e-10, 1.371481e-10, 1.428169e-10, 1.412217e-10, 1.306864e-10, 
    1.311723e-10, 1.328701e-10, 1.320609e-10, 1.343811e-10, 1.349552e-10, 
    1.354227e-10, 1.360215e-10, 1.360863e-10, 1.364417e-10, 1.358595e-10, 
    1.364187e-10, 1.34309e-10, 1.352498e-10, 1.326755e-10, 1.332999e-10, 
    1.330124e-10, 1.326975e-10, 1.336706e-10, 1.347111e-10, 1.347334e-10, 
    1.350679e-10, 1.360126e-10, 1.343906e-10, 1.394415e-10, 1.363117e-10, 
    1.317031e-10, 1.326433e-10, 1.327778e-10, 1.32413e-10, 1.348976e-10, 
    1.339948e-10, 1.36433e-10, 1.35772e-10, 1.368559e-10, 1.363168e-10, 
    1.362375e-10, 1.355468e-10, 1.351176e-10, 1.340361e-10, 1.331593e-10, 
    1.324659e-10, 1.32627e-10, 1.333892e-10, 1.347749e-10, 1.360921e-10, 
    1.358031e-10, 1.367734e-10, 1.342123e-10, 1.352834e-10, 1.348689e-10, 
    1.359509e-10, 1.335855e-10, 1.355986e-10, 1.330732e-10, 1.332937e-10, 
    1.339769e-10, 1.353562e-10, 1.356622e-10, 1.359894e-10, 1.357875e-10, 
    1.348102e-10, 1.346504e-10, 1.339603e-10, 1.337701e-10, 1.332457e-10, 
    1.328124e-10, 1.332083e-10, 1.336247e-10, 1.348106e-10, 1.358836e-10, 
    1.370581e-10, 1.373462e-10, 1.387261e-10, 1.376024e-10, 1.394591e-10, 
    1.378798e-10, 1.40619e-10, 1.357156e-10, 1.378335e-10, 1.34008e-10, 
    1.344177e-10, 1.351601e-10, 1.368704e-10, 1.359458e-10, 1.370274e-10, 
    1.346441e-10, 1.334155e-10, 1.330985e-10, 1.32508e-10, 1.33112e-10, 
    1.330628e-10, 1.336419e-10, 1.334557e-10, 1.3485e-10, 1.341002e-10, 
    1.362356e-10, 1.370188e-10, 1.392424e-10, 1.406139e-10, 1.420165e-10, 
    1.426379e-10, 1.428273e-10, 1.429065e-10,
  1.381445e-10, 1.394321e-10, 1.391812e-10, 1.402237e-10, 1.396449e-10, 
    1.403283e-10, 1.38405e-10, 1.394834e-10, 1.387944e-10, 1.382601e-10, 
    1.422596e-10, 1.402703e-10, 1.443426e-10, 1.430615e-10, 1.462921e-10, 
    1.441429e-10, 1.467277e-10, 1.462298e-10, 1.477312e-10, 1.473001e-10, 
    1.492304e-10, 1.479304e-10, 1.502366e-10, 1.489193e-10, 1.49125e-10, 
    1.478876e-10, 1.406693e-10, 1.420111e-10, 1.4059e-10, 1.407809e-10, 
    1.406952e-10, 1.396568e-10, 1.391353e-10, 1.380463e-10, 1.382437e-10, 
    1.390436e-10, 1.408667e-10, 1.402463e-10, 1.418128e-10, 1.417773e-10, 
    1.435328e-10, 1.427397e-10, 1.457089e-10, 1.448614e-10, 1.473181e-10, 
    1.466981e-10, 1.47289e-10, 1.471096e-10, 1.472913e-10, 1.463825e-10, 
    1.467715e-10, 1.459732e-10, 1.428881e-10, 1.437909e-10, 1.41108e-10, 
    1.395088e-10, 1.384522e-10, 1.377052e-10, 1.378107e-10, 1.380119e-10, 
    1.390483e-10, 1.400267e-10, 1.407749e-10, 1.412767e-10, 1.417722e-10, 
    1.432781e-10, 1.440787e-10, 1.458807e-10, 1.455544e-10, 1.461073e-10, 
    1.466365e-10, 1.475275e-10, 1.473806e-10, 1.477739e-10, 1.460926e-10, 
    1.472088e-10, 1.453688e-10, 1.458707e-10, 1.419074e-10, 1.404135e-10, 
    1.397815e-10, 1.392295e-10, 1.378918e-10, 1.388148e-10, 1.384505e-10, 
    1.39318e-10, 1.398708e-10, 1.395972e-10, 1.412905e-10, 1.406308e-10, 
    1.441262e-10, 1.426146e-10, 1.465747e-10, 1.456213e-10, 1.468037e-10, 
    1.461997e-10, 1.472355e-10, 1.463031e-10, 1.479205e-10, 1.48274e-10, 
    1.480324e-10, 1.489619e-10, 1.462515e-10, 1.47289e-10, 1.395895e-10, 
    1.396342e-10, 1.39842e-10, 1.389297e-10, 1.388739e-10, 1.380409e-10, 
    1.38782e-10, 1.390982e-10, 1.399028e-10, 1.403801e-10, 1.408346e-10, 
    1.418368e-10, 1.42961e-10, 1.445415e-10, 1.45683e-10, 1.464512e-10, 
    1.459799e-10, 1.463959e-10, 1.459309e-10, 1.457132e-10, 1.481415e-10, 
    1.467751e-10, 1.48828e-10, 1.487139e-10, 1.477833e-10, 1.487268e-10, 
    1.396655e-10, 1.394089e-10, 1.385203e-10, 1.392154e-10, 1.379504e-10, 
    1.386577e-10, 1.390654e-10, 1.406446e-10, 1.409929e-10, 1.413164e-10, 
    1.419564e-10, 1.427803e-10, 1.442322e-10, 1.455022e-10, 1.466672e-10, 
    1.465817e-10, 1.466118e-10, 1.468728e-10, 1.462269e-10, 1.46979e-10, 
    1.471055e-10, 1.46775e-10, 1.486987e-10, 1.481476e-10, 1.487115e-10, 
    1.483525e-10, 1.394923e-10, 1.399243e-10, 1.396907e-10, 1.401301e-10, 
    1.398205e-10, 1.412001e-10, 1.416152e-10, 1.43567e-10, 1.427641e-10, 
    1.440431e-10, 1.428936e-10, 1.43097e-10, 1.44085e-10, 1.429556e-10, 
    1.454321e-10, 1.437506e-10, 1.468829e-10, 1.451942e-10, 1.469891e-10, 
    1.466622e-10, 1.472037e-10, 1.476897e-10, 1.483024e-10, 1.494368e-10, 
    1.491736e-10, 1.501251e-10, 1.405697e-10, 1.411326e-10, 1.41083e-10, 
    1.416733e-10, 1.421108e-10, 1.430617e-10, 1.445945e-10, 1.44017e-10, 
    1.450782e-10, 1.452918e-10, 1.4368e-10, 1.446684e-10, 1.415101e-10, 
    1.420177e-10, 1.417153e-10, 1.40614e-10, 1.441501e-10, 1.423291e-10, 
    1.45702e-10, 1.447077e-10, 1.476203e-10, 1.461677e-10, 1.490289e-10, 
    1.50262e-10, 1.514276e-10, 1.527968e-10, 1.414403e-10, 1.410572e-10, 
    1.417436e-10, 1.426965e-10, 1.435837e-10, 1.447683e-10, 1.448897e-10, 
    1.451124e-10, 1.4569e-10, 1.461767e-10, 1.451829e-10, 1.462988e-10, 
    1.421357e-10, 1.443087e-10, 1.409126e-10, 1.419304e-10, 1.426402e-10, 
    1.423285e-10, 1.439511e-10, 1.44335e-10, 1.459015e-10, 1.450905e-10, 
    1.499571e-10, 1.477926e-10, 1.538439e-10, 1.521386e-10, 1.409235e-10, 
    1.41439e-10, 1.432416e-10, 1.423823e-10, 1.448475e-10, 1.454581e-10, 
    1.459555e-10, 1.465928e-10, 1.466617e-10, 1.470402e-10, 1.464203e-10, 
    1.470156e-10, 1.447708e-10, 1.457715e-10, 1.430348e-10, 1.436982e-10, 
    1.433928e-10, 1.430582e-10, 1.440922e-10, 1.451985e-10, 1.452221e-10, 
    1.45578e-10, 1.465836e-10, 1.448575e-10, 1.502381e-10, 1.46902e-10, 
    1.420023e-10, 1.430007e-10, 1.431435e-10, 1.427561e-10, 1.453968e-10, 
    1.444368e-10, 1.470309e-10, 1.463272e-10, 1.474812e-10, 1.469071e-10, 
    1.468227e-10, 1.460875e-10, 1.456308e-10, 1.444807e-10, 1.435488e-10, 
    1.428122e-10, 1.429833e-10, 1.437931e-10, 1.452664e-10, 1.46668e-10, 
    1.463603e-10, 1.473933e-10, 1.446679e-10, 1.458072e-10, 1.453663e-10, 
    1.465176e-10, 1.440017e-10, 1.461428e-10, 1.434574e-10, 1.436917e-10, 
    1.444178e-10, 1.458848e-10, 1.462103e-10, 1.465586e-10, 1.463436e-10, 
    1.453038e-10, 1.451338e-10, 1.444001e-10, 1.441979e-10, 1.436406e-10, 
    1.431802e-10, 1.436009e-10, 1.440434e-10, 1.453042e-10, 1.46446e-10, 
    1.476966e-10, 1.480036e-10, 1.494747e-10, 1.482767e-10, 1.502568e-10, 
    1.485726e-10, 1.514949e-10, 1.462673e-10, 1.48523e-10, 1.444508e-10, 
    1.448864e-10, 1.456762e-10, 1.474968e-10, 1.465122e-10, 1.47664e-10, 
    1.451272e-10, 1.438211e-10, 1.434842e-10, 1.42857e-10, 1.434985e-10, 
    1.434463e-10, 1.440617e-10, 1.438637e-10, 1.453462e-10, 1.445488e-10, 
    1.468207e-10, 1.476548e-10, 1.500253e-10, 1.514893e-10, 1.52988e-10, 
    1.536524e-10, 1.538549e-10, 1.539397e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24532.08, 24551.96, 24548.06, 24564.34, 24555.28, 24565.99, 24536.07, 
    24552.76, 24542.07, 24533.85, 24596.67, 24565.07, 24630.49, 24609.58, 
    24662.55, 24627.2, 24669.81, 24661.51, 24686.72, 24679.43, 24712.44, 
    24690.11, 24730.04, 24707.06, 24710.62, 24689.38, 24571.36, 24592.69, 
    24570.11, 24573.13, 24571.77, 24555.46, 24547.35, 24530.57, 24533.6, 
    24545.93, 24574.49, 24564.7, 24589.53, 24588.96, 24617.23, 24604.38, 
    24652.89, 24639, 24679.74, 24669.32, 24679.25, 24676.22, 24679.29, 
    24664.05, 24670.55, 24657.26, 24606.77, 24621.44, 24578.31, 24553.16, 
    24536.8, 24525.36, 24526.97, 24530.04, 24546, 24561.25, 24573.03, 24581, 
    24588.88, 24613.09, 24626.15, 24655.73, 24650.35, 24659.48, 24668.29, 
    24683.28, 24680.79, 24687.45, 24659.23, 24677.89, 24647.29, 24655.56, 
    24591.04, 24567.33, 24557.41, 24548.81, 24528.21, 24542.39, 24536.78, 
    24550.19, 24558.81, 24554.53, 24581.22, 24570.76, 24626.93, 24602.37, 
    24667.26, 24651.45, 24671.09, 24661.01, 24678.34, 24662.73, 24689.94, 
    24695.97, 24691.85, 24707.79, 24661.87, 24679.25, 24554.41, 24555.11, 
    24558.36, 24544.17, 24543.3, 24530.49, 24541.88, 24546.78, 24559.31, 
    24566.8, 24573.98, 24589.91, 24607.95, 24633.76, 24652.46, 24665.2, 
    24657.37, 24664.28, 24656.56, 24652.96, 24693.71, 24670.61, 24705.48, 
    24703.52, 24687.61, 24703.74, 24555.6, 24551.6, 24537.85, 24548.59, 
    24529.11, 24539.97, 24546.27, 24570.97, 24576.49, 24581.63, 24591.82, 
    24605.03, 24628.67, 24649.49, 24668.8, 24667.37, 24667.88, 24672.24, 
    24661.46, 24674.03, 24676.15, 24670.61, 24703.25, 24693.81, 24703.47, 
    24697.31, 24552.9, 24559.64, 24555.99, 24562.87, 24558.02, 24579.78, 
    24586.38, 24617.78, 24604.77, 24625.56, 24606.86, 24610.15, 24626.25, 
    24607.86, 24648.34, 24620.78, 24672.41, 24644.43, 24674.2, 24668.72, 
    24677.81, 24686.02, 24696.45, 24716.03, 24711.46, 24728.08, 24569.79, 
    24578.71, 24577.92, 24587.31, 24594.29, 24609.58, 24634.64, 24625.14, 
    24642.54, 24646.03, 24619.62, 24635.86, 24584.71, 24592.8, 24587.97, 
    24570.49, 24627.32, 24597.78, 24652.78, 24636.5, 24684.85, 24660.48, 
    24708.95, 24730.49, 24751.19, 24775.84, 24583.61, 24577.51, 24588.42, 
    24603.68, 24618.06, 24637.48, 24639.46, 24643.09, 24652.58, 24660.63, 
    24644.25, 24662.66, 24594.68, 24629.93, 24575.21, 24591.4, 24602.78, 
    24597.77, 24624.06, 24630.36, 24656.07, 24642.74, 24725.13, 24687.77, 
    24794.82, 24764.01, 24575.39, 24583.58, 24612.49, 24598.63, 24638.77, 
    24648.76, 24656.96, 24667.56, 24668.71, 24675.05, 24664.68, 24674.64, 
    24637.52, 24653.92, 24609.14, 24619.92, 24614.95, 24609.52, 24626.37, 
    24644.5, 24644.89, 24650.73, 24667.41, 24638.93, 24730.07, 24672.74, 
    24592.55, 24608.59, 24610.9, 24604.64, 24647.75, 24632.04, 24674.9, 
    24663.13, 24682.49, 24672.82, 24671.41, 24659.15, 24651.6, 24632.76, 
    24617.49, 24605.55, 24608.31, 24621.47, 24645.62, 24668.81, 24663.68, 
    24681.01, 24635.85, 24654.51, 24647.25, 24666.3, 24624.89, 24660.07, 
    24616, 24619.82, 24631.72, 24655.79, 24661.19, 24666.99, 24663.4, 
    24646.23, 24643.45, 24631.43, 24628.11, 24618.98, 24611.5, 24618.34, 
    24625.57, 24646.24, 24665.11, 24686.14, 24691.36, 24716.69, 24696.02, 
    24730.4, 24701.09, 24752.4, 24662.14, 24700.24, 24632.27, 24639.4, 
    24652.35, 24682.76, 24666.21, 24685.59, 24643.34, 24621.93, 24616.44, 
    24606.27, 24616.67, 24615.82, 24625.87, 24622.63, 24646.92, 24633.88, 
    24671.37, 24685.43, 24726.32, 24752.3, 24779.29, 24791.33, 24795.02, 
    24796.57 ;

 GC_ICE1 =
  17606.13, 17637.89, 17631.66, 17657.66, 17643.19, 17660.29, 17612.52, 
    17639.17, 17622.1, 17608.96, 17709.27, 17658.83, 17763.22, 17729.87, 
    17814.27, 17757.98, 17825.83, 17812.62, 17852.74, 17841.13, 17893.65, 
    17858.12, 17921.64, 17885.08, 17890.74, 17856.96, 17668.88, 17702.93, 
    17666.88, 17671.7, 17669.53, 17643.48, 17630.53, 17603.73, 17608.56, 
    17628.26, 17673.87, 17658.23, 17697.88, 17696.97, 17742.07, 17721.57, 
    17798.89, 17776.78, 17841.62, 17825.04, 17840.84, 17836.03, 17840.9, 
    17816.66, 17826.99, 17805.85, 17725.39, 17748.79, 17679.98, 17639.8, 
    17613.68, 17595.4, 17597.97, 17602.88, 17628.37, 17652.72, 17671.54, 
    17684.27, 17696.85, 17735.47, 17756.3, 17803.41, 17794.85, 17809.38, 
    17823.4, 17847.25, 17843.3, 17853.89, 17808.99, 17838.68, 17789.99, 
    17803.15, 17700.29, 17662.43, 17646.6, 17632.86, 17599.95, 17622.6, 
    17613.63, 17635.05, 17648.82, 17642, 17684.62, 17667.91, 17757.54, 
    17718.36, 17821.76, 17796.6, 17827.85, 17811.82, 17839.4, 17814.55, 
    17857.85, 17867.44, 17860.88, 17886.25, 17813.19, 17840.84, 17641.81, 
    17642.92, 17648.11, 17625.44, 17624.06, 17603.6, 17621.79, 17629.61, 
    17649.62, 17661.59, 17673.05, 17698.49, 17727.27, 17768.45, 17798.22, 
    17818.48, 17806.02, 17817.01, 17804.73, 17799.01, 17863.84, 17827.09, 
    17882.57, 17879.45, 17854.14, 17879.8, 17643.7, 17637.31, 17615.35, 
    17632.51, 17601.38, 17618.73, 17628.8, 17668.26, 17677.06, 17685.28, 
    17701.53, 17722.62, 17760.32, 17793.48, 17824.22, 17821.94, 17822.74, 
    17829.7, 17812.54, 17832.53, 17835.91, 17827.09, 17879.03, 17864.01, 
    17879.38, 17869.58, 17639.39, 17650.16, 17644.33, 17655.31, 17647.57, 
    17682.32, 17692.86, 17742.96, 17722.2, 17755.37, 17725.54, 17730.78, 
    17756.47, 17727.13, 17791.65, 17747.74, 17829.97, 17785.44, 17832.8, 
    17824.08, 17838.55, 17851.62, 17868.21, 17899.35, 17892.08, 17918.52, 
    17666.37, 17680.61, 17679.34, 17694.33, 17705.47, 17729.87, 17769.85, 
    17754.69, 17782.41, 17787.98, 17745.89, 17771.79, 17690.19, 17703.1, 
    17695.4, 17667.48, 17758.17, 17711.04, 17798.71, 17772.8, 17849.75, 
    17810.98, 17888.09, 17922.35, 17955.26, 17994.42, 17688.43, 17678.69, 
    17696.12, 17720.46, 17743.39, 17774.37, 17777.52, 17783.3, 17798.4, 
    17811.21, 17785.14, 17814.44, 17706.11, 17762.33, 17675.03, 17700.87, 
    17719.02, 17711.03, 17752.96, 17763.02, 17803.96, 17782.73, 17913.82, 
    17854.39, 18024.5, 17975.65, 17675.3, 17688.39, 17734.52, 17712.4, 
    17776.42, 17792.32, 17805.38, 17822.24, 17824.07, 17834.17, 17817.66, 
    17833.51, 17774.44, 17800.54, 17729.18, 17746.37, 17738.44, 17729.78, 
    17756.65, 17785.55, 17786.16, 17795.46, 17822, 17776.68, 17921.68, 
    17830.48, 17702.7, 17728.3, 17731.98, 17722, 17790.72, 17765.69, 
    17833.92, 17815.19, 17846, 17830.61, 17828.36, 17808.86, 17796.85, 
    17766.85, 17742.49, 17723.44, 17727.85, 17748.84, 17787.32, 17824.24, 
    17816.07, 17843.64, 17771.77, 17801.48, 17789.93, 17820.24, 17754.29, 
    17810.32, 17740.11, 17746.2, 17765.19, 17803.52, 17812.1, 17821.33, 
    17815.63, 17788.29, 17783.86, 17764.73, 17759.42, 17744.87, 17732.93, 
    17743.84, 17755.38, 17788.3, 17818.34, 17851.8, 17860.1, 17900.4, 
    17867.52, 17922.21, 17875.58, 17957.18, 17813.61, 17874.23, 17766.06, 
    17777.43, 17798.04, 17846.42, 17820.1, 17850.92, 17783.69, 17749.57, 
    17740.81, 17724.59, 17741.18, 17739.82, 17755.86, 17750.68, 17789.4, 
    17768.64, 17828.3, 17850.68, 17915.72, 17957.02, 17999.89, 18018.97, 
    18024.82, 18027.28 ;

 GC_LIQ1 =
  5232.775, 5234.804, 5234.406, 5236.067, 5235.142, 5236.235, 5233.183, 
    5234.885, 5233.795, 5232.956, 5239.376, 5236.142, 5242.855, 5240.704, 
    5246.206, 5242.518, 5246.967, 5246.097, 5248.74, 5247.975, 5251.442, 
    5249.096, 5253.291, 5250.876, 5251.25, 5249.019, 5236.784, 5238.967, 
    5236.656, 5236.964, 5236.826, 5235.161, 5234.333, 5232.621, 5232.93, 
    5234.188, 5237.103, 5236.103, 5238.642, 5238.584, 5241.491, 5240.169, 
    5245.193, 5243.738, 5248.007, 5246.915, 5247.956, 5247.639, 5247.959, 
    5246.363, 5247.043, 5245.651, 5240.416, 5241.924, 5237.494, 5234.926, 
    5233.257, 5232.09, 5232.254, 5232.567, 5234.195, 5235.751, 5236.954, 
    5237.768, 5238.576, 5241.065, 5242.409, 5245.49, 5244.927, 5245.884, 
    5246.807, 5248.378, 5248.118, 5248.816, 5245.858, 5247.814, 5244.607, 
    5245.473, 5238.797, 5236.372, 5235.36, 5234.482, 5232.38, 5233.827, 
    5233.254, 5234.623, 5235.502, 5235.066, 5237.79, 5236.722, 5242.489, 
    5239.962, 5246.699, 5245.042, 5247.1, 5246.044, 5247.861, 5246.224, 
    5249.078, 5249.711, 5249.278, 5250.953, 5246.134, 5247.956, 5235.054, 
    5235.125, 5235.456, 5234.008, 5233.92, 5232.613, 5233.775, 5234.274, 
    5235.553, 5236.318, 5237.051, 5238.682, 5240.537, 5243.193, 5245.148, 
    5246.483, 5245.662, 5246.386, 5245.577, 5245.201, 5249.474, 5247.05, 
    5250.71, 5250.504, 5248.833, 5250.527, 5235.175, 5234.767, 5233.364, 
    5234.46, 5232.472, 5233.58, 5234.223, 5236.744, 5237.307, 5237.832, 
    5238.877, 5240.236, 5242.668, 5244.837, 5246.861, 5246.711, 5246.764, 
    5247.222, 5246.092, 5247.408, 5247.631, 5247.05, 5250.476, 5249.484, 
    5250.5, 5249.852, 5234.899, 5235.587, 5235.215, 5235.917, 5235.422, 
    5237.643, 5238.319, 5241.548, 5240.209, 5242.349, 5240.424, 5240.763, 
    5242.42, 5240.527, 5244.716, 5241.856, 5247.239, 5244.307, 5247.426, 
    5246.852, 5247.805, 5248.667, 5249.762, 5251.818, 5251.338, 5253.084, 
    5236.623, 5237.534, 5237.453, 5238.414, 5239.131, 5240.704, 5243.283, 
    5242.305, 5244.108, 5244.475, 5241.738, 5243.409, 5238.147, 5238.978, 
    5238.482, 5236.695, 5242.53, 5239.49, 5245.181, 5243.476, 5248.543, 
    5245.989, 5251.075, 5253.338, 5255.52, 5258.138, 5238.034, 5237.411, 
    5238.529, 5240.098, 5241.576, 5243.579, 5243.786, 5244.167, 5245.161, 
    5246.004, 5244.288, 5246.217, 5239.172, 5242.798, 5237.177, 5238.835, 
    5240.004, 5239.489, 5242.194, 5242.843, 5245.526, 5244.129, 5252.774, 
    5248.85, 5260.183, 5256.872, 5237.194, 5238.032, 5241.004, 5239.578, 
    5243.714, 5244.761, 5245.62, 5246.73, 5246.851, 5247.516, 5246.429, 
    5247.473, 5243.583, 5245.301, 5240.659, 5241.768, 5241.256, 5240.698, 
    5242.432, 5244.314, 5244.355, 5244.967, 5246.714, 5243.731, 5253.294, 
    5247.273, 5238.953, 5240.603, 5240.84, 5240.196, 5244.655, 5243.015, 
    5247.5, 5246.266, 5248.296, 5247.282, 5247.134, 5245.849, 5245.059, 
    5243.09, 5241.518, 5240.29, 5240.574, 5241.928, 5244.431, 5246.862, 
    5246.324, 5248.14, 5243.408, 5245.363, 5244.603, 5246.599, 5242.279, 
    5245.946, 5241.364, 5241.757, 5242.983, 5245.498, 5246.063, 5246.67, 
    5246.295, 5244.496, 5244.204, 5242.953, 5242.61, 5241.671, 5240.901, 
    5241.605, 5242.35, 5244.496, 5246.474, 5248.679, 5249.227, 5251.888, 
    5249.716, 5253.329, 5250.249, 5255.647, 5246.162, 5250.159, 5243.039, 
    5243.78, 5245.137, 5248.324, 5246.589, 5248.621, 5244.192, 5241.975, 
    5241.409, 5240.364, 5241.434, 5241.346, 5242.38, 5242.046, 5244.568, 
    5243.205, 5247.13, 5248.604, 5252.9, 5255.636, 5258.508, 5259.806, 
    5260.205, 5260.372 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.955688e-09, 8.995069e-09, 8.987413e-09, 9.019177e-09, 9.001556e-09, 
    9.022355e-09, 8.963671e-09, 8.996632e-09, 8.97559e-09, 8.959232e-09, 
    9.080819e-09, 9.020593e-09, 9.143371e-09, 9.104964e-09, 9.201444e-09, 
    9.137396e-09, 9.214359e-09, 9.199596e-09, 9.244026e-09, 9.231298e-09, 
    9.288129e-09, 9.249901e-09, 9.317588e-09, 9.278999e-09, 9.285037e-09, 
    9.24864e-09, 9.032712e-09, 9.073321e-09, 9.030306e-09, 9.036097e-09, 
    9.033498e-09, 9.00192e-09, 8.986007e-09, 8.952677e-09, 8.958728e-09, 
    8.983207e-09, 9.038701e-09, 9.019863e-09, 9.067337e-09, 9.066265e-09, 
    9.119118e-09, 9.095288e-09, 9.184119e-09, 9.158872e-09, 9.231829e-09, 
    9.213482e-09, 9.230967e-09, 9.225665e-09, 9.231036e-09, 9.204127e-09, 
    9.215657e-09, 9.191978e-09, 9.099751e-09, 9.126857e-09, 9.046015e-09, 
    8.997406e-09, 8.965117e-09, 8.942204e-09, 8.945443e-09, 8.951619e-09, 
    8.983351e-09, 9.013184e-09, 9.035919e-09, 9.051127e-09, 9.066111e-09, 
    9.11147e-09, 9.135475e-09, 9.189225e-09, 9.179524e-09, 9.195958e-09, 
    9.211656e-09, 9.238013e-09, 9.233675e-09, 9.245287e-09, 9.195523e-09, 
    9.228597e-09, 9.173998e-09, 9.188932e-09, 9.070189e-09, 9.024945e-09, 
    9.005717e-09, 8.988884e-09, 8.947935e-09, 8.976214e-09, 8.965066e-09, 
    8.991586e-09, 9.008438e-09, 9.000104e-09, 9.051543e-09, 9.031544e-09, 
    9.136897e-09, 9.09152e-09, 9.209825e-09, 9.181515e-09, 9.216611e-09, 
    9.198702e-09, 9.229387e-09, 9.201771e-09, 9.249609e-09, 9.260026e-09, 
    9.252907e-09, 9.280251e-09, 9.20024e-09, 9.230968e-09, 8.99987e-09, 
    9.00123e-09, 9.007563e-09, 8.979725e-09, 8.978023e-09, 8.952511e-09, 
    8.975211e-09, 8.984878e-09, 9.009415e-09, 9.02393e-09, 9.037727e-09, 
    9.068063e-09, 9.101943e-09, 9.149317e-09, 9.18335e-09, 9.206164e-09, 
    9.192175e-09, 9.204525e-09, 9.190719e-09, 9.184248e-09, 9.256123e-09, 
    9.215764e-09, 9.276318e-09, 9.272967e-09, 9.245563e-09, 9.273345e-09, 
    9.002184e-09, 8.994362e-09, 8.967203e-09, 8.988457e-09, 8.949733e-09, 
    8.971409e-09, 8.983873e-09, 9.031964e-09, 9.042529e-09, 9.052326e-09, 
    9.071675e-09, 9.096508e-09, 9.140069e-09, 9.17797e-09, 9.212569e-09, 
    9.210034e-09, 9.210926e-09, 9.218656e-09, 9.19951e-09, 9.221799e-09, 
    9.22554e-09, 9.215759e-09, 9.272519e-09, 9.256302e-09, 9.272896e-09, 
    9.262338e-09, 8.996905e-09, 9.010066e-09, 9.002954e-09, 9.016329e-09, 
    9.006906e-09, 9.048804e-09, 9.061366e-09, 9.120142e-09, 9.096019e-09, 
    9.13441e-09, 9.099919e-09, 9.106031e-09, 9.135664e-09, 9.101782e-09, 
    9.175882e-09, 9.125646e-09, 9.218956e-09, 9.168794e-09, 9.2221e-09, 
    9.212419e-09, 9.228446e-09, 9.242802e-09, 9.26086e-09, 9.294181e-09, 
    9.286465e-09, 9.314331e-09, 9.029688e-09, 9.046761e-09, 9.045257e-09, 
    9.063123e-09, 9.076336e-09, 9.104973e-09, 9.150903e-09, 9.133631e-09, 
    9.165339e-09, 9.171704e-09, 9.123532e-09, 9.15311e-09, 9.058186e-09, 
    9.073523e-09, 9.064391e-09, 9.031035e-09, 9.137612e-09, 9.082918e-09, 
    9.183913e-09, 9.154284e-09, 9.240755e-09, 9.197752e-09, 9.282218e-09, 
    9.318327e-09, 9.352308e-09, 9.392024e-09, 9.056078e-09, 9.044477e-09, 
    9.065247e-09, 9.093984e-09, 9.120646e-09, 9.156092e-09, 9.159717e-09, 
    9.166358e-09, 9.183558e-09, 9.198019e-09, 9.168459e-09, 9.201645e-09, 
    9.077082e-09, 9.14236e-09, 9.040092e-09, 9.070889e-09, 9.09229e-09, 
    9.082902e-09, 9.131657e-09, 9.143148e-09, 9.189844e-09, 9.165705e-09, 
    9.309416e-09, 9.245834e-09, 9.422261e-09, 9.372958e-09, 9.040424e-09, 
    9.056038e-09, 9.110376e-09, 9.084522e-09, 9.158457e-09, 9.176657e-09, 
    9.19145e-09, 9.210362e-09, 9.212403e-09, 9.223609e-09, 9.205247e-09, 
    9.222884e-09, 9.156166e-09, 9.185981e-09, 9.104164e-09, 9.124078e-09, 
    9.114917e-09, 9.104868e-09, 9.135881e-09, 9.168924e-09, 9.169629e-09, 
    9.180224e-09, 9.210082e-09, 9.158756e-09, 9.317625e-09, 9.219514e-09, 
    9.073062e-09, 9.103136e-09, 9.10743e-09, 9.095781e-09, 9.174832e-09, 
    9.14619e-09, 9.223336e-09, 9.202486e-09, 9.236648e-09, 9.219672e-09, 
    9.217175e-09, 9.195372e-09, 9.181798e-09, 9.147503e-09, 9.119598e-09, 
    9.09747e-09, 9.102616e-09, 9.126922e-09, 9.170945e-09, 9.212589e-09, 
    9.203467e-09, 9.234052e-09, 9.153096e-09, 9.187043e-09, 9.173923e-09, 
    9.208133e-09, 9.133172e-09, 9.197009e-09, 9.116856e-09, 9.123883e-09, 
    9.14562e-09, 9.189346e-09, 9.199018e-09, 9.209348e-09, 9.202973e-09, 
    9.172062e-09, 9.166998e-09, 9.145092e-09, 9.139044e-09, 9.122353e-09, 
    9.108534e-09, 9.12116e-09, 9.134419e-09, 9.172075e-09, 9.206009e-09, 
    9.243006e-09, 9.25206e-09, 9.29529e-09, 9.2601e-09, 9.318171e-09, 
    9.268803e-09, 9.35426e-09, 9.200707e-09, 9.267349e-09, 9.14661e-09, 
    9.159617e-09, 9.183144e-09, 9.237104e-09, 9.207972e-09, 9.242042e-09, 
    9.166799e-09, 9.127762e-09, 9.11766e-09, 9.098816e-09, 9.118091e-09, 
    9.116524e-09, 9.134968e-09, 9.129041e-09, 9.173325e-09, 9.149537e-09, 
    9.217112e-09, 9.241772e-09, 9.31141e-09, 9.354101e-09, 9.397556e-09, 
    9.41674e-09, 9.422579e-09, 9.425021e-09 ;

 H2OCAN =
  0.05992923, 0.05991429, 0.05991713, 0.05990519, 0.05991171, 0.05990397, 
    0.05992607, 0.05991381, 0.05992156, 0.0599277, 0.05988227, 0.05990463, 
    0.05985794, 0.0598723, 0.0598357, 0.05986036, 0.05983064, 0.0598361, 
    0.05981884, 0.05982378, 0.05980222, 0.05981655, 0.05979044, 0.05980548, 
    0.05980325, 0.05981708, 0.05989985, 0.05988517, 0.05990079, 0.05989868, 
    0.05989955, 0.05991168, 0.05991797, 0.05993015, 0.05992789, 0.05991882, 
    0.05989773, 0.0599047, 0.05988648, 0.05988688, 0.0598669, 0.05987588, 
    0.05984206, 0.05985164, 0.05982357, 0.05983071, 0.05982396, 0.05982597, 
    0.05982393, 0.05983438, 0.05982992, 0.059839, 0.05987426, 0.05986403, 
    0.05989484, 0.05991382, 0.05992559, 0.05993413, 0.05993293, 0.05993069, 
    0.05991877, 0.05990725, 0.05989853, 0.05989273, 0.05988695, 0.05987038, 
    0.05986095, 0.05984026, 0.05984375, 0.05983764, 0.05983141, 0.05982126, 
    0.05982289, 0.05981848, 0.05983761, 0.05982501, 0.05984579, 0.05984016, 
    0.05988643, 0.05990278, 0.05991059, 0.05991662, 0.05993202, 0.05992145, 
    0.05992565, 0.05991543, 0.05990907, 0.05991217, 0.05989257, 0.05990025, 
    0.05986039, 0.05987748, 0.05983213, 0.05984301, 0.05982948, 0.05983634, 
    0.05982465, 0.05983517, 0.05981674, 0.05981283, 0.05981553, 0.05980479, 
    0.05983578, 0.05982406, 0.05991231, 0.05991181, 0.05990936, 0.05992014, 
    0.05992074, 0.05993027, 0.0599217, 0.05991813, 0.05990862, 0.05990317, 
    0.05989792, 0.05988631, 0.05987357, 0.05985551, 0.05984232, 0.05983347, 
    0.05983884, 0.05983411, 0.05983943, 0.05984187, 0.05981437, 0.05982995, 
    0.05980634, 0.05980762, 0.05981841, 0.05980747, 0.05991144, 0.05991435, 
    0.05992476, 0.05991662, 0.05993129, 0.05992322, 0.05991865, 0.05990031, 
    0.05989602, 0.05989236, 0.05988486, 0.05987542, 0.059859, 0.05984449, 
    0.059831, 0.05983197, 0.05983164, 0.05982872, 0.05983608, 0.0598275, 
    0.05982616, 0.05982982, 0.0598078, 0.0598141, 0.05980765, 0.05981173, 
    0.05991338, 0.05990843, 0.05991112, 0.05990612, 0.05990973, 0.05989394, 
    0.05988919, 0.05986677, 0.05987567, 0.05986121, 0.05987412, 0.0598719, 
    0.05986118, 0.05987336, 0.05984549, 0.0598648, 0.05982861, 0.05984845, 
    0.05982738, 0.05983106, 0.05982486, 0.05981942, 0.05981234, 0.05979955, 
    0.05980248, 0.05979156, 0.05990094, 0.05989459, 0.05989496, 0.05988815, 
    0.05988315, 0.05987217, 0.05985478, 0.05986127, 0.05984914, 0.05984677, 
    0.05986508, 0.05985403, 0.05989018, 0.0598845, 0.05988774, 0.05990056, 
    0.05986005, 0.05988087, 0.05984214, 0.05985345, 0.05982022, 0.05983702, 
    0.05980413, 0.05979044, 0.05977655, 0.05976129, 0.0598909, 0.05989525, 
    0.05988728, 0.05987665, 0.0598663, 0.05985279, 0.0598513, 0.05984883, 
    0.05984215, 0.05983662, 0.05984823, 0.05983521, 0.05988358, 0.05985814, 
    0.05989707, 0.05988556, 0.05987718, 0.05988064, 0.05986196, 0.05985761, 
    0.05983997, 0.05984899, 0.05979401, 0.05981854, 0.05974894, 0.05976874, 
    0.05989682, 0.05989082, 0.05987033, 0.05987999, 0.05985179, 0.0598449, 
    0.05983911, 0.05983201, 0.0598311, 0.05982685, 0.05983383, 0.05982705, 
    0.05985277, 0.05984129, 0.05987242, 0.05986499, 0.05986834, 0.05987216, 
    0.05986037, 0.0598481, 0.05984752, 0.05984363, 0.05983318, 0.05985167, 
    0.05979141, 0.05982939, 0.05988429, 0.05987324, 0.05987129, 0.05987561, 
    0.0598456, 0.05985655, 0.05982691, 0.05983489, 0.05982171, 0.0598283, 
    0.05982928, 0.05983764, 0.05984291, 0.05985611, 0.05986672, 0.05987495, 
    0.05987301, 0.05986396, 0.05984727, 0.05983116, 0.05983474, 0.05982271, 
    0.05985385, 0.05984102, 0.05984609, 0.05983277, 0.05986151, 0.05983803, 
    0.0598676, 0.05986495, 0.05985676, 0.05984036, 0.05983623, 0.0598324, 
    0.0598347, 0.05984679, 0.05984862, 0.05985688, 0.05985932, 0.0598655, 
    0.05987076, 0.05986604, 0.05986113, 0.05984665, 0.05983371, 0.05981939, 
    0.05981574, 0.05979966, 0.0598132, 0.05979127, 0.0598106, 0.05977669, 
    0.05983619, 0.05981051, 0.05985628, 0.05985132, 0.05984267, 0.05982197, 
    0.05983283, 0.05981997, 0.05984867, 0.05986381, 0.05986732, 0.0598745, 
    0.05986715, 0.05986774, 0.0598607, 0.05986295, 0.05984617, 0.05985517, 
    0.0598294, 0.05981999, 0.05979282, 0.0597762, 0.05975863, 0.05975101, 
    0.05974865, 0.05974769 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.839474, 3.852424, 3.849903, 3.860369, 3.854561, 3.861418, 3.842096, 
    3.852938, 3.846014, 3.840638, 3.880749, 3.860837, 3.901524, 3.888758, 
    3.920886, 3.899535, 3.925203, 3.92027, 3.935134, 3.930871, 3.949932, 
    3.937103, 3.959843, 3.946865, 3.948893, 3.93668, 3.864838, 3.878265, 
    3.864043, 3.865955, 3.865097, 3.854681, 3.84944, 3.838486, 3.840473, 
    3.848519, 3.866815, 3.860597, 3.876286, 3.875931, 3.893459, 3.885548, 
    3.915103, 3.906687, 3.931049, 3.92491, 3.93076, 3.928986, 3.930783, 
    3.921783, 3.925637, 3.917726, 3.887029, 3.896031, 3.869232, 3.853193, 
    3.842571, 3.835049, 3.836112, 3.838138, 3.848567, 3.858394, 3.865897, 
    3.870923, 3.87588, 3.890917, 3.898896, 3.916806, 3.91357, 3.919054, 
    3.9243, 3.933119, 3.931666, 3.935556, 3.91891, 3.929966, 3.911728, 
    3.916709, 3.877227, 3.862273, 3.855931, 3.850388, 3.836929, 3.846219, 
    3.842554, 3.851278, 3.856829, 3.854083, 3.87106, 3.864452, 3.89937, 
    3.884298, 3.923688, 3.914234, 3.925956, 3.919971, 3.930231, 3.920996, 
    3.937004, 3.940497, 3.93811, 3.947286, 3.920485, 3.93076, 3.854006, 
    3.854454, 3.85654, 3.847374, 3.846814, 3.838431, 3.845889, 3.849069, 
    3.857151, 3.861938, 3.866494, 3.876526, 3.887756, 3.903503, 3.914846, 
    3.922464, 3.917792, 3.921917, 3.917306, 3.915146, 3.939188, 3.925673, 
    3.945965, 3.94484, 3.935648, 3.944967, 3.854768, 3.852191, 3.843257, 
    3.850247, 3.837519, 3.844639, 3.848738, 3.86459, 3.86808, 3.871319, 
    3.877722, 3.885953, 3.900425, 3.913052, 3.924605, 3.923758, 3.924056, 
    3.926641, 3.920241, 3.927692, 3.928943, 3.925672, 3.94469, 3.939249, 
    3.944816, 3.941273, 3.853029, 3.857366, 3.855022, 3.859431, 3.856324, 
    3.870154, 3.874309, 3.893799, 3.88579, 3.898542, 3.887084, 3.889112, 
    3.898958, 3.887703, 3.912354, 3.895628, 3.926741, 3.909991, 3.927793, 
    3.924555, 3.929917, 3.934723, 3.940777, 3.951967, 3.949374, 3.958747, 
    3.863839, 3.869479, 3.868982, 3.874891, 3.879266, 3.888762, 3.904032, 
    3.898284, 3.908841, 3.910962, 3.894926, 3.904767, 3.873257, 3.878333, 
    3.87531, 3.864284, 3.899607, 3.881446, 3.915034, 3.905158, 3.934037, 
    3.919653, 3.947947, 3.960092, 3.97155, 3.984973, 3.87256, 3.868725, 
    3.875594, 3.885115, 3.893967, 3.90576, 3.906968, 3.90918, 3.914916, 
    3.919744, 3.90988, 3.920954, 3.879511, 3.901187, 3.867275, 3.877461, 
    3.884553, 3.881441, 3.897628, 3.901451, 3.917013, 3.908963, 3.957091, 
    3.935739, 3.995219, 3.978525, 3.867385, 3.872547, 3.890555, 3.881978, 
    3.906549, 3.912614, 3.91755, 3.923867, 3.92455, 3.928297, 3.922158, 
    3.928055, 3.905785, 3.915724, 3.888493, 3.895108, 3.892064, 3.888727, 
    3.899033, 3.910035, 3.910271, 3.913803, 3.923771, 3.906648, 3.959853, 
    3.926925, 3.878182, 3.888151, 3.889577, 3.885712, 3.912005, 3.902462, 
    3.928206, 3.921235, 3.932662, 3.92698, 3.926145, 3.918859, 3.914328, 
    3.9029, 3.893619, 3.886272, 3.88798, 3.896053, 3.910709, 3.924612, 
    3.921563, 3.931793, 3.904763, 3.916078, 3.911702, 3.923122, 3.898131, 
    3.919403, 3.892708, 3.895043, 3.902273, 3.916847, 3.920077, 3.923528, 
    3.921398, 3.911081, 3.909394, 3.902097, 3.900084, 3.894534, 3.889944, 
    3.894138, 3.898546, 3.911086, 3.922412, 3.934792, 3.937826, 3.952338, 
    3.940521, 3.960037, 3.943439, 3.972207, 3.92064, 3.942952, 3.902603, 
    3.906935, 3.914777, 3.932814, 3.923069, 3.934468, 3.909327, 3.896332, 
    3.892975, 3.886719, 3.893118, 3.892597, 3.898729, 3.896758, 3.911503, 
    3.903578, 3.926124, 3.934378, 3.957763, 3.972155, 3.986847, 3.993347, 
    3.995327, 3.996155,
  3.319323, 3.332003, 3.329536, 3.339782, 3.334098, 3.340809, 3.321893, 
    3.332504, 3.325729, 3.320467, 3.35973, 3.340241, 3.380096, 3.367593, 
    3.399077, 3.378145, 3.403311, 3.398478, 3.413056, 3.408875, 3.42756, 
    3.414987, 3.437288, 3.424558, 3.426544, 3.414572, 3.344162, 3.357296, 
    3.343383, 3.345254, 3.344415, 3.334213, 3.329077, 3.31836, 3.320305, 
    3.328179, 3.346095, 3.340009, 3.355377, 3.35503, 3.372199, 3.364449, 
    3.393413, 3.385164, 3.40905, 3.403029, 3.408765, 3.407026, 3.408788, 
    3.399962, 3.403741, 3.395985, 3.365898, 3.374717, 3.348464, 3.332747, 
    3.322357, 3.314995, 3.316035, 3.318017, 3.328225, 3.337852, 3.345201, 
    3.350123, 3.35498, 3.369697, 3.377522, 3.395079, 3.391911, 3.397284, 
    3.402431, 3.411078, 3.409655, 3.413467, 3.397146, 3.407984, 3.390106, 
    3.394988, 3.356279, 3.341651, 3.33543, 3.330009, 3.316834, 3.325927, 
    3.32234, 3.330884, 3.336319, 3.333631, 3.350258, 3.343785, 3.377986, 
    3.363221, 3.40183, 3.392562, 3.404056, 3.398188, 3.408245, 3.399193, 
    3.414889, 3.418312, 3.415972, 3.424974, 3.398691, 3.408763, 3.333555, 
    3.333993, 3.336037, 3.327058, 3.32651, 3.318306, 3.325607, 3.328718, 
    3.336636, 3.341323, 3.345784, 3.35561, 3.366608, 3.382039, 3.393162, 
    3.400632, 3.396051, 3.400095, 3.395574, 3.393458, 3.417027, 3.403775, 
    3.423678, 3.422575, 3.413557, 3.4227, 3.334301, 3.331779, 3.323029, 
    3.329875, 3.317414, 3.324382, 3.328392, 3.343915, 3.347339, 3.350509, 
    3.356783, 3.364845, 3.379024, 3.3914, 3.402731, 3.401901, 3.402193, 
    3.404726, 3.398452, 3.405757, 3.406982, 3.403776, 3.422428, 3.417091, 
    3.422552, 3.419077, 3.332599, 3.336845, 3.33455, 3.338866, 3.335823, 
    3.349364, 3.353432, 3.372527, 3.364685, 3.377177, 3.365954, 3.36794, 
    3.377576, 3.366562, 3.390713, 3.374316, 3.404824, 3.388391, 3.405856, 
    3.402682, 3.40794, 3.412651, 3.41859, 3.429563, 3.42702, 3.436216, 
    3.343185, 3.348705, 3.348223, 3.35401, 3.358294, 3.367599, 3.38256, 
    3.376929, 3.387276, 3.389354, 3.37364, 3.383278, 3.352407, 3.357375, 
    3.354419, 3.343618, 3.37822, 3.360425, 3.393345, 3.383665, 3.411978, 
    3.39787, 3.42562, 3.437526, 3.448781, 3.461946, 3.351725, 3.34797, 
    3.3547, 3.36402, 3.372697, 3.384254, 3.38544, 3.387607, 3.393232, 
    3.397964, 3.388289, 3.399152, 3.35852, 3.37977, 3.346548, 3.356519, 
    3.363472, 3.360425, 3.376287, 3.380033, 3.395283, 3.387396, 3.434581, 
    3.413641, 3.47201, 3.455619, 3.346658, 3.351714, 3.369352, 3.360951, 
    3.385028, 3.390972, 3.395814, 3.402004, 3.402676, 3.406349, 3.400332, 
    3.406113, 3.384278, 3.394023, 3.367337, 3.373815, 3.370835, 3.367566, 
    3.377663, 3.38844, 3.388677, 3.392137, 3.40189, 3.385126, 3.437279, 
    3.404986, 3.357234, 3.366993, 3.368397, 3.364611, 3.390376, 3.381022, 
    3.406261, 3.399427, 3.410632, 3.40506, 3.40424, 3.397097, 3.392654, 
    3.38145, 3.372355, 3.365161, 3.366833, 3.37474, 3.389102, 3.402734, 
    3.399744, 3.409779, 3.383278, 3.394367, 3.390076, 3.401276, 3.376778, 
    3.397611, 3.371466, 3.373754, 3.380837, 3.395116, 3.398291, 3.401672, 
    3.399587, 3.389468, 3.387815, 3.380666, 3.378691, 3.373256, 3.368758, 
    3.372866, 3.377182, 3.389475, 3.400578, 3.412717, 3.415696, 3.429916, 
    3.418328, 3.437459, 3.421175, 3.449408, 3.398831, 3.42071, 3.381162, 
    3.385407, 3.393089, 3.410772, 3.401223, 3.412396, 3.387751, 3.37501, 
    3.371727, 3.365597, 3.371868, 3.371358, 3.377366, 3.375435, 3.389884, 
    3.382117, 3.404218, 3.412309, 3.435249, 3.449367, 3.463794, 3.470175, 
    3.472119, 3.472932,
  3.010891, 3.024971, 3.02223, 3.033613, 3.027295, 3.034755, 3.013742, 
    3.02553, 3.018001, 3.012157, 3.055793, 3.034122, 3.078022, 3.064518, 
    3.09849, 3.075921, 3.103057, 3.097839, 3.113567, 3.109055, 3.129234, 
    3.115651, 3.139735, 3.125987, 3.128134, 3.115203, 3.038475, 3.053089, 
    3.037611, 3.039691, 3.038758, 3.027425, 3.021726, 3.009818, 3.011977, 
    3.020725, 3.040627, 3.033861, 3.050936, 3.050549, 3.069506, 3.061021, 
    3.092375, 3.083477, 3.109243, 3.102748, 3.108938, 3.10706, 3.108962, 
    3.09944, 3.103517, 3.095149, 3.062634, 3.072222, 3.043257, 3.025806, 
    3.014258, 3.006083, 3.007237, 3.00944, 3.020776, 3.031464, 3.039628, 
    3.045097, 3.050494, 3.066821, 3.075247, 3.094176, 3.090754, 3.096553, 
    3.102103, 3.111434, 3.109897, 3.114013, 3.096401, 3.108097, 3.088806, 
    3.094074, 3.051959, 3.035685, 3.028785, 3.022757, 3.008126, 3.018224, 
    3.01424, 3.023725, 3.029762, 3.026775, 3.045247, 3.038056, 3.075747, 
    3.059659, 3.101455, 3.091456, 3.103855, 3.097524, 3.108377, 3.098608, 
    3.115546, 3.119244, 3.116717, 3.126433, 3.098067, 3.108937, 3.026691, 
    3.027178, 3.029448, 3.019479, 3.01887, 3.009758, 3.017866, 3.021323, 
    3.030113, 3.035321, 3.040277, 3.051197, 3.063425, 3.080113, 3.092104, 
    3.100161, 3.095219, 3.099581, 3.094705, 3.092421, 3.117858, 3.103555, 
    3.125034, 3.123843, 3.114111, 3.123977, 3.02752, 3.024718, 3.015004, 
    3.022604, 3.008767, 3.016506, 3.020963, 3.038205, 3.042004, 3.045529, 
    3.052499, 3.061462, 3.076862, 3.090205, 3.102426, 3.101529, 3.101845, 
    3.104579, 3.097809, 3.105691, 3.107015, 3.103554, 3.123683, 3.117923, 
    3.123817, 3.120066, 3.025629, 3.030346, 3.027797, 3.032592, 3.029213, 
    3.04426, 3.048782, 3.069864, 3.061285, 3.074873, 3.062694, 3.064903, 
    3.075311, 3.063368, 3.089468, 3.071795, 3.104685, 3.086968, 3.105798, 
    3.102373, 3.108045, 3.113132, 3.119541, 3.13139, 3.128644, 3.138573, 
    3.037389, 3.043526, 3.042985, 3.049417, 3.054179, 3.064522, 3.080672, 
    3.074601, 3.085754, 3.087997, 3.071056, 3.081448, 3.047638, 3.053164, 
    3.049873, 3.037872, 3.075998, 3.056553, 3.092302, 3.081861, 3.112406, 
    3.097187, 3.127132, 3.139997, 3.152144, 3.166379, 3.046879, 3.042705, 
    3.050183, 3.060549, 3.070043, 3.082497, 3.083774, 3.086113, 3.092177, 
    3.097283, 3.086852, 3.098564, 3.054446, 3.077667, 3.041127, 3.052214, 
    3.059937, 3.056548, 3.073908, 3.077945, 3.094394, 3.085883, 3.136817, 
    3.114206, 3.177253, 3.159539, 3.041247, 3.046865, 3.06644, 3.057133, 
    3.083331, 3.089742, 3.094963, 3.101644, 3.102367, 3.106332, 3.099837, 
    3.106075, 3.082524, 3.093032, 3.064229, 3.071247, 3.068034, 3.064484, 
    3.075392, 3.087016, 3.087265, 3.091, 3.10154, 3.083436, 3.139742, 
    3.104877, 3.052999, 3.063856, 3.065408, 3.061199, 3.089099, 3.079014, 
    3.106235, 3.098861, 3.110951, 3.104939, 3.104055, 3.096347, 3.091556, 
    3.079476, 3.069675, 3.06181, 3.063669, 3.072245, 3.087728, 3.102432, 
    3.099206, 3.110031, 3.081444, 3.093406, 3.088778, 3.100857, 3.07444, 
    3.09692, 3.068714, 3.071179, 3.078814, 3.094218, 3.097636, 3.101286, 
    3.099033, 3.088122, 3.086338, 3.078629, 3.076503, 3.070642, 3.065796, 
    3.070223, 3.074878, 3.088127, 3.100105, 3.113204, 3.116416, 3.131782, 
    3.119268, 3.139937, 3.122355, 3.152838, 3.098229, 3.121842, 3.079163, 
    3.083739, 3.09203, 3.11111, 3.1008, 3.112861, 3.086268, 3.072539, 
    3.068996, 3.062296, 3.069147, 3.068597, 3.075071, 3.07299, 3.088568, 
    3.080192, 3.104032, 3.112766, 3.137531, 3.152784, 3.168369, 3.175267, 
    3.177368, 3.178247,
  2.88864, 2.903944, 2.900964, 2.913344, 2.906471, 2.914585, 2.891737, 
    2.904553, 2.896366, 2.890014, 2.937405, 2.913897, 2.961275, 2.946599, 
    2.983575, 2.958988, 2.988553, 2.982863, 3.000012, 2.995091, 3.017113, 
    3.002285, 3.028578, 3.013566, 3.015911, 3.001797, 2.918632, 2.934543, 
    2.917692, 2.919956, 2.91894, 2.906613, 2.900418, 2.887472, 2.889819, 
    2.899328, 2.920974, 2.913612, 2.932193, 2.931772, 2.952001, 2.942912, 
    2.976908, 2.967213, 2.995296, 2.988214, 2.994963, 2.992916, 2.99499, 
    2.984609, 2.989053, 2.979931, 2.944613, 2.954957, 2.923836, 2.904855, 
    2.892298, 2.883414, 2.884669, 2.887062, 2.899384, 2.911005, 2.919886, 
    2.925838, 2.931712, 2.949082, 2.958253, 2.978872, 2.975142, 2.981463, 
    2.98751, 2.997687, 2.99601, 3.0005, 2.981295, 2.994048, 2.973019, 
    2.978759, 2.933314, 2.915596, 2.908094, 2.901537, 2.885634, 2.896609, 
    2.892279, 2.902588, 2.909154, 2.905905, 2.926001, 2.918176, 2.958797, 
    2.941477, 2.986804, 2.975907, 2.989421, 2.982519, 2.994353, 2.983701, 
    3.002172, 3.006207, 3.003449, 3.014052, 2.983111, 2.994964, 2.905814, 
    2.906344, 2.908813, 2.897974, 2.897312, 2.887408, 2.896219, 2.899978, 
    2.909535, 2.9152, 2.920593, 2.932478, 2.945448, 2.963552, 2.976612, 
    2.985393, 2.980006, 2.984762, 2.979446, 2.976957, 3.004695, 2.989095, 
    3.012525, 3.011225, 3.000607, 3.011371, 2.906716, 2.903669, 2.893108, 
    2.90137, 2.886331, 2.894742, 2.899587, 2.91834, 2.922472, 2.926308, 
    2.933896, 2.943376, 2.960011, 2.974545, 2.987862, 2.986885, 2.987229, 
    2.99021, 2.98283, 2.991423, 2.992867, 2.989093, 3.011051, 3.004764, 
    3.011197, 3.007102, 2.904659, 2.909789, 2.907016, 2.912232, 2.908557, 
    2.924929, 2.929851, 2.952392, 2.94319, 2.957845, 2.944676, 2.947006, 
    2.958325, 2.945386, 2.973742, 2.954495, 2.990326, 2.971021, 2.991539, 
    2.987805, 2.99399, 2.999538, 3.00653, 3.019465, 3.016466, 3.027308, 
    2.91745, 2.924129, 2.92354, 2.93054, 2.935699, 2.946603, 2.964159, 
    2.957547, 2.969694, 2.972138, 2.953687, 2.965005, 2.928604, 2.934622, 
    2.931037, 2.917977, 2.95907, 2.938203, 2.976829, 2.965455, 2.998747, 
    2.982153, 3.014816, 3.028867, 3.042136, 3.057704, 2.927778, 2.923234, 
    2.931373, 2.942415, 2.952584, 2.966147, 2.967538, 2.970085, 2.976692, 
    2.982256, 2.970892, 2.983652, 2.935984, 2.960887, 2.921519, 2.933587, 
    2.94177, 2.938196, 2.956792, 2.961189, 2.97911, 2.969835, 3.025395, 
    3.000712, 3.069598, 3.050223, 2.921648, 2.927762, 2.948664, 2.938813, 
    2.967054, 2.97404, 2.979728, 2.987012, 2.987798, 2.992122, 2.98504, 
    2.991842, 2.966177, 2.977624, 2.946294, 2.953895, 2.950396, 2.946563, 
    2.958408, 2.971071, 2.971341, 2.975411, 2.986905, 2.967169, 3.028594, 
    2.990543, 2.93444, 2.945903, 2.94754, 2.943099, 2.973339, 2.962353, 
    2.992016, 2.983976, 2.997159, 2.990602, 2.989639, 2.981237, 2.976015, 
    2.962857, 2.952184, 2.943743, 2.945704, 2.954983, 2.971846, 2.98787, 
    2.984354, 2.996155, 2.964999, 2.978032, 2.97299, 2.986152, 2.957372, 
    2.981869, 2.951137, 2.953821, 2.962136, 2.978919, 2.982641, 2.986621, 
    2.984164, 2.972275, 2.970331, 2.961933, 2.959618, 2.953236, 2.947961, 
    2.95278, 2.957849, 2.97228, 2.985334, 2.999618, 3.003121, 3.019897, 
    3.006236, 3.028807, 3.009611, 3.042901, 2.983292, 3.009046, 2.962514, 
    2.967499, 2.976534, 2.997336, 2.98609, 2.999245, 2.970255, 2.955303, 
    2.951444, 2.944256, 2.951608, 2.95101, 2.958058, 2.955792, 2.97276, 
    2.963636, 2.989615, 2.999141, 3.026171, 3.042838, 3.059876, 3.067424, 
    3.069723, 3.070685,
  2.94331, 2.959417, 2.956279, 2.969319, 2.962078, 2.970627, 2.946568, 
    2.960059, 2.95144, 2.944756, 2.994787, 2.969902, 3.020844, 3.004816, 
    3.045234, 3.018345, 3.050684, 3.044453, 3.063145, 3.057845, 3.081308, 
    3.065558, 3.093498, 3.077538, 3.08003, 3.06504, 2.974892, 2.991678, 
    2.973901, 2.976288, 2.975217, 2.962228, 2.955704, 2.942082, 2.94455, 
    2.954557, 2.977362, 2.969601, 2.989196, 2.988752, 3.010713, 3.000792, 
    3.037936, 3.027334, 3.05807, 3.050312, 3.057706, 3.055462, 3.057735, 
    3.046365, 3.051231, 3.041244, 3.002648, 3.013942, 2.98038, 2.960377, 
    2.947159, 2.937815, 2.939134, 2.941651, 2.954616, 2.966854, 2.976214, 
    2.982491, 2.988688, 3.007527, 3.017542, 3.040086, 3.036004, 3.042921, 
    3.049541, 3.060678, 3.058852, 3.063663, 3.042737, 3.056703, 3.033681, 
    3.039961, 2.990381, 2.971693, 2.963788, 2.956882, 2.940149, 2.951695, 
    2.947138, 2.957989, 2.964904, 2.961482, 2.982663, 2.974411, 3.018137, 
    2.999226, 3.048768, 3.036841, 3.051634, 3.044076, 3.057037, 3.04537, 
    3.065438, 3.069721, 3.066794, 3.078054, 3.044725, 3.057706, 2.961386, 
    2.961944, 2.964544, 2.953132, 2.952435, 2.942014, 2.951284, 2.95524, 
    2.965305, 2.971275, 2.97696, 2.989497, 3.00356, 3.023331, 3.037613, 
    3.047223, 3.041326, 3.046532, 3.040714, 3.03799, 3.068116, 3.051277, 
    3.076432, 3.07505, 3.063777, 3.075206, 2.962336, 2.959126, 2.948011, 
    2.956706, 2.940882, 2.94973, 2.95483, 2.974585, 2.97894, 2.982987, 
    2.990993, 3.001299, 3.019462, 3.035351, 3.049927, 3.048856, 3.049233, 
    3.052498, 3.044417, 3.053827, 3.05541, 3.051274, 3.074865, 3.068189, 
    3.075021, 3.070672, 2.960169, 2.965573, 2.962652, 2.968148, 2.964275, 
    2.981533, 2.986726, 3.011141, 3.001096, 3.017096, 3.002717, 3.00526, 
    3.017622, 3.003492, 3.034474, 3.013438, 3.052625, 3.031498, 3.053954, 
    3.049864, 3.056639, 3.062643, 3.070064, 3.083807, 3.080619, 3.092148, 
    2.973646, 2.980689, 2.980067, 2.987452, 2.992925, 3.00482, 3.023995, 
    3.01677, 3.030046, 3.032718, 3.012553, 3.02492, 2.98541, 2.99176, 
    2.987977, 2.974202, 3.018435, 2.995656, 3.03785, 3.025411, 3.061803, 
    3.043677, 3.078866, 3.093806, 3.10793, 3.124524, 2.984538, 2.979745, 
    2.988331, 3.000251, 3.01135, 3.026169, 3.027688, 3.030474, 3.0377, 
    3.043789, 3.031356, 3.045317, 2.993237, 3.02042, 2.977936, 2.990669, 
    2.999547, 2.995648, 3.015945, 3.020749, 3.040346, 3.030199, 3.090113, 
    3.063889, 3.137215, 3.116547, 2.978072, 2.984521, 3.00707, 2.99632, 
    3.02716, 3.034799, 3.041021, 3.048995, 3.049857, 3.054593, 3.046836, 
    3.054285, 3.0262, 3.038719, 3.004483, 3.012782, 3.008961, 3.004776, 
    3.01771, 3.031552, 3.031847, 3.036299, 3.048882, 3.027285, 3.093517, 
    3.052865, 2.991568, 3.004057, 3.005843, 3.000996, 3.034032, 3.022022, 
    3.054477, 3.045672, 3.060111, 3.052928, 3.051872, 3.042673, 3.03696, 
    3.022572, 3.010913, 3.001699, 3.003839, 3.013969, 3.0324, 3.049936, 
    3.046086, 3.059011, 3.024913, 3.039167, 3.033651, 3.048054, 3.016579, 
    3.043367, 3.009769, 3.0127, 3.021784, 3.040137, 3.04421, 3.048567, 
    3.045877, 3.032869, 3.030742, 3.021562, 3.019033, 3.012061, 3.006302, 
    3.011564, 3.0171, 3.032874, 3.047158, 3.062727, 3.066445, 3.084268, 
    3.069754, 3.093744, 3.073339, 3.108747, 3.044924, 3.072738, 3.022197, 
    3.027646, 3.037527, 3.060306, 3.047986, 3.062331, 3.030659, 3.01432, 
    3.010105, 3.002258, 3.010284, 3.00963, 3.017329, 3.014853, 3.033399, 
    3.023423, 3.051846, 3.062221, 3.090938, 3.108678, 3.12684, 3.134893, 
    3.137349, 3.138376,
  2.96992, 2.988319, 2.984731, 2.999652, 2.991363, 3.00115, 2.973638, 
    2.989053, 2.979201, 2.971569, 3.028873, 3.000319, 3.058882, 3.04041, 
    3.087076, 3.055999, 3.09339, 3.086172, 3.107955, 3.101695, 3.129773, 
    3.11085, 3.144451, 3.125239, 3.128236, 3.110228, 3.006037, 3.025301, 
    3.004901, 3.007638, 3.006409, 2.991534, 2.984074, 2.968518, 2.971334, 
    2.982763, 3.008869, 2.999974, 3.022449, 3.021939, 3.047201, 3.035779, 
    3.078629, 3.066374, 3.101956, 3.092959, 3.101532, 3.098929, 3.101567, 
    3.088385, 3.094024, 3.082456, 3.037914, 3.050922, 3.01233, 2.989418, 
    2.974312, 2.963651, 2.965156, 2.968026, 2.98283, 2.996829, 3.007552, 
    3.014751, 3.021866, 3.043532, 3.055073, 3.081116, 3.076394, 3.084398, 
    3.092066, 3.104996, 3.102863, 3.108577, 3.084185, 3.100369, 3.073709, 
    3.080972, 3.02381, 3.00237, 2.99332, 2.98542, 2.966313, 2.979493, 
    2.974289, 2.986686, 2.994597, 2.990681, 3.014949, 3.005486, 3.055759, 
    3.033978, 3.09117, 3.077362, 3.094491, 3.085735, 3.100757, 3.087234, 
    3.110706, 3.115848, 3.112333, 3.125859, 3.086486, 3.101533, 2.990571, 
    2.99121, 2.994185, 2.981134, 2.980338, 2.968441, 2.979023, 2.983544, 
    2.995056, 3.001892, 3.008407, 3.022794, 3.038964, 3.061753, 3.078255, 
    3.08938, 3.082552, 3.088579, 3.081843, 3.078691, 3.11392, 3.094077, 
    3.123909, 3.122248, 3.108713, 3.122436, 2.991658, 2.987987, 2.975285, 
    2.985219, 2.967149, 2.977248, 2.983075, 3.005684, 3.010679, 3.015321, 
    3.024513, 3.036362, 3.057287, 3.075639, 3.092512, 3.091272, 3.091708, 
    3.095493, 3.08613, 3.097034, 3.098869, 3.094074, 3.122026, 3.114008, 
    3.122213, 3.116989, 2.989179, 2.995363, 2.992019, 2.99831, 2.993877, 
    3.013652, 3.019612, 3.047694, 3.036129, 3.054559, 3.037994, 3.040921, 
    3.055165, 3.038886, 3.074625, 3.050341, 3.09564, 3.071185, 3.097181, 
    3.092439, 3.100295, 3.107352, 3.116259, 3.13278, 3.128944, 3.142823, 
    3.004609, 3.012683, 3.01197, 3.020446, 3.026733, 3.040414, 3.062519, 
    3.054183, 3.069507, 3.072595, 3.049322, 3.063586, 3.018101, 3.025394, 
    3.021049, 3.005246, 3.056103, 3.029872, 3.078529, 3.064153, 3.106345, 
    3.085273, 3.126835, 3.144822, 3.161329, 3.180762, 3.0171, 3.011601, 
    3.021455, 3.035156, 3.047935, 3.065028, 3.066783, 3.070001, 3.078356, 
    3.085402, 3.071021, 3.087172, 3.027092, 3.058392, 3.009526, 3.02414, 
    3.034346, 3.029863, 3.053231, 3.058772, 3.081417, 3.069684, 3.140372, 
    3.108848, 3.195661, 3.171414, 3.009683, 3.017081, 3.043005, 3.030636, 
    3.066173, 3.075, 3.082199, 3.091433, 3.092431, 3.097921, 3.088932, 
    3.097565, 3.065065, 3.079535, 3.040026, 3.049585, 3.045182, 3.040363, 
    3.055267, 3.071247, 3.071588, 3.076735, 3.091301, 3.066318, 3.144474, 
    3.095918, 3.025173, 3.039536, 3.041592, 3.036014, 3.074114, 3.060241, 
    3.097787, 3.087583, 3.104324, 3.095991, 3.094767, 3.08411, 3.0775, 
    3.060875, 3.047431, 3.036822, 3.039284, 3.050953, 3.072227, 3.092523, 
    3.088063, 3.103048, 3.063579, 3.080053, 3.073673, 3.090343, 3.053962, 
    3.084914, 3.046113, 3.04949, 3.059966, 3.081176, 3.08589, 3.090937, 
    3.087821, 3.07277, 3.070312, 3.059711, 3.056792, 3.048754, 3.04212, 
    3.048181, 3.054563, 3.072775, 3.089305, 3.107453, 3.111914, 3.133334, 
    3.115886, 3.144747, 3.120193, 3.162284, 3.086717, 3.11947, 3.060443, 
    3.066734, 3.078156, 3.104551, 3.090264, 3.106979, 3.070215, 3.051358, 
    3.0465, 3.037466, 3.046707, 3.045954, 3.054826, 3.051971, 3.073382, 
    3.061858, 3.094737, 3.106846, 3.141365, 3.162204, 3.183479, 3.192933, 
    3.195818, 3.197025,
  3.254737, 3.278214, 3.273626, 3.292734, 3.282109, 3.294657, 3.259472, 
    3.279153, 3.266564, 3.256837, 3.3299, 3.29359, 3.367675, 3.344384, 
    3.40347, 3.364032, 3.411527, 3.402317, 3.430173, 3.422149, 3.458259, 
    3.433888, 3.477261, 3.452407, 3.456274, 3.43309, 3.300935, 3.325425, 
    3.299475, 3.302993, 3.301413, 3.282329, 3.272787, 3.252954, 3.256538, 
    3.271112, 3.304577, 3.293148, 3.321856, 3.321218, 3.352931, 3.338563, 
    3.392715, 3.377157, 3.422483, 3.410977, 3.421941, 3.418609, 3.421985, 
    3.405139, 3.412338, 3.397584, 3.341246, 3.357622, 3.309032, 3.279619, 
    3.260331, 3.246767, 3.248678, 3.252328, 3.271198, 3.289113, 3.302883, 
    3.312152, 3.321126, 3.348311, 3.362862, 3.395878, 3.389873, 3.400056, 
    3.409836, 3.426378, 3.423645, 3.43097, 3.399785, 3.420452, 3.386461, 
    3.395695, 3.323559, 3.296224, 3.284615, 3.274507, 3.250149, 3.266937, 
    3.260301, 3.276125, 3.286251, 3.281236, 3.312406, 3.300226, 3.363728, 
    3.336303, 3.408693, 3.391104, 3.412934, 3.401761, 3.420948, 3.403671, 
    3.433704, 3.440311, 3.435794, 3.453207, 3.402718, 3.421942, 3.281096, 
    3.281913, 3.285723, 3.269032, 3.268015, 3.252856, 3.266338, 3.27211, 
    3.286839, 3.295609, 3.303983, 3.322288, 3.342566, 3.371306, 3.392239, 
    3.406408, 3.397706, 3.405386, 3.396803, 3.392793, 3.437833, 3.412405, 
    3.450692, 3.448552, 3.431145, 3.448793, 3.282487, 3.277789, 3.261571, 
    3.274251, 3.251212, 3.264074, 3.27151, 3.300481, 3.306906, 3.312885, 
    3.324439, 3.339296, 3.365659, 3.388914, 3.410406, 3.408823, 3.40938, 
    3.414215, 3.402264, 3.416184, 3.418532, 3.412401, 3.448265, 3.437946, 
    3.448506, 3.44178, 3.279314, 3.287233, 3.28295, 3.291012, 3.285329, 
    3.310735, 3.318309, 3.353553, 3.339003, 3.362213, 3.341346, 3.345027, 
    3.362978, 3.342467, 3.387626, 3.35689, 3.414403, 3.383258, 3.416373, 
    3.410313, 3.420356, 3.4294, 3.44084, 3.462145, 3.457189, 3.475149, 
    3.299099, 3.309487, 3.308569, 3.31935, 3.327218, 3.344388, 3.372275, 
    3.361737, 3.381129, 3.385048, 3.355605, 3.373627, 3.31642, 3.325542, 
    3.320105, 3.299917, 3.364163, 3.331152, 3.392587, 3.374345, 3.428108, 
    3.401172, 3.454467, 3.477742, 3.499917, 3.526191, 3.31517, 3.308093, 
    3.320613, 3.337782, 3.353856, 3.375453, 3.377676, 3.381756, 3.392366, 
    3.401337, 3.38305, 3.403592, 3.327668, 3.367056, 3.305423, 3.323972, 
    3.336765, 3.331141, 3.360537, 3.367536, 3.396261, 3.381354, 3.471971, 
    3.431318, 3.546055, 3.513531, 3.305624, 3.315145, 3.347648, 3.33211, 
    3.376903, 3.388102, 3.397256, 3.409029, 3.410303, 3.41732, 3.405836, 
    3.416864, 3.375499, 3.393867, 3.343901, 3.355936, 3.350389, 3.344325, 
    3.363107, 3.383337, 3.383769, 3.390306, 3.408861, 3.377086, 3.477291, 
    3.414758, 3.325265, 3.343285, 3.34587, 3.338859, 3.386976, 3.369393, 
    3.417148, 3.404116, 3.425517, 3.414851, 3.413287, 3.399691, 3.391278, 
    3.370196, 3.353222, 3.339874, 3.342968, 3.357662, 3.384581, 3.41042, 
    3.404728, 3.423882, 3.373617, 3.394526, 3.386416, 3.407636, 3.361459, 
    3.400715, 3.351561, 3.355817, 3.369046, 3.395954, 3.401958, 3.408395, 
    3.40442, 3.385269, 3.38215, 3.368722, 3.365034, 3.35489, 3.346535, 
    3.354167, 3.362218, 3.385276, 3.406312, 3.429529, 3.435256, 3.462861, 
    3.440361, 3.477646, 3.445904, 3.501205, 3.403012, 3.444973, 3.369649, 
    3.377614, 3.392113, 3.425807, 3.407536, 3.428921, 3.382027, 3.358173, 
    3.352048, 3.340683, 3.352309, 3.351361, 3.36255, 3.358947, 3.386047, 
    3.371439, 3.413249, 3.428751, 3.473259, 3.501097, 3.529877, 3.542453, 
    3.546262, 3.547857,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016906, 3.972589, 
    4.084889, 4.009922, 4.10039, 4.08268, 4.136661, 4.120983, 4.192374, 
    4.143956, 4.230834, 4.180657, 4.188393, 4.142387, 3.892786, 3.937095, 
    3.890204, 3.896427, 3.893631, 3.860096, 3.843496, 3.80934, 3.815479, 
    3.840593, 3.899234, 3.879051, 3.93047, 3.929288, 3.98876, 3.961638, 
    4.064354, 4.034962, 4.121634, 4.099329, 4.120579, 4.114101, 4.120664, 
    4.088092, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821991, 3.798779, 3.802037, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078352, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077834, 4.117682, 4.052496, 
    4.070027, 3.933629, 3.884468, 3.86409, 3.846481, 3.804548, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085274, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083447, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835236, 3.809173, 3.832339, 3.842322, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023888, 4.063449, 
    4.09053, 4.073862, 4.088567, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846035, 3.806363, 3.828434, 3.841284, 3.891984, 3.903367, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095176, 4.09625, 
    4.105584, 4.082578, 4.109397, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172877, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865338, 
    3.910178, 3.923903, 3.98994, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007905, 3.968978, 4.054699, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226528, 
    3.889541, 3.907957, 3.906323, 3.925829, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937313, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132616, 
    4.080487, 4.184773, 4.231818, 4.277537, 4.332245, 3.918106, 3.905478, 
    3.928166, 3.960172, 3.990517, 4.031764, 4.035936, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941267, 4.015718, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071106, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034484, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971678, 3.994471, 3.983939, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.095249, 4.034829, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975393, 3.962193, 4.05347, 4.020208, 
    4.111265, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021752, 3.989313, 3.964099, 3.969922, 3.997757, 4.048942, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.067799, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994244, 4.01954, 4.070521, 4.081992, 4.094354, 
    4.086711, 4.050242, 4.044355, 4.018919, 4.011841, 3.99248, 3.976649, 
    3.991108, 4.006452, 4.050255, 4.090346, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084011, 4.165854, 4.0207, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044124, 3.998729, 
    3.987085, 3.96562, 3.98758, 3.985781, 4.007087, 4.000206, 4.051712, 
    4.024145, 4.103716, 4.133875, 4.222682, 4.279995, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24814.02, 24834.45, 24830.45, 24847.17, 24837.86, 24848.86, 24818.13, 
    24835.27, 24824.29, 24815.84, 24880.38, 24847.92, 24915.13, 24893.65, 
    24948.09, 24911.76, 24955.55, 24947.02, 24972.93, 24965.44, 24999.37, 
    24976.41, 25017.45, 24993.83, 24997.49, 24975.66, 24854.38, 24876.3, 
    24853.1, 24856.2, 24854.8, 24838.05, 24829.71, 24812.47, 24815.58, 
    24828.25, 24857.59, 24847.53, 24873.05, 24872.47, 24901.51, 24888.31, 
    24938.16, 24923.88, 24965.75, 24955.04, 24965.25, 24962.14, 24965.29, 
    24949.63, 24956.31, 24942.65, 24890.77, 24905.84, 24861.53, 24835.68, 
    24818.87, 24807.12, 24808.77, 24811.93, 24828.33, 24843.99, 24856.1, 
    24864.29, 24872.38, 24897.26, 24910.68, 24941.07, 24935.54, 24944.93, 
    24953.98, 24969.39, 24966.84, 24973.68, 24944.68, 24963.86, 24932.41, 
    24940.91, 24874.6, 24850.24, 24840.05, 24831.21, 24810.04, 24824.62, 
    24818.85, 24832.62, 24841.48, 24837.09, 24864.51, 24853.76, 24911.48, 
    24886.24, 24952.92, 24936.68, 24956.86, 24946.51, 24964.32, 24948.27, 
    24976.24, 24982.44, 24978.2, 24994.59, 24947.39, 24965.25, 24836.97, 
    24837.69, 24841.02, 24826.44, 24825.55, 24812.39, 24824.09, 24829.12, 
    24842, 24849.7, 24857.07, 24873.44, 24891.98, 24918.5, 24937.72, 
    24950.81, 24942.76, 24949.86, 24941.93, 24938.23, 24980.11, 24956.37, 
    24992.21, 24990.19, 24973.84, 24990.42, 24838.19, 24834.08, 24819.95, 
    24830.99, 24810.96, 24822.12, 24828.6, 24853.98, 24859.65, 24864.93, 
    24875.4, 24888.98, 24913.27, 24934.66, 24954.51, 24953.04, 24953.56, 
    24958.05, 24946.97, 24959.88, 24962.07, 24956.37, 24989.92, 24980.21, 
    24990.15, 24983.81, 24835.41, 24842.34, 24838.59, 24845.66, 24840.68, 
    24863.03, 24869.82, 24902.08, 24888.71, 24910.08, 24890.86, 24894.24, 
    24910.79, 24891.89, 24933.48, 24905.16, 24958.23, 24929.47, 24960.06, 
    24954.43, 24963.77, 24972.21, 24982.93, 25003.05, 24998.35, 25015.43, 
    24852.77, 24861.93, 24861.12, 24870.77, 24877.94, 24893.65, 24919.4, 
    24909.64, 24927.52, 24931.11, 24903.97, 24920.65, 24868.1, 24876.41, 
    24871.45, 24853.49, 24911.88, 24881.53, 24938.04, 24921.31, 24971, 
    24945.96, 24995.78, 25017.91, 25039.19, 25064.53, 24866.96, 24860.7, 
    24871.92, 24887.59, 24902.36, 24922.32, 24924.36, 24928.09, 24937.84, 
    24946.12, 24929.28, 24948.2, 24878.35, 24914.56, 24858.34, 24874.98, 
    24886.66, 24881.52, 24908.53, 24915.01, 24941.43, 24927.72, 25012.4, 
    24974, 25084.04, 25052.37, 24858.52, 24866.94, 24896.65, 24882.4, 
    24923.65, 24933.92, 24942.35, 24953.24, 24954.42, 24960.94, 24950.28, 
    24960.52, 24922.37, 24939.22, 24893.21, 24904.28, 24899.17, 24893.6, 
    24910.9, 24929.54, 24929.94, 24935.94, 24953.08, 24923.82, 25017.48, 
    24958.56, 24876.16, 24892.64, 24895.02, 24888.58, 24932.88, 24916.73, 
    24960.78, 24948.68, 24968.58, 24958.64, 24957.19, 24944.59, 24936.84, 
    24917.47, 24901.78, 24889.51, 24892.35, 24905.87, 24930.68, 24954.53, 
    24949.25, 24967.06, 24920.65, 24939.83, 24932.37, 24951.95, 24909.38, 
    24945.54, 24900.25, 24904.17, 24916.41, 24941.14, 24946.69, 24952.65, 
    24948.97, 24931.31, 24928.45, 24916.11, 24912.69, 24903.32, 24895.63, 
    24902.65, 24910.08, 24931.32, 24950.72, 24972.33, 24977.69, 25003.73, 
    24982.48, 25017.82, 24987.7, 25040.43, 24947.66, 24986.82, 24916.97, 
    24924.3, 24937.61, 24968.86, 24951.85, 24971.76, 24928.34, 24906.34, 
    24900.7, 24890.25, 24900.94, 24900.06, 24910.39, 24907.06, 24932.03, 
    24918.63, 24957.15, 24971.6, 25013.63, 25040.33, 25068.08, 25080.45, 
    25084.25, 25085.84 ;

 HCSOI =
  24814.02, 24834.45, 24830.45, 24847.17, 24837.86, 24848.86, 24818.13, 
    24835.27, 24824.29, 24815.84, 24880.38, 24847.92, 24915.13, 24893.65, 
    24948.09, 24911.76, 24955.55, 24947.02, 24972.93, 24965.44, 24999.37, 
    24976.41, 25017.45, 24993.83, 24997.49, 24975.66, 24854.38, 24876.3, 
    24853.1, 24856.2, 24854.8, 24838.05, 24829.71, 24812.47, 24815.58, 
    24828.25, 24857.59, 24847.53, 24873.05, 24872.47, 24901.51, 24888.31, 
    24938.16, 24923.88, 24965.75, 24955.04, 24965.25, 24962.14, 24965.29, 
    24949.63, 24956.31, 24942.65, 24890.77, 24905.84, 24861.53, 24835.68, 
    24818.87, 24807.12, 24808.77, 24811.93, 24828.33, 24843.99, 24856.1, 
    24864.29, 24872.38, 24897.26, 24910.68, 24941.07, 24935.54, 24944.93, 
    24953.98, 24969.39, 24966.84, 24973.68, 24944.68, 24963.86, 24932.41, 
    24940.91, 24874.6, 24850.24, 24840.05, 24831.21, 24810.04, 24824.62, 
    24818.85, 24832.62, 24841.48, 24837.09, 24864.51, 24853.76, 24911.48, 
    24886.24, 24952.92, 24936.68, 24956.86, 24946.51, 24964.32, 24948.27, 
    24976.24, 24982.44, 24978.2, 24994.59, 24947.39, 24965.25, 24836.97, 
    24837.69, 24841.02, 24826.44, 24825.55, 24812.39, 24824.09, 24829.12, 
    24842, 24849.7, 24857.07, 24873.44, 24891.98, 24918.5, 24937.72, 
    24950.81, 24942.76, 24949.86, 24941.93, 24938.23, 24980.11, 24956.37, 
    24992.21, 24990.19, 24973.84, 24990.42, 24838.19, 24834.08, 24819.95, 
    24830.99, 24810.96, 24822.12, 24828.6, 24853.98, 24859.65, 24864.93, 
    24875.4, 24888.98, 24913.27, 24934.66, 24954.51, 24953.04, 24953.56, 
    24958.05, 24946.97, 24959.88, 24962.07, 24956.37, 24989.92, 24980.21, 
    24990.15, 24983.81, 24835.41, 24842.34, 24838.59, 24845.66, 24840.68, 
    24863.03, 24869.82, 24902.08, 24888.71, 24910.08, 24890.86, 24894.24, 
    24910.79, 24891.89, 24933.48, 24905.16, 24958.23, 24929.47, 24960.06, 
    24954.43, 24963.77, 24972.21, 24982.93, 25003.05, 24998.35, 25015.43, 
    24852.77, 24861.93, 24861.12, 24870.77, 24877.94, 24893.65, 24919.4, 
    24909.64, 24927.52, 24931.11, 24903.97, 24920.65, 24868.1, 24876.41, 
    24871.45, 24853.49, 24911.88, 24881.53, 24938.04, 24921.31, 24971, 
    24945.96, 24995.78, 25017.91, 25039.19, 25064.53, 24866.96, 24860.7, 
    24871.92, 24887.59, 24902.36, 24922.32, 24924.36, 24928.09, 24937.84, 
    24946.12, 24929.28, 24948.2, 24878.35, 24914.56, 24858.34, 24874.98, 
    24886.66, 24881.52, 24908.53, 24915.01, 24941.43, 24927.72, 25012.4, 
    24974, 25084.04, 25052.37, 24858.52, 24866.94, 24896.65, 24882.4, 
    24923.65, 24933.92, 24942.35, 24953.24, 24954.42, 24960.94, 24950.28, 
    24960.52, 24922.37, 24939.22, 24893.21, 24904.28, 24899.17, 24893.6, 
    24910.9, 24929.54, 24929.94, 24935.94, 24953.08, 24923.82, 25017.48, 
    24958.56, 24876.16, 24892.64, 24895.02, 24888.58, 24932.88, 24916.73, 
    24960.78, 24948.68, 24968.58, 24958.64, 24957.19, 24944.59, 24936.84, 
    24917.47, 24901.78, 24889.51, 24892.35, 24905.87, 24930.68, 24954.53, 
    24949.25, 24967.06, 24920.65, 24939.83, 24932.37, 24951.95, 24909.38, 
    24945.54, 24900.25, 24904.17, 24916.41, 24941.14, 24946.69, 24952.65, 
    24948.97, 24931.31, 24928.45, 24916.11, 24912.69, 24903.32, 24895.63, 
    24902.65, 24910.08, 24931.32, 24950.72, 24972.33, 24977.69, 25003.73, 
    24982.48, 25017.82, 24987.7, 25040.43, 24947.66, 24986.82, 24916.97, 
    24924.3, 24937.61, 24968.86, 24951.85, 24971.76, 24928.34, 24906.34, 
    24900.7, 24890.25, 24900.94, 24900.06, 24910.39, 24907.06, 24932.03, 
    24918.63, 24957.15, 24971.6, 25013.63, 25040.33, 25068.08, 25080.45, 
    25084.25, 25085.84 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.35703e-08, 6.384985e-08, 6.379551e-08, 6.402099e-08, 6.389591e-08, 
    6.404356e-08, 6.362697e-08, 6.386096e-08, 6.371158e-08, 6.359546e-08, 
    6.445858e-08, 6.403105e-08, 6.490264e-08, 6.462999e-08, 6.531489e-08, 
    6.486022e-08, 6.540657e-08, 6.530176e-08, 6.561717e-08, 6.552681e-08, 
    6.593026e-08, 6.565888e-08, 6.613939e-08, 6.586544e-08, 6.59083e-08, 
    6.564993e-08, 6.411708e-08, 6.440536e-08, 6.410001e-08, 6.414111e-08, 
    6.412267e-08, 6.38985e-08, 6.378554e-08, 6.354892e-08, 6.359188e-08, 
    6.376565e-08, 6.41596e-08, 6.402587e-08, 6.436288e-08, 6.435527e-08, 
    6.473046e-08, 6.45613e-08, 6.519191e-08, 6.501268e-08, 6.553059e-08, 
    6.540034e-08, 6.552447e-08, 6.548683e-08, 6.552496e-08, 6.533394e-08, 
    6.541578e-08, 6.524769e-08, 6.459298e-08, 6.47854e-08, 6.421152e-08, 
    6.386645e-08, 6.363724e-08, 6.347459e-08, 6.349758e-08, 6.354141e-08, 
    6.376668e-08, 6.397845e-08, 6.413985e-08, 6.424781e-08, 6.435418e-08, 
    6.467617e-08, 6.484658e-08, 6.522815e-08, 6.515928e-08, 6.527594e-08, 
    6.538738e-08, 6.557449e-08, 6.554369e-08, 6.562612e-08, 6.527286e-08, 
    6.550764e-08, 6.512006e-08, 6.522607e-08, 6.438312e-08, 6.406194e-08, 
    6.392545e-08, 6.380596e-08, 6.351526e-08, 6.371601e-08, 6.363688e-08, 
    6.382514e-08, 6.394477e-08, 6.38856e-08, 6.425076e-08, 6.41088e-08, 
    6.485669e-08, 6.453455e-08, 6.537438e-08, 6.517342e-08, 6.542255e-08, 
    6.529542e-08, 6.551326e-08, 6.531721e-08, 6.565681e-08, 6.573075e-08, 
    6.568022e-08, 6.587433e-08, 6.530634e-08, 6.552447e-08, 6.388395e-08, 
    6.389359e-08, 6.393855e-08, 6.374094e-08, 6.372885e-08, 6.354775e-08, 
    6.370889e-08, 6.377751e-08, 6.39517e-08, 6.405474e-08, 6.415268e-08, 
    6.436803e-08, 6.460854e-08, 6.494484e-08, 6.518644e-08, 6.53484e-08, 
    6.524908e-08, 6.533676e-08, 6.523875e-08, 6.519281e-08, 6.570305e-08, 
    6.541654e-08, 6.584641e-08, 6.582263e-08, 6.562809e-08, 6.58253e-08, 
    6.390037e-08, 6.384484e-08, 6.365205e-08, 6.380292e-08, 6.352803e-08, 
    6.36819e-08, 6.377039e-08, 6.411177e-08, 6.418676e-08, 6.425632e-08, 
    6.439367e-08, 6.456996e-08, 6.48792e-08, 6.514825e-08, 6.539386e-08, 
    6.537586e-08, 6.53822e-08, 6.543707e-08, 6.530116e-08, 6.545939e-08, 
    6.548594e-08, 6.541651e-08, 6.581944e-08, 6.570433e-08, 6.582212e-08, 
    6.574717e-08, 6.386289e-08, 6.395633e-08, 6.390584e-08, 6.400078e-08, 
    6.39339e-08, 6.423132e-08, 6.432049e-08, 6.473773e-08, 6.456649e-08, 
    6.483902e-08, 6.459417e-08, 6.463756e-08, 6.484792e-08, 6.46074e-08, 
    6.513343e-08, 6.477681e-08, 6.543921e-08, 6.508311e-08, 6.546152e-08, 
    6.53928e-08, 6.550658e-08, 6.560848e-08, 6.573668e-08, 6.597322e-08, 
    6.591844e-08, 6.611626e-08, 6.409562e-08, 6.421681e-08, 6.420614e-08, 
    6.433297e-08, 6.442676e-08, 6.463005e-08, 6.49561e-08, 6.483349e-08, 
    6.505858e-08, 6.510377e-08, 6.47618e-08, 6.497177e-08, 6.429792e-08, 
    6.44068e-08, 6.434197e-08, 6.410518e-08, 6.486175e-08, 6.447348e-08, 
    6.519043e-08, 6.498011e-08, 6.559395e-08, 6.528868e-08, 6.588829e-08, 
    6.614464e-08, 6.638587e-08, 6.66678e-08, 6.428295e-08, 6.42006e-08, 
    6.434804e-08, 6.455205e-08, 6.474131e-08, 6.499293e-08, 6.501867e-08, 
    6.506582e-08, 6.518791e-08, 6.529058e-08, 6.508073e-08, 6.531631e-08, 
    6.443206e-08, 6.489545e-08, 6.416948e-08, 6.438809e-08, 6.454002e-08, 
    6.447337e-08, 6.481947e-08, 6.490105e-08, 6.523254e-08, 6.506118e-08, 
    6.608137e-08, 6.563001e-08, 6.688245e-08, 6.653246e-08, 6.417183e-08, 
    6.428267e-08, 6.466841e-08, 6.448487e-08, 6.500973e-08, 6.513893e-08, 
    6.524394e-08, 6.53782e-08, 6.539269e-08, 6.547224e-08, 6.534189e-08, 
    6.546708e-08, 6.499347e-08, 6.520511e-08, 6.462431e-08, 6.476568e-08, 
    6.470064e-08, 6.46293e-08, 6.484947e-08, 6.508403e-08, 6.508903e-08, 
    6.516425e-08, 6.537621e-08, 6.501185e-08, 6.613964e-08, 6.544317e-08, 
    6.440352e-08, 6.461701e-08, 6.464749e-08, 6.456479e-08, 6.512597e-08, 
    6.492264e-08, 6.54703e-08, 6.532228e-08, 6.55648e-08, 6.544429e-08, 
    6.542655e-08, 6.527178e-08, 6.517542e-08, 6.493197e-08, 6.473388e-08, 
    6.457679e-08, 6.461332e-08, 6.478587e-08, 6.509838e-08, 6.5394e-08, 
    6.532925e-08, 6.554637e-08, 6.497167e-08, 6.521266e-08, 6.511952e-08, 
    6.536237e-08, 6.483023e-08, 6.528341e-08, 6.471441e-08, 6.476429e-08, 
    6.49186e-08, 6.522901e-08, 6.529767e-08, 6.5371e-08, 6.532575e-08, 
    6.510631e-08, 6.507035e-08, 6.491485e-08, 6.487192e-08, 6.475343e-08, 
    6.465533e-08, 6.474496e-08, 6.483909e-08, 6.51064e-08, 6.534729e-08, 
    6.560993e-08, 6.56742e-08, 6.598109e-08, 6.573129e-08, 6.614352e-08, 
    6.579306e-08, 6.639972e-08, 6.530966e-08, 6.578274e-08, 6.492562e-08, 
    6.501796e-08, 6.518498e-08, 6.556804e-08, 6.536123e-08, 6.560308e-08, 
    6.506895e-08, 6.479183e-08, 6.472012e-08, 6.458635e-08, 6.472317e-08, 
    6.471205e-08, 6.484298e-08, 6.480091e-08, 6.511527e-08, 6.494641e-08, 
    6.542611e-08, 6.560117e-08, 6.609553e-08, 6.639859e-08, 6.670707e-08, 
    6.684326e-08, 6.688472e-08, 6.690204e-08 ;

 HR_vr =
  2.667178e-07, 2.67426e-07, 2.672884e-07, 2.678591e-07, 2.675426e-07, 
    2.679162e-07, 2.668614e-07, 2.674541e-07, 2.670758e-07, 2.667815e-07, 
    2.689654e-07, 2.678846e-07, 2.700857e-07, 2.69398e-07, 2.711239e-07, 
    2.699788e-07, 2.713545e-07, 2.710908e-07, 2.71884e-07, 2.716569e-07, 
    2.726703e-07, 2.719888e-07, 2.731948e-07, 2.725075e-07, 2.726152e-07, 
    2.719663e-07, 2.681022e-07, 2.688309e-07, 2.68059e-07, 2.68163e-07, 
    2.681163e-07, 2.675491e-07, 2.672631e-07, 2.666636e-07, 2.667725e-07, 
    2.672128e-07, 2.682097e-07, 2.678715e-07, 2.687235e-07, 2.687043e-07, 
    2.696515e-07, 2.692246e-07, 2.708143e-07, 2.70363e-07, 2.716664e-07, 
    2.713388e-07, 2.71651e-07, 2.715563e-07, 2.716522e-07, 2.711718e-07, 
    2.713777e-07, 2.709547e-07, 2.693046e-07, 2.697901e-07, 2.68341e-07, 
    2.67468e-07, 2.668874e-07, 2.664751e-07, 2.665334e-07, 2.666446e-07, 
    2.672153e-07, 2.677515e-07, 2.681597e-07, 2.684327e-07, 2.687015e-07, 
    2.695146e-07, 2.699444e-07, 2.709056e-07, 2.707322e-07, 2.710258e-07, 
    2.713062e-07, 2.717767e-07, 2.716993e-07, 2.719065e-07, 2.710181e-07, 
    2.716087e-07, 2.706334e-07, 2.709003e-07, 2.687748e-07, 2.679627e-07, 
    2.676174e-07, 2.673148e-07, 2.665783e-07, 2.67087e-07, 2.668865e-07, 
    2.673634e-07, 2.676662e-07, 2.675165e-07, 2.684401e-07, 2.680812e-07, 
    2.699698e-07, 2.691571e-07, 2.712735e-07, 2.707677e-07, 2.713947e-07, 
    2.710748e-07, 2.716228e-07, 2.711297e-07, 2.719836e-07, 2.721694e-07, 
    2.720424e-07, 2.725299e-07, 2.711023e-07, 2.71651e-07, 2.675123e-07, 
    2.675367e-07, 2.676505e-07, 2.671502e-07, 2.671195e-07, 2.666606e-07, 
    2.67069e-07, 2.672428e-07, 2.676838e-07, 2.679445e-07, 2.681922e-07, 
    2.687365e-07, 2.693439e-07, 2.701921e-07, 2.708005e-07, 2.712081e-07, 
    2.709582e-07, 2.711789e-07, 2.709322e-07, 2.708166e-07, 2.720998e-07, 
    2.713796e-07, 2.724598e-07, 2.724e-07, 2.719114e-07, 2.724068e-07, 
    2.675538e-07, 2.674133e-07, 2.66925e-07, 2.673071e-07, 2.666106e-07, 
    2.670006e-07, 2.672247e-07, 2.680888e-07, 2.682784e-07, 2.684542e-07, 
    2.688013e-07, 2.692465e-07, 2.700266e-07, 2.707044e-07, 2.713225e-07, 
    2.712773e-07, 2.712932e-07, 2.714312e-07, 2.710893e-07, 2.714873e-07, 
    2.715541e-07, 2.713795e-07, 2.72392e-07, 2.721029e-07, 2.723988e-07, 
    2.722105e-07, 2.674589e-07, 2.676955e-07, 2.675677e-07, 2.67808e-07, 
    2.676387e-07, 2.683911e-07, 2.686164e-07, 2.696699e-07, 2.692377e-07, 
    2.699253e-07, 2.693076e-07, 2.694171e-07, 2.699478e-07, 2.69341e-07, 
    2.706672e-07, 2.697684e-07, 2.714366e-07, 2.705404e-07, 2.714927e-07, 
    2.713199e-07, 2.71606e-07, 2.718621e-07, 2.721842e-07, 2.72778e-07, 
    2.726406e-07, 2.731368e-07, 2.680479e-07, 2.683544e-07, 2.683274e-07, 
    2.686479e-07, 2.688849e-07, 2.693981e-07, 2.702204e-07, 2.699113e-07, 
    2.704786e-07, 2.705924e-07, 2.697305e-07, 2.702599e-07, 2.685594e-07, 
    2.688345e-07, 2.686707e-07, 2.680721e-07, 2.699826e-07, 2.690029e-07, 
    2.708106e-07, 2.702809e-07, 2.718256e-07, 2.710579e-07, 2.725649e-07, 
    2.73208e-07, 2.738124e-07, 2.745181e-07, 2.685215e-07, 2.683134e-07, 
    2.68686e-07, 2.692013e-07, 2.696788e-07, 2.703132e-07, 2.703781e-07, 
    2.704968e-07, 2.708042e-07, 2.710626e-07, 2.705344e-07, 2.711274e-07, 
    2.688983e-07, 2.700675e-07, 2.682347e-07, 2.687873e-07, 2.691709e-07, 
    2.690026e-07, 2.69876e-07, 2.700816e-07, 2.709166e-07, 2.704851e-07, 
    2.730494e-07, 2.719163e-07, 2.750547e-07, 2.741795e-07, 2.682406e-07, 
    2.685208e-07, 2.694949e-07, 2.690316e-07, 2.703555e-07, 2.70681e-07, 
    2.709453e-07, 2.712831e-07, 2.713196e-07, 2.715196e-07, 2.711918e-07, 
    2.715067e-07, 2.703146e-07, 2.708476e-07, 2.693836e-07, 2.697403e-07, 
    2.695762e-07, 2.693963e-07, 2.699516e-07, 2.705428e-07, 2.705553e-07, 
    2.707447e-07, 2.712783e-07, 2.703609e-07, 2.731956e-07, 2.714466e-07, 
    2.688262e-07, 2.693653e-07, 2.694422e-07, 2.692334e-07, 2.706483e-07, 
    2.701361e-07, 2.715148e-07, 2.711424e-07, 2.717523e-07, 2.714494e-07, 
    2.714048e-07, 2.710154e-07, 2.707728e-07, 2.701596e-07, 2.696601e-07, 
    2.692637e-07, 2.693559e-07, 2.697913e-07, 2.705789e-07, 2.713229e-07, 
    2.7116e-07, 2.71706e-07, 2.702596e-07, 2.708666e-07, 2.706321e-07, 
    2.712433e-07, 2.699031e-07, 2.710447e-07, 2.69611e-07, 2.697368e-07, 
    2.701259e-07, 2.709077e-07, 2.710805e-07, 2.71265e-07, 2.711512e-07, 
    2.705988e-07, 2.705083e-07, 2.701164e-07, 2.700082e-07, 2.697094e-07, 
    2.694619e-07, 2.696881e-07, 2.699254e-07, 2.705991e-07, 2.712054e-07, 
    2.718658e-07, 2.720273e-07, 2.727978e-07, 2.721707e-07, 2.732053e-07, 
    2.723259e-07, 2.738472e-07, 2.711107e-07, 2.723e-07, 2.701436e-07, 
    2.703763e-07, 2.707969e-07, 2.717605e-07, 2.712404e-07, 2.718486e-07, 
    2.705047e-07, 2.698063e-07, 2.696254e-07, 2.692878e-07, 2.696331e-07, 
    2.69605e-07, 2.699352e-07, 2.698291e-07, 2.706214e-07, 2.70196e-07, 
    2.714036e-07, 2.718438e-07, 2.730849e-07, 2.738443e-07, 2.746163e-07, 
    2.749568e-07, 2.750604e-07, 2.751036e-07,
  2.414499e-07, 2.423604e-07, 2.421834e-07, 2.429173e-07, 2.425103e-07, 
    2.429907e-07, 2.416346e-07, 2.423965e-07, 2.419102e-07, 2.415319e-07, 
    2.443397e-07, 2.4295e-07, 2.457811e-07, 2.448964e-07, 2.47117e-07, 
    2.456434e-07, 2.474139e-07, 2.470746e-07, 2.480955e-07, 2.478031e-07, 
    2.491075e-07, 2.482304e-07, 2.49783e-07, 2.488981e-07, 2.490366e-07, 
    2.482014e-07, 2.432299e-07, 2.441668e-07, 2.431743e-07, 2.43308e-07, 
    2.43248e-07, 2.425187e-07, 2.421509e-07, 2.413803e-07, 2.415202e-07, 
    2.420862e-07, 2.433681e-07, 2.429332e-07, 2.440289e-07, 2.440042e-07, 
    2.452226e-07, 2.446734e-07, 2.467187e-07, 2.461379e-07, 2.478153e-07, 
    2.473938e-07, 2.477955e-07, 2.476737e-07, 2.477971e-07, 2.471788e-07, 
    2.474438e-07, 2.468994e-07, 2.447763e-07, 2.454008e-07, 2.435369e-07, 
    2.424143e-07, 2.41668e-07, 2.41138e-07, 2.41213e-07, 2.413558e-07, 
    2.420896e-07, 2.427789e-07, 2.433039e-07, 2.436549e-07, 2.440006e-07, 
    2.450462e-07, 2.455992e-07, 2.468361e-07, 2.46613e-07, 2.469909e-07, 
    2.473518e-07, 2.479574e-07, 2.478577e-07, 2.481244e-07, 2.46981e-07, 
    2.47741e-07, 2.46486e-07, 2.468294e-07, 2.440945e-07, 2.430505e-07, 
    2.426063e-07, 2.422175e-07, 2.412706e-07, 2.419246e-07, 2.416668e-07, 
    2.422799e-07, 2.426693e-07, 2.424767e-07, 2.436645e-07, 2.432029e-07, 
    2.45632e-07, 2.445865e-07, 2.473097e-07, 2.466588e-07, 2.474657e-07, 
    2.470541e-07, 2.477592e-07, 2.471246e-07, 2.482236e-07, 2.484628e-07, 
    2.482994e-07, 2.489269e-07, 2.470894e-07, 2.477955e-07, 2.424713e-07, 
    2.425028e-07, 2.426491e-07, 2.420057e-07, 2.419664e-07, 2.413765e-07, 
    2.419014e-07, 2.421249e-07, 2.426919e-07, 2.430271e-07, 2.433456e-07, 
    2.440457e-07, 2.448268e-07, 2.45918e-07, 2.46701e-07, 2.472256e-07, 
    2.46904e-07, 2.471879e-07, 2.468705e-07, 2.467217e-07, 2.483731e-07, 
    2.474462e-07, 2.488366e-07, 2.487598e-07, 2.481307e-07, 2.487684e-07, 
    2.425248e-07, 2.423441e-07, 2.417162e-07, 2.422076e-07, 2.413122e-07, 
    2.418135e-07, 2.421016e-07, 2.432126e-07, 2.434565e-07, 2.436826e-07, 
    2.44129e-07, 2.447015e-07, 2.457051e-07, 2.465773e-07, 2.473728e-07, 
    2.473145e-07, 2.473351e-07, 2.475127e-07, 2.470726e-07, 2.475849e-07, 
    2.476708e-07, 2.474461e-07, 2.487495e-07, 2.483773e-07, 2.487581e-07, 
    2.485158e-07, 2.424028e-07, 2.427069e-07, 2.425426e-07, 2.428515e-07, 
    2.426339e-07, 2.436012e-07, 2.438911e-07, 2.452461e-07, 2.446903e-07, 
    2.455747e-07, 2.447802e-07, 2.44921e-07, 2.456035e-07, 2.448231e-07, 
    2.465292e-07, 2.453729e-07, 2.475196e-07, 2.463661e-07, 2.475918e-07, 
    2.473694e-07, 2.477377e-07, 2.480673e-07, 2.484819e-07, 2.492464e-07, 
    2.490694e-07, 2.497083e-07, 2.431601e-07, 2.435541e-07, 2.435195e-07, 
    2.439317e-07, 2.442364e-07, 2.448967e-07, 2.459545e-07, 2.455569e-07, 
    2.462867e-07, 2.464332e-07, 2.453243e-07, 2.460053e-07, 2.438178e-07, 
    2.441715e-07, 2.43961e-07, 2.431912e-07, 2.456485e-07, 2.443882e-07, 
    2.46714e-07, 2.460323e-07, 2.480203e-07, 2.470322e-07, 2.48972e-07, 
    2.497999e-07, 2.505784e-07, 2.514871e-07, 2.437691e-07, 2.435015e-07, 
    2.439807e-07, 2.446433e-07, 2.452578e-07, 2.460739e-07, 2.461574e-07, 
    2.463102e-07, 2.467058e-07, 2.470384e-07, 2.463585e-07, 2.471217e-07, 
    2.442535e-07, 2.457578e-07, 2.434002e-07, 2.441108e-07, 2.446043e-07, 
    2.443878e-07, 2.455114e-07, 2.45776e-07, 2.468504e-07, 2.462952e-07, 
    2.495956e-07, 2.481369e-07, 2.521785e-07, 2.51051e-07, 2.434079e-07, 
    2.437682e-07, 2.450211e-07, 2.444252e-07, 2.461284e-07, 2.465471e-07, 
    2.468873e-07, 2.473221e-07, 2.47369e-07, 2.476265e-07, 2.472045e-07, 
    2.476098e-07, 2.460756e-07, 2.467615e-07, 2.44878e-07, 2.453368e-07, 
    2.451258e-07, 2.448942e-07, 2.456087e-07, 2.463692e-07, 2.463854e-07, 
    2.466291e-07, 2.473154e-07, 2.461353e-07, 2.497836e-07, 2.475322e-07, 
    2.44161e-07, 2.448542e-07, 2.449533e-07, 2.446848e-07, 2.465051e-07, 
    2.45846e-07, 2.476202e-07, 2.471411e-07, 2.47926e-07, 2.47536e-07, 
    2.474787e-07, 2.469775e-07, 2.466653e-07, 2.458762e-07, 2.452336e-07, 
    2.447237e-07, 2.448423e-07, 2.454023e-07, 2.464157e-07, 2.473732e-07, 
    2.471636e-07, 2.478664e-07, 2.46005e-07, 2.46786e-07, 2.464842e-07, 
    2.472709e-07, 2.455463e-07, 2.47015e-07, 2.451705e-07, 2.453323e-07, 
    2.458329e-07, 2.468389e-07, 2.470613e-07, 2.472987e-07, 2.471523e-07, 
    2.464414e-07, 2.463249e-07, 2.458207e-07, 2.456815e-07, 2.452971e-07, 
    2.449787e-07, 2.452696e-07, 2.45575e-07, 2.464417e-07, 2.47222e-07, 
    2.48072e-07, 2.482799e-07, 2.492717e-07, 2.484644e-07, 2.497961e-07, 
    2.48664e-07, 2.506229e-07, 2.471e-07, 2.486307e-07, 2.458557e-07, 
    2.461551e-07, 2.466963e-07, 2.479364e-07, 2.472671e-07, 2.480498e-07, 
    2.463203e-07, 2.454216e-07, 2.45189e-07, 2.447547e-07, 2.451989e-07, 
    2.451628e-07, 2.455876e-07, 2.454511e-07, 2.464705e-07, 2.459231e-07, 
    2.474772e-07, 2.480436e-07, 2.496414e-07, 2.506193e-07, 2.516137e-07, 
    2.520523e-07, 2.521858e-07, 2.522416e-07,
  2.259464e-07, 2.269437e-07, 2.267498e-07, 2.275538e-07, 2.271079e-07, 
    2.276343e-07, 2.261486e-07, 2.269832e-07, 2.264505e-07, 2.260362e-07, 
    2.291128e-07, 2.275897e-07, 2.306933e-07, 2.297232e-07, 2.321591e-07, 
    2.305424e-07, 2.324848e-07, 2.321125e-07, 2.332329e-07, 2.32912e-07, 
    2.343441e-07, 2.33381e-07, 2.350859e-07, 2.341142e-07, 2.342663e-07, 
    2.333492e-07, 2.278964e-07, 2.289232e-07, 2.278355e-07, 2.27982e-07, 
    2.279162e-07, 2.271171e-07, 2.267142e-07, 2.258701e-07, 2.260234e-07, 
    2.266433e-07, 2.280478e-07, 2.275712e-07, 2.287721e-07, 2.28745e-07, 
    2.300808e-07, 2.294787e-07, 2.31722e-07, 2.310848e-07, 2.329254e-07, 
    2.324628e-07, 2.329037e-07, 2.3277e-07, 2.329054e-07, 2.322268e-07, 
    2.325176e-07, 2.319203e-07, 2.295915e-07, 2.302763e-07, 2.282329e-07, 
    2.270027e-07, 2.261852e-07, 2.256048e-07, 2.256869e-07, 2.258433e-07, 
    2.26647e-07, 2.274022e-07, 2.279775e-07, 2.283622e-07, 2.287411e-07, 
    2.298875e-07, 2.304939e-07, 2.318508e-07, 2.316061e-07, 2.320207e-07, 
    2.324167e-07, 2.330813e-07, 2.32972e-07, 2.332647e-07, 2.320098e-07, 
    2.328439e-07, 2.314666e-07, 2.318434e-07, 2.28844e-07, 2.276998e-07, 
    2.272131e-07, 2.267871e-07, 2.2575e-07, 2.264663e-07, 2.261839e-07, 
    2.268555e-07, 2.272821e-07, 2.270712e-07, 2.283727e-07, 2.278668e-07, 
    2.305298e-07, 2.293834e-07, 2.323705e-07, 2.316563e-07, 2.325417e-07, 
    2.3209e-07, 2.328638e-07, 2.321674e-07, 2.333736e-07, 2.336361e-07, 
    2.334568e-07, 2.341458e-07, 2.321288e-07, 2.329037e-07, 2.270652e-07, 
    2.270996e-07, 2.272599e-07, 2.265552e-07, 2.265121e-07, 2.258659e-07, 
    2.264409e-07, 2.266856e-07, 2.273068e-07, 2.276741e-07, 2.280232e-07, 
    2.287905e-07, 2.296468e-07, 2.308435e-07, 2.317026e-07, 2.322782e-07, 
    2.319253e-07, 2.322369e-07, 2.318885e-07, 2.317253e-07, 2.335378e-07, 
    2.325203e-07, 2.340467e-07, 2.339623e-07, 2.332716e-07, 2.339718e-07, 
    2.271238e-07, 2.269258e-07, 2.262381e-07, 2.267763e-07, 2.257955e-07, 
    2.263446e-07, 2.266602e-07, 2.278774e-07, 2.281447e-07, 2.283925e-07, 
    2.288818e-07, 2.295095e-07, 2.3061e-07, 2.315668e-07, 2.324398e-07, 
    2.323758e-07, 2.323983e-07, 2.325933e-07, 2.321103e-07, 2.326725e-07, 
    2.327668e-07, 2.325202e-07, 2.33951e-07, 2.335424e-07, 2.339605e-07, 
    2.336945e-07, 2.269902e-07, 2.273233e-07, 2.271433e-07, 2.274818e-07, 
    2.272433e-07, 2.283034e-07, 2.28621e-07, 2.301066e-07, 2.294971e-07, 
    2.30467e-07, 2.295957e-07, 2.297501e-07, 2.304986e-07, 2.296428e-07, 
    2.315141e-07, 2.302456e-07, 2.326008e-07, 2.313351e-07, 2.326801e-07, 
    2.32436e-07, 2.328402e-07, 2.33202e-07, 2.336572e-07, 2.344966e-07, 
    2.343023e-07, 2.35004e-07, 2.278199e-07, 2.282517e-07, 2.282137e-07, 
    2.286656e-07, 2.289996e-07, 2.297234e-07, 2.308836e-07, 2.304474e-07, 
    2.31248e-07, 2.314087e-07, 2.301923e-07, 2.309393e-07, 2.285407e-07, 
    2.289285e-07, 2.286976e-07, 2.278539e-07, 2.305479e-07, 2.29166e-07, 
    2.317168e-07, 2.309689e-07, 2.331504e-07, 2.320659e-07, 2.341953e-07, 
    2.351045e-07, 2.359598e-07, 2.369585e-07, 2.284874e-07, 2.28194e-07, 
    2.287193e-07, 2.294457e-07, 2.301194e-07, 2.310146e-07, 2.311061e-07, 
    2.312737e-07, 2.317079e-07, 2.320727e-07, 2.313267e-07, 2.321642e-07, 
    2.290183e-07, 2.306678e-07, 2.280831e-07, 2.288618e-07, 2.294029e-07, 
    2.291656e-07, 2.303976e-07, 2.306878e-07, 2.318664e-07, 2.312573e-07, 
    2.348801e-07, 2.332784e-07, 2.377184e-07, 2.364791e-07, 2.280915e-07, 
    2.284864e-07, 2.298599e-07, 2.292065e-07, 2.310743e-07, 2.315337e-07, 
    2.31907e-07, 2.323841e-07, 2.324356e-07, 2.327182e-07, 2.322551e-07, 
    2.326999e-07, 2.310165e-07, 2.31769e-07, 2.29703e-07, 2.302061e-07, 
    2.299747e-07, 2.297208e-07, 2.305043e-07, 2.313385e-07, 2.313563e-07, 
    2.316237e-07, 2.323768e-07, 2.310819e-07, 2.350867e-07, 2.326147e-07, 
    2.289169e-07, 2.296769e-07, 2.297855e-07, 2.294911e-07, 2.314876e-07, 
    2.307645e-07, 2.327113e-07, 2.321854e-07, 2.330469e-07, 2.326189e-07, 
    2.325559e-07, 2.320059e-07, 2.316634e-07, 2.307977e-07, 2.300929e-07, 
    2.295339e-07, 2.296639e-07, 2.30278e-07, 2.313895e-07, 2.324402e-07, 
    2.322101e-07, 2.329815e-07, 2.30939e-07, 2.317958e-07, 2.314647e-07, 
    2.323278e-07, 2.304358e-07, 2.32047e-07, 2.300237e-07, 2.302012e-07, 
    2.307502e-07, 2.318538e-07, 2.320979e-07, 2.323585e-07, 2.321977e-07, 
    2.314177e-07, 2.312899e-07, 2.307369e-07, 2.305841e-07, 2.301626e-07, 
    2.298134e-07, 2.301324e-07, 2.304673e-07, 2.31418e-07, 2.322743e-07, 
    2.332072e-07, 2.334354e-07, 2.345244e-07, 2.336379e-07, 2.351004e-07, 
    2.338571e-07, 2.360087e-07, 2.321404e-07, 2.338206e-07, 2.307752e-07, 
    2.311036e-07, 2.316974e-07, 2.330583e-07, 2.323238e-07, 2.331828e-07, 
    2.312849e-07, 2.302991e-07, 2.30044e-07, 2.295678e-07, 2.300549e-07, 
    2.300153e-07, 2.304812e-07, 2.303315e-07, 2.314496e-07, 2.308491e-07, 
    2.325543e-07, 2.331761e-07, 2.349304e-07, 2.360048e-07, 2.370976e-07, 
    2.375798e-07, 2.377265e-07, 2.377878e-07,
  2.166373e-07, 2.176638e-07, 2.174643e-07, 2.182921e-07, 2.178329e-07, 
    2.18375e-07, 2.168454e-07, 2.177046e-07, 2.171561e-07, 2.167297e-07, 
    2.198984e-07, 2.18329e-07, 2.215279e-07, 2.205274e-07, 2.230404e-07, 
    2.213723e-07, 2.233766e-07, 2.229922e-07, 2.241491e-07, 2.238177e-07, 
    2.252972e-07, 2.24302e-07, 2.260639e-07, 2.250595e-07, 2.252167e-07, 
    2.242692e-07, 2.186449e-07, 2.19703e-07, 2.185822e-07, 2.187331e-07, 
    2.186654e-07, 2.178424e-07, 2.174276e-07, 2.165588e-07, 2.167165e-07, 
    2.173547e-07, 2.188009e-07, 2.1831e-07, 2.195471e-07, 2.195192e-07, 
    2.208962e-07, 2.202754e-07, 2.225892e-07, 2.219317e-07, 2.238315e-07, 
    2.233538e-07, 2.238091e-07, 2.236711e-07, 2.238109e-07, 2.231102e-07, 
    2.234105e-07, 2.227939e-07, 2.203917e-07, 2.210978e-07, 2.189915e-07, 
    2.177247e-07, 2.168831e-07, 2.162858e-07, 2.163703e-07, 2.165312e-07, 
    2.173584e-07, 2.18136e-07, 2.187284e-07, 2.191248e-07, 2.195152e-07, 
    2.206969e-07, 2.213223e-07, 2.227222e-07, 2.224696e-07, 2.228975e-07, 
    2.233063e-07, 2.239925e-07, 2.238796e-07, 2.241819e-07, 2.228862e-07, 
    2.237474e-07, 2.223257e-07, 2.227145e-07, 2.196214e-07, 2.184425e-07, 
    2.179413e-07, 2.175026e-07, 2.164352e-07, 2.171724e-07, 2.168818e-07, 
    2.175731e-07, 2.180123e-07, 2.17795e-07, 2.191356e-07, 2.186145e-07, 
    2.213593e-07, 2.201772e-07, 2.232586e-07, 2.225214e-07, 2.234353e-07, 
    2.22969e-07, 2.23768e-07, 2.230489e-07, 2.242944e-07, 2.245656e-07, 
    2.243803e-07, 2.250921e-07, 2.23009e-07, 2.238091e-07, 2.17789e-07, 
    2.178244e-07, 2.179895e-07, 2.172639e-07, 2.172195e-07, 2.165545e-07, 
    2.171462e-07, 2.173982e-07, 2.180377e-07, 2.18416e-07, 2.187756e-07, 
    2.19566e-07, 2.204488e-07, 2.216828e-07, 2.225692e-07, 2.231633e-07, 
    2.22799e-07, 2.231206e-07, 2.227611e-07, 2.225926e-07, 2.24464e-07, 
    2.234133e-07, 2.249897e-07, 2.249025e-07, 2.241891e-07, 2.249123e-07, 
    2.178493e-07, 2.176454e-07, 2.169375e-07, 2.174915e-07, 2.164821e-07, 
    2.170471e-07, 2.17372e-07, 2.186254e-07, 2.189007e-07, 2.19156e-07, 
    2.196602e-07, 2.203072e-07, 2.214419e-07, 2.224291e-07, 2.233301e-07, 
    2.232641e-07, 2.232873e-07, 2.234886e-07, 2.2299e-07, 2.235704e-07, 
    2.236678e-07, 2.234131e-07, 2.248908e-07, 2.244687e-07, 2.249007e-07, 
    2.246258e-07, 2.177117e-07, 2.180547e-07, 2.178693e-07, 2.182179e-07, 
    2.179724e-07, 2.190642e-07, 2.193915e-07, 2.209228e-07, 2.202944e-07, 
    2.212945e-07, 2.20396e-07, 2.205552e-07, 2.213271e-07, 2.204446e-07, 
    2.223747e-07, 2.210662e-07, 2.234964e-07, 2.2219e-07, 2.235782e-07, 
    2.233262e-07, 2.237435e-07, 2.241172e-07, 2.245873e-07, 2.254547e-07, 
    2.252539e-07, 2.259791e-07, 2.185661e-07, 2.19011e-07, 2.189718e-07, 
    2.194373e-07, 2.197816e-07, 2.205277e-07, 2.217241e-07, 2.212742e-07, 
    2.221001e-07, 2.222659e-07, 2.210112e-07, 2.217816e-07, 2.193087e-07, 
    2.197083e-07, 2.194704e-07, 2.186012e-07, 2.213779e-07, 2.199531e-07, 
    2.225838e-07, 2.218122e-07, 2.240639e-07, 2.229442e-07, 2.251433e-07, 
    2.260831e-07, 2.269674e-07, 2.280007e-07, 2.192537e-07, 2.189515e-07, 
    2.194927e-07, 2.202414e-07, 2.20936e-07, 2.218593e-07, 2.219537e-07, 
    2.221267e-07, 2.225746e-07, 2.229512e-07, 2.221813e-07, 2.230456e-07, 
    2.19801e-07, 2.215016e-07, 2.188372e-07, 2.196397e-07, 2.201973e-07, 
    2.199527e-07, 2.212228e-07, 2.215221e-07, 2.227383e-07, 2.221096e-07, 
    2.258512e-07, 2.241962e-07, 2.287873e-07, 2.275047e-07, 2.188459e-07, 
    2.192527e-07, 2.206684e-07, 2.199949e-07, 2.219209e-07, 2.223949e-07, 
    2.227801e-07, 2.232726e-07, 2.233258e-07, 2.236175e-07, 2.231394e-07, 
    2.235986e-07, 2.218612e-07, 2.226377e-07, 2.205066e-07, 2.210254e-07, 
    2.207867e-07, 2.20525e-07, 2.213329e-07, 2.221935e-07, 2.222118e-07, 
    2.224878e-07, 2.232653e-07, 2.219287e-07, 2.260648e-07, 2.235109e-07, 
    2.196963e-07, 2.204798e-07, 2.205917e-07, 2.202882e-07, 2.223473e-07, 
    2.216013e-07, 2.236104e-07, 2.230675e-07, 2.23957e-07, 2.23515e-07, 
    2.2345e-07, 2.228822e-07, 2.225287e-07, 2.216355e-07, 2.209087e-07, 
    2.203322e-07, 2.204663e-07, 2.210995e-07, 2.222461e-07, 2.233306e-07, 
    2.23093e-07, 2.238894e-07, 2.217812e-07, 2.226653e-07, 2.223237e-07, 
    2.232145e-07, 2.212623e-07, 2.229248e-07, 2.208373e-07, 2.210203e-07, 
    2.215865e-07, 2.227253e-07, 2.229772e-07, 2.232462e-07, 2.230802e-07, 
    2.222752e-07, 2.221433e-07, 2.215728e-07, 2.214152e-07, 2.209805e-07, 
    2.206205e-07, 2.209494e-07, 2.212948e-07, 2.222755e-07, 2.231592e-07, 
    2.241225e-07, 2.243582e-07, 2.254835e-07, 2.245675e-07, 2.26079e-07, 
    2.24794e-07, 2.270182e-07, 2.230211e-07, 2.247562e-07, 2.216123e-07, 
    2.219511e-07, 2.225638e-07, 2.239689e-07, 2.232103e-07, 2.240974e-07, 
    2.221381e-07, 2.211213e-07, 2.208582e-07, 2.203673e-07, 2.208694e-07, 
    2.208286e-07, 2.213091e-07, 2.211547e-07, 2.223081e-07, 2.216886e-07, 
    2.234484e-07, 2.240904e-07, 2.259031e-07, 2.270141e-07, 2.281447e-07, 
    2.286437e-07, 2.287956e-07, 2.288591e-07,
  2.081374e-07, 2.091062e-07, 2.089178e-07, 2.096996e-07, 2.092658e-07, 
    2.097778e-07, 2.083337e-07, 2.091447e-07, 2.086269e-07, 2.082245e-07, 
    2.112181e-07, 2.097344e-07, 2.127605e-07, 2.118132e-07, 2.141942e-07, 
    2.126131e-07, 2.145132e-07, 2.141484e-07, 2.152463e-07, 2.149317e-07, 
    2.16337e-07, 2.153915e-07, 2.170659e-07, 2.161111e-07, 2.162604e-07, 
    2.153603e-07, 2.100328e-07, 2.110333e-07, 2.099736e-07, 2.101162e-07, 
    2.100522e-07, 2.092748e-07, 2.088832e-07, 2.080633e-07, 2.082121e-07, 
    2.088143e-07, 2.101803e-07, 2.097164e-07, 2.108857e-07, 2.108593e-07, 
    2.121622e-07, 2.115746e-07, 2.137663e-07, 2.13143e-07, 2.149448e-07, 
    2.144914e-07, 2.149235e-07, 2.147925e-07, 2.149252e-07, 2.142604e-07, 
    2.145452e-07, 2.139603e-07, 2.116847e-07, 2.123531e-07, 2.103605e-07, 
    2.091637e-07, 2.083693e-07, 2.078058e-07, 2.078854e-07, 2.080373e-07, 
    2.088178e-07, 2.09552e-07, 2.101118e-07, 2.104863e-07, 2.108555e-07, 
    2.119737e-07, 2.125657e-07, 2.138924e-07, 2.136528e-07, 2.140586e-07, 
    2.144463e-07, 2.150976e-07, 2.149904e-07, 2.152774e-07, 2.140479e-07, 
    2.148649e-07, 2.135164e-07, 2.138851e-07, 2.109561e-07, 2.098416e-07, 
    2.093683e-07, 2.08954e-07, 2.079467e-07, 2.086422e-07, 2.08368e-07, 
    2.090205e-07, 2.094352e-07, 2.092301e-07, 2.104966e-07, 2.100041e-07, 
    2.126008e-07, 2.114817e-07, 2.144011e-07, 2.13702e-07, 2.145687e-07, 
    2.141264e-07, 2.148845e-07, 2.142022e-07, 2.153843e-07, 2.156418e-07, 
    2.154658e-07, 2.16142e-07, 2.141643e-07, 2.149235e-07, 2.092243e-07, 
    2.092578e-07, 2.094136e-07, 2.087286e-07, 2.086867e-07, 2.080592e-07, 
    2.086175e-07, 2.088554e-07, 2.094592e-07, 2.098166e-07, 2.101563e-07, 
    2.109036e-07, 2.117387e-07, 2.129072e-07, 2.137473e-07, 2.143107e-07, 
    2.139652e-07, 2.142702e-07, 2.139292e-07, 2.137694e-07, 2.155453e-07, 
    2.145479e-07, 2.160447e-07, 2.159618e-07, 2.152843e-07, 2.159712e-07, 
    2.092813e-07, 2.090887e-07, 2.084206e-07, 2.089434e-07, 2.079909e-07, 
    2.08524e-07, 2.088307e-07, 2.100144e-07, 2.102746e-07, 2.105159e-07, 
    2.109926e-07, 2.116047e-07, 2.12679e-07, 2.136145e-07, 2.144689e-07, 
    2.144063e-07, 2.144283e-07, 2.146193e-07, 2.141463e-07, 2.14697e-07, 
    2.147894e-07, 2.145477e-07, 2.159507e-07, 2.155498e-07, 2.159601e-07, 
    2.15699e-07, 2.091513e-07, 2.094753e-07, 2.093002e-07, 2.096294e-07, 
    2.093975e-07, 2.104292e-07, 2.107386e-07, 2.121875e-07, 2.115926e-07, 
    2.125394e-07, 2.116888e-07, 2.118395e-07, 2.125704e-07, 2.117347e-07, 
    2.135629e-07, 2.123233e-07, 2.146267e-07, 2.133879e-07, 2.147044e-07, 
    2.144652e-07, 2.148612e-07, 2.15216e-07, 2.156624e-07, 2.164866e-07, 
    2.162957e-07, 2.169853e-07, 2.099584e-07, 2.103788e-07, 2.103418e-07, 
    2.107819e-07, 2.111075e-07, 2.118134e-07, 2.129463e-07, 2.125202e-07, 
    2.133026e-07, 2.134597e-07, 2.12271e-07, 2.130008e-07, 2.106603e-07, 
    2.110382e-07, 2.108131e-07, 2.099916e-07, 2.126184e-07, 2.112697e-07, 
    2.137612e-07, 2.130298e-07, 2.151654e-07, 2.141029e-07, 2.161907e-07, 
    2.170842e-07, 2.179256e-07, 2.189098e-07, 2.106083e-07, 2.103226e-07, 
    2.108342e-07, 2.115425e-07, 2.121999e-07, 2.130744e-07, 2.131638e-07, 
    2.133278e-07, 2.137524e-07, 2.141095e-07, 2.133796e-07, 2.14199e-07, 
    2.11126e-07, 2.127355e-07, 2.102146e-07, 2.109733e-07, 2.115007e-07, 
    2.112693e-07, 2.124715e-07, 2.12755e-07, 2.139076e-07, 2.133116e-07, 
    2.168637e-07, 2.15291e-07, 2.196595e-07, 2.184372e-07, 2.102227e-07, 
    2.106073e-07, 2.119466e-07, 2.113092e-07, 2.131328e-07, 2.13582e-07, 
    2.139473e-07, 2.144144e-07, 2.144648e-07, 2.147417e-07, 2.14288e-07, 
    2.147237e-07, 2.130762e-07, 2.138122e-07, 2.117934e-07, 2.122845e-07, 
    2.120586e-07, 2.118108e-07, 2.125757e-07, 2.133911e-07, 2.134085e-07, 
    2.136701e-07, 2.144076e-07, 2.131401e-07, 2.17067e-07, 2.146406e-07, 
    2.110268e-07, 2.117681e-07, 2.11874e-07, 2.115867e-07, 2.135369e-07, 
    2.1283e-07, 2.147349e-07, 2.142198e-07, 2.150639e-07, 2.146444e-07, 
    2.145827e-07, 2.140441e-07, 2.137089e-07, 2.128624e-07, 2.12174e-07, 
    2.116284e-07, 2.117552e-07, 2.123547e-07, 2.13441e-07, 2.144694e-07, 
    2.142441e-07, 2.149997e-07, 2.130004e-07, 2.138385e-07, 2.135145e-07, 
    2.143593e-07, 2.125089e-07, 2.140847e-07, 2.121064e-07, 2.122797e-07, 
    2.12816e-07, 2.138954e-07, 2.141342e-07, 2.143893e-07, 2.142319e-07, 
    2.134686e-07, 2.133436e-07, 2.128029e-07, 2.126537e-07, 2.12242e-07, 
    2.119012e-07, 2.122126e-07, 2.125396e-07, 2.134689e-07, 2.143069e-07, 
    2.152211e-07, 2.154448e-07, 2.165141e-07, 2.156437e-07, 2.170805e-07, 
    2.15859e-07, 2.179741e-07, 2.14176e-07, 2.15823e-07, 2.128404e-07, 
    2.131614e-07, 2.137422e-07, 2.150752e-07, 2.143553e-07, 2.151972e-07, 
    2.133386e-07, 2.123754e-07, 2.121262e-07, 2.116616e-07, 2.121369e-07, 
    2.120982e-07, 2.125531e-07, 2.124069e-07, 2.134997e-07, 2.129126e-07, 
    2.145812e-07, 2.151906e-07, 2.16913e-07, 2.179701e-07, 2.190468e-07, 
    2.195225e-07, 2.196673e-07, 2.197279e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.35703e-08, 6.384985e-08, 6.379551e-08, 6.402099e-08, 6.389591e-08, 
    6.404356e-08, 6.362697e-08, 6.386096e-08, 6.371158e-08, 6.359546e-08, 
    6.445858e-08, 6.403105e-08, 6.490264e-08, 6.462999e-08, 6.531489e-08, 
    6.486022e-08, 6.540657e-08, 6.530176e-08, 6.561717e-08, 6.552681e-08, 
    6.593026e-08, 6.565888e-08, 6.613939e-08, 6.586544e-08, 6.59083e-08, 
    6.564993e-08, 6.411708e-08, 6.440536e-08, 6.410001e-08, 6.414111e-08, 
    6.412267e-08, 6.38985e-08, 6.378554e-08, 6.354892e-08, 6.359188e-08, 
    6.376565e-08, 6.41596e-08, 6.402587e-08, 6.436288e-08, 6.435527e-08, 
    6.473046e-08, 6.45613e-08, 6.519191e-08, 6.501268e-08, 6.553059e-08, 
    6.540034e-08, 6.552447e-08, 6.548683e-08, 6.552496e-08, 6.533394e-08, 
    6.541578e-08, 6.524769e-08, 6.459298e-08, 6.47854e-08, 6.421152e-08, 
    6.386645e-08, 6.363724e-08, 6.347459e-08, 6.349758e-08, 6.354141e-08, 
    6.376668e-08, 6.397845e-08, 6.413985e-08, 6.424781e-08, 6.435418e-08, 
    6.467617e-08, 6.484658e-08, 6.522815e-08, 6.515928e-08, 6.527594e-08, 
    6.538738e-08, 6.557449e-08, 6.554369e-08, 6.562612e-08, 6.527286e-08, 
    6.550764e-08, 6.512006e-08, 6.522607e-08, 6.438312e-08, 6.406194e-08, 
    6.392545e-08, 6.380596e-08, 6.351526e-08, 6.371601e-08, 6.363688e-08, 
    6.382514e-08, 6.394477e-08, 6.38856e-08, 6.425076e-08, 6.41088e-08, 
    6.485669e-08, 6.453455e-08, 6.537438e-08, 6.517342e-08, 6.542255e-08, 
    6.529542e-08, 6.551326e-08, 6.531721e-08, 6.565681e-08, 6.573075e-08, 
    6.568022e-08, 6.587433e-08, 6.530634e-08, 6.552447e-08, 6.388395e-08, 
    6.389359e-08, 6.393855e-08, 6.374094e-08, 6.372885e-08, 6.354775e-08, 
    6.370889e-08, 6.377751e-08, 6.39517e-08, 6.405474e-08, 6.415268e-08, 
    6.436803e-08, 6.460854e-08, 6.494484e-08, 6.518644e-08, 6.53484e-08, 
    6.524908e-08, 6.533676e-08, 6.523875e-08, 6.519281e-08, 6.570305e-08, 
    6.541654e-08, 6.584641e-08, 6.582263e-08, 6.562809e-08, 6.58253e-08, 
    6.390037e-08, 6.384484e-08, 6.365205e-08, 6.380292e-08, 6.352803e-08, 
    6.36819e-08, 6.377039e-08, 6.411177e-08, 6.418676e-08, 6.425632e-08, 
    6.439367e-08, 6.456996e-08, 6.48792e-08, 6.514825e-08, 6.539386e-08, 
    6.537586e-08, 6.53822e-08, 6.543707e-08, 6.530116e-08, 6.545939e-08, 
    6.548594e-08, 6.541651e-08, 6.581944e-08, 6.570433e-08, 6.582212e-08, 
    6.574717e-08, 6.386289e-08, 6.395633e-08, 6.390584e-08, 6.400078e-08, 
    6.39339e-08, 6.423132e-08, 6.432049e-08, 6.473773e-08, 6.456649e-08, 
    6.483902e-08, 6.459417e-08, 6.463756e-08, 6.484792e-08, 6.46074e-08, 
    6.513343e-08, 6.477681e-08, 6.543921e-08, 6.508311e-08, 6.546152e-08, 
    6.53928e-08, 6.550658e-08, 6.560848e-08, 6.573668e-08, 6.597322e-08, 
    6.591844e-08, 6.611626e-08, 6.409562e-08, 6.421681e-08, 6.420614e-08, 
    6.433297e-08, 6.442676e-08, 6.463005e-08, 6.49561e-08, 6.483349e-08, 
    6.505858e-08, 6.510377e-08, 6.47618e-08, 6.497177e-08, 6.429792e-08, 
    6.44068e-08, 6.434197e-08, 6.410518e-08, 6.486175e-08, 6.447348e-08, 
    6.519043e-08, 6.498011e-08, 6.559395e-08, 6.528868e-08, 6.588829e-08, 
    6.614464e-08, 6.638587e-08, 6.66678e-08, 6.428295e-08, 6.42006e-08, 
    6.434804e-08, 6.455205e-08, 6.474131e-08, 6.499293e-08, 6.501867e-08, 
    6.506582e-08, 6.518791e-08, 6.529058e-08, 6.508073e-08, 6.531631e-08, 
    6.443206e-08, 6.489545e-08, 6.416948e-08, 6.438809e-08, 6.454002e-08, 
    6.447337e-08, 6.481947e-08, 6.490105e-08, 6.523254e-08, 6.506118e-08, 
    6.608137e-08, 6.563001e-08, 6.688245e-08, 6.653246e-08, 6.417183e-08, 
    6.428267e-08, 6.466841e-08, 6.448487e-08, 6.500973e-08, 6.513893e-08, 
    6.524394e-08, 6.53782e-08, 6.539269e-08, 6.547224e-08, 6.534189e-08, 
    6.546708e-08, 6.499347e-08, 6.520511e-08, 6.462431e-08, 6.476568e-08, 
    6.470064e-08, 6.46293e-08, 6.484947e-08, 6.508403e-08, 6.508903e-08, 
    6.516425e-08, 6.537621e-08, 6.501185e-08, 6.613964e-08, 6.544317e-08, 
    6.440352e-08, 6.461701e-08, 6.464749e-08, 6.456479e-08, 6.512597e-08, 
    6.492264e-08, 6.54703e-08, 6.532228e-08, 6.55648e-08, 6.544429e-08, 
    6.542655e-08, 6.527178e-08, 6.517542e-08, 6.493197e-08, 6.473388e-08, 
    6.457679e-08, 6.461332e-08, 6.478587e-08, 6.509838e-08, 6.5394e-08, 
    6.532925e-08, 6.554637e-08, 6.497167e-08, 6.521266e-08, 6.511952e-08, 
    6.536237e-08, 6.483023e-08, 6.528341e-08, 6.471441e-08, 6.476429e-08, 
    6.49186e-08, 6.522901e-08, 6.529767e-08, 6.5371e-08, 6.532575e-08, 
    6.510631e-08, 6.507035e-08, 6.491485e-08, 6.487192e-08, 6.475343e-08, 
    6.465533e-08, 6.474496e-08, 6.483909e-08, 6.51064e-08, 6.534729e-08, 
    6.560993e-08, 6.56742e-08, 6.598109e-08, 6.573129e-08, 6.614352e-08, 
    6.579306e-08, 6.639972e-08, 6.530966e-08, 6.578274e-08, 6.492562e-08, 
    6.501796e-08, 6.518498e-08, 6.556804e-08, 6.536123e-08, 6.560308e-08, 
    6.506895e-08, 6.479183e-08, 6.472012e-08, 6.458635e-08, 6.472317e-08, 
    6.471205e-08, 6.484298e-08, 6.480091e-08, 6.511527e-08, 6.494641e-08, 
    6.542611e-08, 6.560117e-08, 6.609553e-08, 6.639859e-08, 6.670707e-08, 
    6.684326e-08, 6.688472e-08, 6.690204e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  8.582233e-13, 8.605457e-13, 8.600946e-13, 8.61966e-13, 8.609284e-13, 
    8.621533e-13, 8.586947e-13, 8.606376e-13, 8.593977e-13, 8.58433e-13, 
    8.655925e-13, 8.620496e-13, 8.692698e-13, 8.670143e-13, 8.726766e-13, 
    8.689185e-13, 8.734338e-13, 8.725691e-13, 8.751727e-13, 8.744272e-13, 
    8.777522e-13, 8.755167e-13, 8.794752e-13, 8.77219e-13, 8.775718e-13, 
    8.754428e-13, 8.627638e-13, 8.651514e-13, 8.62622e-13, 8.629628e-13, 
    8.628101e-13, 8.609495e-13, 8.600109e-13, 8.580462e-13, 8.584032e-13, 
    8.598464e-13, 8.631159e-13, 8.620071e-13, 8.648021e-13, 8.647391e-13, 
    8.678461e-13, 8.664457e-13, 8.716615e-13, 8.701809e-13, 8.744583e-13, 
    8.733831e-13, 8.744077e-13, 8.740972e-13, 8.744117e-13, 8.728347e-13, 
    8.735105e-13, 8.721225e-13, 8.667079e-13, 8.683005e-13, 8.635468e-13, 
    8.606823e-13, 8.587798e-13, 8.574282e-13, 8.576193e-13, 8.579834e-13, 
    8.598548e-13, 8.616137e-13, 8.629528e-13, 8.638481e-13, 8.6473e-13, 
    8.673951e-13, 8.688061e-13, 8.719605e-13, 8.713922e-13, 8.723554e-13, 
    8.732762e-13, 8.748203e-13, 8.745663e-13, 8.752462e-13, 8.723305e-13, 
    8.742684e-13, 8.710687e-13, 8.719439e-13, 8.64967e-13, 8.623064e-13, 
    8.611724e-13, 8.601812e-13, 8.577662e-13, 8.594341e-13, 8.587766e-13, 
    8.60341e-13, 8.613341e-13, 8.60843e-13, 8.638726e-13, 8.626952e-13, 
    8.688898e-13, 8.662237e-13, 8.731688e-13, 8.715089e-13, 8.735666e-13, 
    8.72517e-13, 8.743149e-13, 8.726968e-13, 8.754994e-13, 8.761088e-13, 
    8.756923e-13, 8.772928e-13, 8.726071e-13, 8.744074e-13, 8.608291e-13, 
    8.609092e-13, 8.612826e-13, 8.596411e-13, 8.595408e-13, 8.580363e-13, 
    8.593753e-13, 8.59945e-13, 8.613918e-13, 8.622466e-13, 8.630591e-13, 
    8.648445e-13, 8.668363e-13, 8.696193e-13, 8.716165e-13, 8.729544e-13, 
    8.721343e-13, 8.728583e-13, 8.720488e-13, 8.716694e-13, 8.758803e-13, 
    8.735166e-13, 8.770627e-13, 8.768667e-13, 8.752623e-13, 8.768888e-13, 
    8.609655e-13, 8.605046e-13, 8.58903e-13, 8.601565e-13, 8.578724e-13, 
    8.591509e-13, 8.598855e-13, 8.627192e-13, 8.63342e-13, 8.639184e-13, 
    8.650572e-13, 8.665174e-13, 8.690765e-13, 8.713006e-13, 8.733298e-13, 
    8.731813e-13, 8.732336e-13, 8.736864e-13, 8.725642e-13, 8.738706e-13, 
    8.740895e-13, 8.735166e-13, 8.768404e-13, 8.758914e-13, 8.768625e-13, 
    8.762447e-13, 8.606545e-13, 8.6143e-13, 8.61011e-13, 8.617988e-13, 
    8.612435e-13, 8.637105e-13, 8.644496e-13, 8.679055e-13, 8.664885e-13, 
    8.68744e-13, 8.667179e-13, 8.670769e-13, 8.688164e-13, 8.668277e-13, 
    8.71178e-13, 8.682285e-13, 8.73704e-13, 8.707614e-13, 8.738882e-13, 
    8.733211e-13, 8.742602e-13, 8.751007e-13, 8.761581e-13, 8.78107e-13, 
    8.77656e-13, 8.792853e-13, 8.625859e-13, 8.635906e-13, 8.635026e-13, 
    8.64554e-13, 8.653311e-13, 8.670152e-13, 8.697128e-13, 8.686989e-13, 
    8.705605e-13, 8.709338e-13, 8.681058e-13, 8.698421e-13, 8.642631e-13, 
    8.651649e-13, 8.646285e-13, 8.626649e-13, 8.689319e-13, 8.657175e-13, 
    8.716494e-13, 8.699114e-13, 8.749808e-13, 8.724604e-13, 8.774076e-13, 
    8.795176e-13, 8.81504e-13, 8.8382e-13, 8.641393e-13, 8.634568e-13, 
    8.646792e-13, 8.663683e-13, 8.679359e-13, 8.700174e-13, 8.702305e-13, 
    8.706201e-13, 8.716289e-13, 8.724769e-13, 8.707427e-13, 8.726895e-13, 
    8.65373e-13, 8.692109e-13, 8.631982e-13, 8.650098e-13, 8.66269e-13, 
    8.657173e-13, 8.685831e-13, 8.692578e-13, 8.719969e-13, 8.705819e-13, 
    8.789965e-13, 8.752774e-13, 8.855835e-13, 8.827082e-13, 8.632181e-13, 
    8.641372e-13, 8.673321e-13, 8.658126e-13, 8.701565e-13, 8.712243e-13, 
    8.720918e-13, 8.732001e-13, 8.733201e-13, 8.739765e-13, 8.729007e-13, 
    8.739342e-13, 8.700218e-13, 8.717709e-13, 8.669677e-13, 8.681375e-13, 
    8.675997e-13, 8.670091e-13, 8.688312e-13, 8.707699e-13, 8.708122e-13, 
    8.714328e-13, 8.731807e-13, 8.701742e-13, 8.794746e-13, 8.737338e-13, 
    8.651389e-13, 8.669062e-13, 8.671594e-13, 8.664749e-13, 8.711172e-13, 
    8.694361e-13, 8.739606e-13, 8.727388e-13, 8.747405e-13, 8.73746e-13, 
    8.735996e-13, 8.723216e-13, 8.715254e-13, 8.695131e-13, 8.678743e-13, 
    8.665743e-13, 8.668767e-13, 8.683045e-13, 8.708886e-13, 8.733305e-13, 
    8.727957e-13, 8.745885e-13, 8.698418e-13, 8.718328e-13, 8.710635e-13, 
    8.730696e-13, 8.686718e-13, 8.724148e-13, 8.677136e-13, 8.681264e-13, 
    8.694028e-13, 8.719672e-13, 8.725355e-13, 8.731406e-13, 8.727674e-13, 
    8.709544e-13, 8.706574e-13, 8.69372e-13, 8.690165e-13, 8.680366e-13, 
    8.672246e-13, 8.679663e-13, 8.687447e-13, 8.709555e-13, 8.729448e-13, 
    8.751125e-13, 8.75643e-13, 8.781703e-13, 8.761121e-13, 8.795063e-13, 
    8.766191e-13, 8.816153e-13, 8.726327e-13, 8.765359e-13, 8.694611e-13, 
    8.702247e-13, 8.716036e-13, 8.747661e-13, 8.730603e-13, 8.750555e-13, 
    8.706459e-13, 8.683533e-13, 8.677608e-13, 8.666532e-13, 8.677861e-13, 
    8.67694e-13, 8.687776e-13, 8.684295e-13, 8.710288e-13, 8.69633e-13, 
    8.735957e-13, 8.750399e-13, 8.791143e-13, 8.816076e-13, 8.841439e-13, 
    8.852622e-13, 8.856025e-13, 8.857447e-13 ;

 LITR1C =
  3.066807e-05, 3.066795e-05, 3.066797e-05, 3.066788e-05, 3.066793e-05, 
    3.066787e-05, 3.066804e-05, 3.066794e-05, 3.066801e-05, 3.066806e-05, 
    3.06677e-05, 3.066787e-05, 3.066751e-05, 3.066762e-05, 3.066734e-05, 
    3.066753e-05, 3.06673e-05, 3.066735e-05, 3.066722e-05, 3.066725e-05, 
    3.066708e-05, 3.06672e-05, 3.0667e-05, 3.066711e-05, 3.06671e-05, 
    3.06672e-05, 3.066784e-05, 3.066772e-05, 3.066784e-05, 3.066783e-05, 
    3.066783e-05, 3.066793e-05, 3.066798e-05, 3.066807e-05, 3.066806e-05, 
    3.066798e-05, 3.066782e-05, 3.066788e-05, 3.066774e-05, 3.066774e-05, 
    3.066758e-05, 3.066765e-05, 3.066739e-05, 3.066747e-05, 3.066725e-05, 
    3.06673e-05, 3.066725e-05, 3.066727e-05, 3.066725e-05, 3.066733e-05, 
    3.06673e-05, 3.066737e-05, 3.066764e-05, 3.066756e-05, 3.06678e-05, 
    3.066794e-05, 3.066804e-05, 3.066811e-05, 3.06681e-05, 3.066808e-05, 
    3.066798e-05, 3.06679e-05, 3.066783e-05, 3.066778e-05, 3.066774e-05, 
    3.06676e-05, 3.066754e-05, 3.066738e-05, 3.06674e-05, 3.066736e-05, 
    3.066731e-05, 3.066723e-05, 3.066724e-05, 3.066721e-05, 3.066736e-05, 
    3.066726e-05, 3.066742e-05, 3.066738e-05, 3.066773e-05, 3.066786e-05, 
    3.066792e-05, 3.066797e-05, 3.066809e-05, 3.0668e-05, 3.066804e-05, 
    3.066796e-05, 3.066791e-05, 3.066794e-05, 3.066778e-05, 3.066784e-05, 
    3.066753e-05, 3.066766e-05, 3.066731e-05, 3.06674e-05, 3.06673e-05, 
    3.066735e-05, 3.066726e-05, 3.066734e-05, 3.06672e-05, 3.066717e-05, 
    3.066719e-05, 3.066711e-05, 3.066734e-05, 3.066725e-05, 3.066794e-05, 
    3.066793e-05, 3.066791e-05, 3.066799e-05, 3.0668e-05, 3.066807e-05, 
    3.066801e-05, 3.066798e-05, 3.066791e-05, 3.066786e-05, 3.066782e-05, 
    3.066773e-05, 3.066763e-05, 3.066749e-05, 3.066739e-05, 3.066732e-05, 
    3.066737e-05, 3.066733e-05, 3.066737e-05, 3.066739e-05, 3.066718e-05, 
    3.06673e-05, 3.066712e-05, 3.066713e-05, 3.066721e-05, 3.066713e-05, 
    3.066793e-05, 3.066795e-05, 3.066803e-05, 3.066797e-05, 3.066808e-05, 
    3.066802e-05, 3.066798e-05, 3.066784e-05, 3.066781e-05, 3.066778e-05, 
    3.066772e-05, 3.066765e-05, 3.066752e-05, 3.066741e-05, 3.066731e-05, 
    3.066731e-05, 3.066731e-05, 3.066729e-05, 3.066735e-05, 3.066728e-05, 
    3.066727e-05, 3.06673e-05, 3.066713e-05, 3.066718e-05, 3.066713e-05, 
    3.066716e-05, 3.066794e-05, 3.066791e-05, 3.066792e-05, 3.066788e-05, 
    3.066791e-05, 3.066779e-05, 3.066775e-05, 3.066758e-05, 3.066765e-05, 
    3.066754e-05, 3.066764e-05, 3.066762e-05, 3.066753e-05, 3.066763e-05, 
    3.066742e-05, 3.066756e-05, 3.066729e-05, 3.066744e-05, 3.066728e-05, 
    3.066731e-05, 3.066726e-05, 3.066722e-05, 3.066716e-05, 3.066707e-05, 
    3.066709e-05, 3.066701e-05, 3.066785e-05, 3.06678e-05, 3.06678e-05, 
    3.066775e-05, 3.066771e-05, 3.066762e-05, 3.066749e-05, 3.066754e-05, 
    3.066744e-05, 3.066743e-05, 3.066757e-05, 3.066748e-05, 3.066776e-05, 
    3.066772e-05, 3.066774e-05, 3.066784e-05, 3.066753e-05, 3.066769e-05, 
    3.066739e-05, 3.066748e-05, 3.066722e-05, 3.066735e-05, 3.06671e-05, 
    3.0667e-05, 3.06669e-05, 3.066678e-05, 3.066777e-05, 3.06678e-05, 
    3.066774e-05, 3.066766e-05, 3.066758e-05, 3.066747e-05, 3.066746e-05, 
    3.066744e-05, 3.066739e-05, 3.066735e-05, 3.066744e-05, 3.066734e-05, 
    3.066771e-05, 3.066751e-05, 3.066782e-05, 3.066772e-05, 3.066766e-05, 
    3.066769e-05, 3.066755e-05, 3.066751e-05, 3.066738e-05, 3.066744e-05, 
    3.066702e-05, 3.066721e-05, 3.066669e-05, 3.066684e-05, 3.066782e-05, 
    3.066777e-05, 3.066761e-05, 3.066768e-05, 3.066747e-05, 3.066741e-05, 
    3.066737e-05, 3.066731e-05, 3.066731e-05, 3.066727e-05, 3.066733e-05, 
    3.066728e-05, 3.066747e-05, 3.066739e-05, 3.066763e-05, 3.066757e-05, 
    3.066759e-05, 3.066762e-05, 3.066753e-05, 3.066744e-05, 3.066743e-05, 
    3.06674e-05, 3.066731e-05, 3.066747e-05, 3.0667e-05, 3.066729e-05, 
    3.066772e-05, 3.066763e-05, 3.066762e-05, 3.066765e-05, 3.066742e-05, 
    3.06675e-05, 3.066727e-05, 3.066734e-05, 3.066724e-05, 3.066728e-05, 
    3.066729e-05, 3.066736e-05, 3.06674e-05, 3.06675e-05, 3.066758e-05, 
    3.066764e-05, 3.066763e-05, 3.066756e-05, 3.066743e-05, 3.066731e-05, 
    3.066734e-05, 3.066724e-05, 3.066748e-05, 3.066738e-05, 3.066742e-05, 
    3.066732e-05, 3.066754e-05, 3.066735e-05, 3.066759e-05, 3.066757e-05, 
    3.06675e-05, 3.066738e-05, 3.066735e-05, 3.066732e-05, 3.066734e-05, 
    3.066743e-05, 3.066744e-05, 3.066751e-05, 3.066752e-05, 3.066757e-05, 
    3.066761e-05, 3.066758e-05, 3.066754e-05, 3.066743e-05, 3.066732e-05, 
    3.066722e-05, 3.066719e-05, 3.066706e-05, 3.066717e-05, 3.0667e-05, 
    3.066714e-05, 3.066689e-05, 3.066734e-05, 3.066715e-05, 3.06675e-05, 
    3.066746e-05, 3.066739e-05, 3.066723e-05, 3.066732e-05, 3.066722e-05, 
    3.066744e-05, 3.066756e-05, 3.066759e-05, 3.066764e-05, 3.066759e-05, 
    3.066759e-05, 3.066754e-05, 3.066755e-05, 3.066742e-05, 3.066749e-05, 
    3.06673e-05, 3.066722e-05, 3.066702e-05, 3.066689e-05, 3.066676e-05, 
    3.066671e-05, 3.066669e-05, 3.066668e-05 ;

 LITR1C_TO_SOIL1C =
  5.716177e-13, 5.731643e-13, 5.728639e-13, 5.741101e-13, 5.734191e-13, 
    5.742348e-13, 5.719316e-13, 5.732254e-13, 5.723998e-13, 5.717573e-13, 
    5.76525e-13, 5.741657e-13, 5.789739e-13, 5.774718e-13, 5.812425e-13, 
    5.787399e-13, 5.817468e-13, 5.811709e-13, 5.829048e-13, 5.824083e-13, 
    5.846225e-13, 5.831339e-13, 5.857699e-13, 5.842674e-13, 5.845024e-13, 
    5.830846e-13, 5.746414e-13, 5.762313e-13, 5.74547e-13, 5.747738e-13, 
    5.746721e-13, 5.734332e-13, 5.728081e-13, 5.714998e-13, 5.717375e-13, 
    5.726986e-13, 5.748759e-13, 5.741375e-13, 5.759987e-13, 5.759567e-13, 
    5.780258e-13, 5.770932e-13, 5.805666e-13, 5.795805e-13, 5.82429e-13, 
    5.81713e-13, 5.823953e-13, 5.821885e-13, 5.82398e-13, 5.813478e-13, 
    5.817978e-13, 5.808736e-13, 5.772678e-13, 5.783284e-13, 5.751627e-13, 
    5.732553e-13, 5.719883e-13, 5.710882e-13, 5.712155e-13, 5.71458e-13, 
    5.727042e-13, 5.738754e-13, 5.747672e-13, 5.753634e-13, 5.759507e-13, 
    5.777255e-13, 5.786651e-13, 5.807657e-13, 5.803872e-13, 5.810286e-13, 
    5.816418e-13, 5.826701e-13, 5.82501e-13, 5.829537e-13, 5.81012e-13, 
    5.823026e-13, 5.801718e-13, 5.807546e-13, 5.761085e-13, 5.743368e-13, 
    5.735815e-13, 5.729215e-13, 5.713133e-13, 5.72424e-13, 5.719862e-13, 
    5.73028e-13, 5.736892e-13, 5.733623e-13, 5.753797e-13, 5.745957e-13, 
    5.787208e-13, 5.769454e-13, 5.815703e-13, 5.804649e-13, 5.818352e-13, 
    5.811362e-13, 5.823335e-13, 5.81256e-13, 5.831223e-13, 5.835281e-13, 
    5.832508e-13, 5.843166e-13, 5.811962e-13, 5.823951e-13, 5.73353e-13, 
    5.734063e-13, 5.736549e-13, 5.725619e-13, 5.724951e-13, 5.714932e-13, 
    5.723849e-13, 5.727643e-13, 5.737277e-13, 5.74297e-13, 5.74838e-13, 
    5.76027e-13, 5.773534e-13, 5.792066e-13, 5.805366e-13, 5.814275e-13, 
    5.808814e-13, 5.813636e-13, 5.808245e-13, 5.805718e-13, 5.83376e-13, 
    5.818019e-13, 5.841633e-13, 5.840328e-13, 5.829644e-13, 5.840475e-13, 
    5.734438e-13, 5.731369e-13, 5.720703e-13, 5.729051e-13, 5.71384e-13, 
    5.722354e-13, 5.727246e-13, 5.746116e-13, 5.750264e-13, 5.754103e-13, 
    5.761686e-13, 5.77141e-13, 5.788451e-13, 5.803263e-13, 5.816776e-13, 
    5.815786e-13, 5.816134e-13, 5.819149e-13, 5.811677e-13, 5.820376e-13, 
    5.821834e-13, 5.818019e-13, 5.840153e-13, 5.833833e-13, 5.840301e-13, 
    5.836187e-13, 5.732367e-13, 5.737531e-13, 5.734741e-13, 5.739987e-13, 
    5.73629e-13, 5.752718e-13, 5.757639e-13, 5.780653e-13, 5.771217e-13, 
    5.786237e-13, 5.772745e-13, 5.775136e-13, 5.786719e-13, 5.773476e-13, 
    5.802446e-13, 5.782804e-13, 5.819267e-13, 5.799672e-13, 5.820494e-13, 
    5.816717e-13, 5.822971e-13, 5.828568e-13, 5.83561e-13, 5.848588e-13, 
    5.845584e-13, 5.856434e-13, 5.745229e-13, 5.751919e-13, 5.751334e-13, 
    5.758335e-13, 5.76351e-13, 5.774724e-13, 5.792689e-13, 5.785937e-13, 
    5.798333e-13, 5.800819e-13, 5.781987e-13, 5.79355e-13, 5.756398e-13, 
    5.762403e-13, 5.75883e-13, 5.745754e-13, 5.787489e-13, 5.766083e-13, 
    5.805585e-13, 5.794011e-13, 5.82777e-13, 5.810985e-13, 5.84393e-13, 
    5.857981e-13, 5.871208e-13, 5.886632e-13, 5.755573e-13, 5.751028e-13, 
    5.759168e-13, 5.770417e-13, 5.780856e-13, 5.794717e-13, 5.796136e-13, 
    5.79873e-13, 5.805448e-13, 5.811095e-13, 5.799547e-13, 5.812511e-13, 
    5.763789e-13, 5.789346e-13, 5.749306e-13, 5.76137e-13, 5.769756e-13, 
    5.766082e-13, 5.785166e-13, 5.789659e-13, 5.807899e-13, 5.798476e-13, 
    5.854511e-13, 5.829745e-13, 5.898375e-13, 5.879228e-13, 5.749439e-13, 
    5.755559e-13, 5.776835e-13, 5.766716e-13, 5.795644e-13, 5.802754e-13, 
    5.808531e-13, 5.815911e-13, 5.816711e-13, 5.821081e-13, 5.813918e-13, 
    5.8208e-13, 5.794746e-13, 5.806394e-13, 5.774409e-13, 5.782199e-13, 
    5.778617e-13, 5.774684e-13, 5.786818e-13, 5.799728e-13, 5.800009e-13, 
    5.804142e-13, 5.815782e-13, 5.795761e-13, 5.857694e-13, 5.819465e-13, 
    5.76223e-13, 5.773998e-13, 5.775685e-13, 5.771127e-13, 5.802041e-13, 
    5.790846e-13, 5.820976e-13, 5.812839e-13, 5.82617e-13, 5.819547e-13, 
    5.818572e-13, 5.810062e-13, 5.804759e-13, 5.791359e-13, 5.780446e-13, 
    5.771789e-13, 5.773803e-13, 5.783311e-13, 5.800519e-13, 5.81678e-13, 
    5.813218e-13, 5.825157e-13, 5.793548e-13, 5.806806e-13, 5.801683e-13, 
    5.815043e-13, 5.785756e-13, 5.810682e-13, 5.779375e-13, 5.782124e-13, 
    5.790624e-13, 5.807701e-13, 5.811486e-13, 5.815515e-13, 5.81303e-13, 
    5.800957e-13, 5.798979e-13, 5.790419e-13, 5.788052e-13, 5.781527e-13, 
    5.776119e-13, 5.781058e-13, 5.786242e-13, 5.800964e-13, 5.814211e-13, 
    5.828647e-13, 5.832179e-13, 5.849009e-13, 5.835303e-13, 5.857906e-13, 
    5.83868e-13, 5.871951e-13, 5.812133e-13, 5.838126e-13, 5.791013e-13, 
    5.796097e-13, 5.80528e-13, 5.826339e-13, 5.81498e-13, 5.828266e-13, 
    5.798902e-13, 5.783636e-13, 5.77969e-13, 5.772314e-13, 5.779858e-13, 
    5.779245e-13, 5.786461e-13, 5.784143e-13, 5.801453e-13, 5.792157e-13, 
    5.818546e-13, 5.828163e-13, 5.855295e-13, 5.871899e-13, 5.888789e-13, 
    5.896236e-13, 5.898502e-13, 5.899449e-13 ;

 LITR1C_vr =
  0.001751178, 0.001751172, 0.001751173, 0.001751167, 0.00175117, 
    0.001751167, 0.001751177, 0.001751171, 0.001751175, 0.001751178, 
    0.001751157, 0.001751167, 0.001751147, 0.001751153, 0.001751137, 
    0.001751148, 0.001751135, 0.001751137, 0.00175113, 0.001751132, 
    0.001751122, 0.001751129, 0.001751117, 0.001751124, 0.001751123, 
    0.001751129, 0.001751165, 0.001751158, 0.001751166, 0.001751165, 
    0.001751165, 0.00175117, 0.001751173, 0.001751179, 0.001751178, 
    0.001751174, 0.001751164, 0.001751167, 0.001751159, 0.00175116, 
    0.001751151, 0.001751155, 0.00175114, 0.001751144, 0.001751132, 
    0.001751135, 0.001751132, 0.001751133, 0.001751132, 0.001751136, 
    0.001751134, 0.001751138, 0.001751154, 0.001751149, 0.001751163, 
    0.001751171, 0.001751177, 0.001751181, 0.00175118, 0.001751179, 
    0.001751174, 0.001751169, 0.001751165, 0.001751162, 0.00175116, 
    0.001751152, 0.001751148, 0.001751139, 0.00175114, 0.001751138, 
    0.001751135, 0.001751131, 0.001751131, 0.001751129, 0.001751138, 
    0.001751132, 0.001751141, 0.001751139, 0.001751159, 0.001751167, 
    0.00175117, 0.001751173, 0.00175118, 0.001751175, 0.001751177, 
    0.001751172, 0.001751169, 0.001751171, 0.001751162, 0.001751165, 
    0.001751148, 0.001751155, 0.001751135, 0.00175114, 0.001751134, 
    0.001751137, 0.001751132, 0.001751137, 0.001751129, 0.001751127, 
    0.001751128, 0.001751124, 0.001751137, 0.001751132, 0.001751171, 
    0.001751171, 0.001751169, 0.001751174, 0.001751174, 0.001751179, 
    0.001751175, 0.001751173, 0.001751169, 0.001751167, 0.001751164, 
    0.001751159, 0.001751153, 0.001751146, 0.00175114, 0.001751136, 
    0.001751138, 0.001751136, 0.001751139, 0.00175114, 0.001751128, 
    0.001751134, 0.001751124, 0.001751125, 0.001751129, 0.001751125, 
    0.00175117, 0.001751172, 0.001751176, 0.001751173, 0.001751179, 
    0.001751176, 0.001751174, 0.001751165, 0.001751164, 0.001751162, 
    0.001751159, 0.001751154, 0.001751147, 0.001751141, 0.001751135, 
    0.001751135, 0.001751135, 0.001751134, 0.001751137, 0.001751133, 
    0.001751133, 0.001751134, 0.001751125, 0.001751128, 0.001751125, 
    0.001751127, 0.001751171, 0.001751169, 0.00175117, 0.001751168, 
    0.00175117, 0.001751162, 0.00175116, 0.00175115, 0.001751155, 
    0.001751148, 0.001751154, 0.001751153, 0.001751148, 0.001751154, 
    0.001751141, 0.00175115, 0.001751134, 0.001751142, 0.001751133, 
    0.001751135, 0.001751132, 0.00175113, 0.001751127, 0.001751121, 
    0.001751123, 0.001751118, 0.001751166, 0.001751163, 0.001751163, 
    0.00175116, 0.001751158, 0.001751153, 0.001751145, 0.001751148, 
    0.001751143, 0.001751142, 0.00175115, 0.001751145, 0.001751161, 
    0.001751158, 0.00175116, 0.001751165, 0.001751148, 0.001751157, 
    0.00175114, 0.001751145, 0.00175113, 0.001751137, 0.001751123, 
    0.001751117, 0.001751111, 0.001751105, 0.001751161, 0.001751163, 
    0.00175116, 0.001751155, 0.00175115, 0.001751144, 0.001751144, 
    0.001751143, 0.00175114, 0.001751137, 0.001751142, 0.001751137, 
    0.001751158, 0.001751147, 0.001751164, 0.001751159, 0.001751155, 
    0.001751157, 0.001751148, 0.001751147, 0.001751139, 0.001751143, 
    0.001751119, 0.001751129, 0.0017511, 0.001751108, 0.001751164, 
    0.001751161, 0.001751152, 0.001751157, 0.001751144, 0.001751141, 
    0.001751138, 0.001751135, 0.001751135, 0.001751133, 0.001751136, 
    0.001751133, 0.001751144, 0.001751139, 0.001751153, 0.00175115, 
    0.001751151, 0.001751153, 0.001751148, 0.001751142, 0.001751142, 
    0.00175114, 0.001751135, 0.001751144, 0.001751117, 0.001751134, 
    0.001751158, 0.001751153, 0.001751153, 0.001751155, 0.001751141, 
    0.001751146, 0.001751133, 0.001751137, 0.001751131, 0.001751134, 
    0.001751134, 0.001751138, 0.00175114, 0.001751146, 0.001751151, 
    0.001751154, 0.001751153, 0.001751149, 0.001751142, 0.001751135, 
    0.001751137, 0.001751131, 0.001751145, 0.001751139, 0.001751141, 
    0.001751136, 0.001751148, 0.001751138, 0.001751151, 0.00175115, 
    0.001751146, 0.001751139, 0.001751137, 0.001751135, 0.001751137, 
    0.001751142, 0.001751143, 0.001751146, 0.001751147, 0.00175115, 
    0.001751152, 0.00175115, 0.001751148, 0.001751142, 0.001751136, 
    0.00175113, 0.001751128, 0.001751121, 0.001751127, 0.001751117, 
    0.001751125, 0.001751111, 0.001751137, 0.001751126, 0.001751146, 
    0.001751144, 0.00175114, 0.001751131, 0.001751136, 0.00175113, 
    0.001751143, 0.001751149, 0.001751151, 0.001751154, 0.001751151, 
    0.001751151, 0.001751148, 0.001751149, 0.001751142, 0.001751146, 
    0.001751134, 0.00175113, 0.001751118, 0.001751111, 0.001751104, 
    0.001751101, 0.0017511, 0.001751099,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732905e-07, 9.732868e-07, 9.732875e-07, 9.732845e-07, 9.732862e-07, 
    9.732843e-07, 9.732897e-07, 9.732867e-07, 9.732886e-07, 9.732902e-07, 
    9.732787e-07, 9.732844e-07, 9.732729e-07, 9.732764e-07, 9.732674e-07, 
    9.732735e-07, 9.732662e-07, 9.732677e-07, 9.732635e-07, 9.732647e-07, 
    9.732594e-07, 9.732629e-07, 9.732566e-07, 9.732602e-07, 9.732596e-07, 
    9.73263e-07, 9.732832e-07, 9.732795e-07, 9.732835e-07, 9.732829e-07, 
    9.732831e-07, 9.732861e-07, 9.732877e-07, 9.732908e-07, 9.732902e-07, 
    9.732879e-07, 9.732827e-07, 9.732845e-07, 9.7328e-07, 9.732801e-07, 
    9.732752e-07, 9.732773e-07, 9.73269e-07, 9.732714e-07, 9.732646e-07, 
    9.732663e-07, 9.732647e-07, 9.732652e-07, 9.732647e-07, 9.732672e-07, 
    9.732661e-07, 9.732684e-07, 9.73277e-07, 9.732744e-07, 9.73282e-07, 
    9.732865e-07, 9.732896e-07, 9.732918e-07, 9.732914e-07, 9.732909e-07, 
    9.732879e-07, 9.732851e-07, 9.732829e-07, 9.732815e-07, 9.732801e-07, 
    9.732759e-07, 9.732736e-07, 9.732686e-07, 9.732695e-07, 9.73268e-07, 
    9.732665e-07, 9.73264e-07, 9.732645e-07, 9.732634e-07, 9.73268e-07, 
    9.732649e-07, 9.732701e-07, 9.732686e-07, 9.732797e-07, 9.732839e-07, 
    9.732858e-07, 9.732873e-07, 9.732912e-07, 9.732886e-07, 9.732896e-07, 
    9.732871e-07, 9.732855e-07, 9.732863e-07, 9.732815e-07, 9.732834e-07, 
    9.732735e-07, 9.732778e-07, 9.732667e-07, 9.732693e-07, 9.732661e-07, 
    9.732677e-07, 9.732648e-07, 9.732674e-07, 9.732629e-07, 9.73262e-07, 
    9.732627e-07, 9.732601e-07, 9.732676e-07, 9.732647e-07, 9.732863e-07, 
    9.732862e-07, 9.732856e-07, 9.732883e-07, 9.732884e-07, 9.732908e-07, 
    9.732887e-07, 9.732878e-07, 9.732854e-07, 9.73284e-07, 9.732828e-07, 
    9.7328e-07, 9.732768e-07, 9.732723e-07, 9.732692e-07, 9.73267e-07, 
    9.732684e-07, 9.732672e-07, 9.732685e-07, 9.73269e-07, 9.732623e-07, 
    9.732661e-07, 9.732605e-07, 9.732607e-07, 9.732634e-07, 9.732607e-07, 
    9.732861e-07, 9.732869e-07, 9.732894e-07, 9.732875e-07, 9.732911e-07, 
    9.73289e-07, 9.732878e-07, 9.732834e-07, 9.732823e-07, 9.732814e-07, 
    9.732796e-07, 9.732772e-07, 9.732732e-07, 9.732696e-07, 9.732664e-07, 
    9.732667e-07, 9.732665e-07, 9.732659e-07, 9.732677e-07, 9.732655e-07, 
    9.732652e-07, 9.732661e-07, 9.732609e-07, 9.732623e-07, 9.732607e-07, 
    9.732618e-07, 9.732867e-07, 9.732854e-07, 9.732861e-07, 9.732848e-07, 
    9.732856e-07, 9.732818e-07, 9.732805e-07, 9.732751e-07, 9.732773e-07, 
    9.732737e-07, 9.73277e-07, 9.732764e-07, 9.732736e-07, 9.732768e-07, 
    9.732698e-07, 9.732745e-07, 9.732659e-07, 9.732705e-07, 9.732655e-07, 
    9.732664e-07, 9.732649e-07, 9.732636e-07, 9.732619e-07, 9.732588e-07, 
    9.732595e-07, 9.732569e-07, 9.732836e-07, 9.732819e-07, 9.732821e-07, 
    9.732804e-07, 9.732792e-07, 9.732764e-07, 9.732722e-07, 9.732738e-07, 
    9.732709e-07, 9.732702e-07, 9.732747e-07, 9.73272e-07, 9.732809e-07, 
    9.732794e-07, 9.732803e-07, 9.732834e-07, 9.732735e-07, 9.732786e-07, 
    9.73269e-07, 9.732719e-07, 9.732638e-07, 9.732678e-07, 9.732599e-07, 
    9.732565e-07, 9.732533e-07, 9.732497e-07, 9.732811e-07, 9.732821e-07, 
    9.732802e-07, 9.732775e-07, 9.732751e-07, 9.732717e-07, 9.732713e-07, 
    9.732707e-07, 9.732692e-07, 9.732678e-07, 9.732705e-07, 9.732674e-07, 
    9.73279e-07, 9.73273e-07, 9.732826e-07, 9.732797e-07, 9.732777e-07, 
    9.732786e-07, 9.732739e-07, 9.732729e-07, 9.732686e-07, 9.732707e-07, 
    9.732573e-07, 9.732634e-07, 9.732469e-07, 9.732514e-07, 9.732826e-07, 
    9.732811e-07, 9.73276e-07, 9.732784e-07, 9.732714e-07, 9.732697e-07, 
    9.732684e-07, 9.732667e-07, 9.732664e-07, 9.732654e-07, 9.732671e-07, 
    9.732654e-07, 9.732717e-07, 9.732689e-07, 9.732765e-07, 9.732747e-07, 
    9.732755e-07, 9.732765e-07, 9.732736e-07, 9.732705e-07, 9.732704e-07, 
    9.732694e-07, 9.732667e-07, 9.732714e-07, 9.732566e-07, 9.732657e-07, 
    9.732795e-07, 9.732767e-07, 9.732762e-07, 9.732773e-07, 9.732699e-07, 
    9.732726e-07, 9.732654e-07, 9.732673e-07, 9.732642e-07, 9.732657e-07, 
    9.73266e-07, 9.73268e-07, 9.732693e-07, 9.732724e-07, 9.732751e-07, 
    9.732772e-07, 9.732767e-07, 9.732744e-07, 9.732703e-07, 9.732664e-07, 
    9.732672e-07, 9.732644e-07, 9.73272e-07, 9.732688e-07, 9.732701e-07, 
    9.732669e-07, 9.732738e-07, 9.732679e-07, 9.732754e-07, 9.732747e-07, 
    9.732727e-07, 9.732686e-07, 9.732677e-07, 9.732668e-07, 9.732673e-07, 
    9.732702e-07, 9.732706e-07, 9.732727e-07, 9.732732e-07, 9.732748e-07, 
    9.732762e-07, 9.73275e-07, 9.732737e-07, 9.732702e-07, 9.73267e-07, 
    9.732636e-07, 9.732627e-07, 9.732587e-07, 9.73262e-07, 9.732565e-07, 
    9.732612e-07, 9.732532e-07, 9.732676e-07, 9.732613e-07, 9.732726e-07, 
    9.732713e-07, 9.732692e-07, 9.732642e-07, 9.732669e-07, 9.732637e-07, 
    9.732707e-07, 9.732744e-07, 9.732753e-07, 9.732771e-07, 9.732753e-07, 
    9.732754e-07, 9.732737e-07, 9.732743e-07, 9.732701e-07, 9.732723e-07, 
    9.73266e-07, 9.732637e-07, 9.732572e-07, 9.732532e-07, 9.732491e-07, 
    9.732474e-07, 9.732469e-07, 9.732466e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  4.215557e-25, -2.254833e-25, 6.862535e-26, -6.47039e-25, 2.450906e-25, 
    2.695996e-25, -1.470543e-25, 1.666616e-25, 2.254833e-25, 1.911706e-25, 
    -1.470543e-26, 1.078398e-25, -3.333231e-25, -4.019485e-25, -3.431268e-25, 
    -2.843051e-25, 8.333079e-26, -5.931191e-25, -9.803622e-26, 5.98021e-25, 
    -3.039123e-25, -7.842898e-26, 1.862688e-25, -2.156797e-25, -4.313593e-25, 
    7.646825e-25, -2.843051e-25, -3.921449e-26, -1.470543e-25, 1.078398e-25, 
    -8.333079e-25, 6.568427e-25, -9.313441e-25, 1.372507e-25, 1.666616e-25, 
    -6.2253e-25, 2.009742e-25, 2.009742e-25, 1.372507e-25, 4.607703e-25, 
    -2.646978e-25, -5.391992e-25, 7.352717e-25, 1.102908e-24, 1.764652e-25, 
    -3.137159e-25, 3.725376e-25, -1.078398e-25, -2.843051e-25, 4.901811e-25, 
    -6.862535e-25, -3.725376e-25, -1.176435e-25, 9.999695e-25, 7.352717e-26, 
    -2.941087e-26, 2.058761e-25, -2.941087e-26, -5.244938e-25, 3.235195e-25, 
    7.25468e-25, -1.764652e-25, 4.705739e-25, -6.127264e-25, 9.068351e-25, 
    7.156644e-25, 7.156644e-25, 1.56858e-25, 1.156827e-24, 9.999695e-25, 
    -8.82326e-26, 2.892069e-25, 4.41163e-25, 2.990105e-25, 1.960724e-25, 
    5.882173e-25, 6.078246e-25, -3.431268e-26, 4.313593e-25, 5.882173e-25, 
    -7.107626e-25, 6.764499e-25, -6.519409e-25, 1.960724e-26, -1.81367e-25, 
    -4.705739e-25, 3.333231e-25, 2.303851e-25, 5.048866e-25, -5.686101e-25, 
    6.47039e-25, 1.009773e-24, -1.274471e-25, 3.480286e-25, 6.862535e-25, 
    6.911554e-25, 3.970467e-25, -5.490028e-25, -4.607703e-25, -9.803622e-26, 
    3.921449e-25, 2.450906e-25, 4.803775e-25, 1.176435e-25, 5.98021e-25, 
    3.38225e-25, 1.274471e-25, 5.490028e-25, -7.842898e-26, 5.490028e-25, 
    -2.695996e-25, 1.960724e-26, 5.097883e-25, 2.646978e-25, 6.862535e-26, 
    -2.941087e-26, -2.352869e-25, -2.794032e-25, 4.117521e-25, -3.970467e-25, 
    -3.774394e-25, 3.186177e-25, 3.725376e-25, 1.960724e-25, 3.529304e-25, 
    -4.215557e-25, 3.921449e-25, 9.019333e-25, 1.519561e-25, -2.156797e-25, 
    -3.431268e-25, 5.097883e-25, 6.764499e-25, 6.813517e-25, 6.078246e-25, 
    7.303698e-25, -8.529151e-25, -1.56858e-25, 4.558684e-25, -1.274471e-25, 
    4.313593e-25, 6.862535e-26, -1.176435e-25, 2.450905e-26, 1.078398e-25, 
    -4.41163e-25, 4.117521e-25, 7.058608e-25, -1.960724e-26, 8.529151e-25, 
    -1.02938e-25, 6.568427e-25, -3.333231e-25, 4.999847e-25, 6.568427e-25, 
    2.646978e-25, 3.921449e-26, 1.274471e-25, 4.509666e-25, -2.941087e-26, 
    4.509666e-25, 3.725376e-25, -3.62734e-25, 3.725376e-25, -3.431268e-26, 
    -2.941087e-25, 9.411477e-25, 6.47039e-25, -3.137159e-25, -1.862688e-25, 
    -3.578322e-25, 6.764499e-25, 5.19592e-25, 9.313441e-25, -4.705739e-25, 
    -7.842898e-26, 4.313593e-25, -3.137159e-25, 7.205662e-25, -7.842898e-26, 
    -1.470543e-25, -3.529304e-25, -1.911706e-25, 4.117521e-25, -4.215557e-25, 
    4.901811e-26, -7.842898e-26, 2.254833e-25, -2.107779e-25, 7.695843e-25, 
    1.323489e-25, 4.117521e-25, 1.470543e-26, 2.450905e-26, -4.607703e-25, 
    2.745014e-25, -3.970467e-25, -2.59796e-25, 3.431268e-26, -3.774394e-25, 
    -7.156644e-25, -3.039123e-25, -8.82326e-26, -7.450753e-25, 3.676358e-25, 
    3.480286e-25, 9.803622e-26, 4.117521e-25, 2.548942e-25, 1.862688e-25, 
    3.333231e-25, 4.65672e-25, -1.225453e-25, -3.529304e-25, 1.960724e-26, 
    8.82326e-26, -8.333079e-26, 5.882173e-26, -2.156797e-25, -2.548942e-25, 
    7.058608e-25, -1.014675e-24, 3.725376e-25, 2.794032e-25, -1.176435e-25, 
    7.352717e-25, -8.382097e-25, 7.842898e-26, -2.205815e-25, 3.529304e-25, 
    1.666616e-25, 1.372507e-25, 5.98021e-25, 5.784137e-25, 3.431268e-25, 
    4.068503e-25, -1.519561e-25, -5.391992e-26, -3.431268e-26, 1.960724e-26, 
    5.833155e-25, 6.2253e-25, -1.666616e-25, 4.215557e-25, -4.264576e-25, 
    4.41163e-25, -1.911706e-25, 2.254833e-25, -3.872431e-25, -4.901811e-26, 
    -7.842898e-26, -4.215557e-25, -7.401734e-25, 5.784137e-25, 2.695996e-25, 
    -2.892069e-25, -1.56858e-25, 1.960724e-25, 3.235195e-25, -3.921449e-25, 
    4.558684e-25, -6.862535e-26, 4.607703e-25, -4.65672e-25, 4.019485e-25, 
    -3.921449e-25, 1.274471e-25, 6.666463e-25, 1.862688e-25, 6.421373e-25, 
    2.548942e-25, 1.176435e-24, 1.078398e-25, 5.342974e-25, -1.225453e-25, 
    1.862688e-25, 7.107626e-25, 9.803622e-27, -3.431268e-25, -3.235195e-25, 
    7.597807e-25, 4.999847e-25, 5.882173e-25, -3.921449e-25, 1.764652e-25, 
    -5.882173e-25, 1.078398e-25, -6.372354e-26, -3.039123e-25, 3.333231e-25, 
    3.921449e-25, -1.960724e-25, 8.82326e-26, -6.862535e-26, 4.019485e-25, 
    5.293956e-25, -3.676358e-25, -1.862688e-25, 3.970467e-25, 1.666616e-25, 
    -1.323489e-25, -1.56858e-25, 1.02938e-24, -6.372354e-26, -3.431268e-25, 
    3.039123e-25, -2.450905e-26, 7.597807e-25, 7.842898e-25, -5.588064e-25, 
    -1.274471e-25, 3.284213e-25, 2.156797e-25, -3.823413e-25, -6.862535e-26, 
    -7.842898e-26, 1.862688e-25, -1.044086e-24, -6.862535e-25, -8.82326e-26, 
    1.176435e-25, 3.039123e-25, 8.137007e-25, 6.421373e-25, -2.548942e-25, 
    1.205845e-24, 4.509666e-25, 5.097883e-25, 1.372507e-25, 3.431268e-26, 
    -1.56858e-25, -3.921449e-25, 9.019333e-25, 6.372354e-26, 3.431268e-25, 
    6.176282e-25, 3.823413e-25, 1.862688e-25,
  9.436745e-32, 9.436708e-32, 9.436715e-32, 9.436685e-32, 9.436702e-32, 
    9.436682e-32, 9.436738e-32, 9.436706e-32, 9.436726e-32, 9.436742e-32, 
    9.436626e-32, 9.436684e-32, 9.436568e-32, 9.436604e-32, 9.436513e-32, 
    9.436574e-32, 9.436501e-32, 9.436515e-32, 9.436473e-32, 9.436485e-32, 
    9.436432e-32, 9.436468e-32, 9.436404e-32, 9.436441e-32, 9.436435e-32, 
    9.436469e-32, 9.436672e-32, 9.436634e-32, 9.436674e-32, 9.436669e-32, 
    9.436671e-32, 9.436701e-32, 9.436716e-32, 9.436748e-32, 9.436742e-32, 
    9.436719e-32, 9.436666e-32, 9.436684e-32, 9.436639e-32, 9.436641e-32, 
    9.436591e-32, 9.436613e-32, 9.43653e-32, 9.436553e-32, 9.436485e-32, 
    9.436502e-32, 9.436485e-32, 9.436491e-32, 9.436485e-32, 9.436511e-32, 
    9.4365e-32, 9.436522e-32, 9.436609e-32, 9.436584e-32, 9.436659e-32, 
    9.436705e-32, 9.436736e-32, 9.436758e-32, 9.436755e-32, 9.436749e-32, 
    9.436719e-32, 9.436691e-32, 9.436669e-32, 9.436655e-32, 9.436641e-32, 
    9.436598e-32, 9.436575e-32, 9.436525e-32, 9.436534e-32, 9.436518e-32, 
    9.436504e-32, 9.436479e-32, 9.436483e-32, 9.436472e-32, 9.436519e-32, 
    9.436488e-32, 9.436539e-32, 9.436525e-32, 9.436637e-32, 9.436679e-32, 
    9.436698e-32, 9.436713e-32, 9.436752e-32, 9.436725e-32, 9.436736e-32, 
    9.436711e-32, 9.436695e-32, 9.436703e-32, 9.436654e-32, 9.436673e-32, 
    9.436574e-32, 9.436617e-32, 9.436505e-32, 9.436532e-32, 9.436499e-32, 
    9.436516e-32, 9.436487e-32, 9.436513e-32, 9.436468e-32, 9.436458e-32, 
    9.436465e-32, 9.43644e-32, 9.436514e-32, 9.436485e-32, 9.436703e-32, 
    9.436702e-32, 9.436696e-32, 9.436722e-32, 9.436723e-32, 9.436748e-32, 
    9.436726e-32, 9.436717e-32, 9.436694e-32, 9.436681e-32, 9.436668e-32, 
    9.436639e-32, 9.436607e-32, 9.436562e-32, 9.43653e-32, 9.436509e-32, 
    9.436522e-32, 9.436511e-32, 9.436524e-32, 9.43653e-32, 9.436462e-32, 
    9.4365e-32, 9.436443e-32, 9.436446e-32, 9.436472e-32, 9.436446e-32, 
    9.436701e-32, 9.436708e-32, 9.436734e-32, 9.436714e-32, 9.436751e-32, 
    9.43673e-32, 9.436718e-32, 9.436673e-32, 9.436663e-32, 9.436654e-32, 
    9.436635e-32, 9.436612e-32, 9.436571e-32, 9.436535e-32, 9.436503e-32, 
    9.436505e-32, 9.436504e-32, 9.436497e-32, 9.436515e-32, 9.436494e-32, 
    9.436491e-32, 9.4365e-32, 9.436447e-32, 9.436462e-32, 9.436446e-32, 
    9.436456e-32, 9.436706e-32, 9.436693e-32, 9.4367e-32, 9.436688e-32, 
    9.436696e-32, 9.436657e-32, 9.436645e-32, 9.436589e-32, 9.436612e-32, 
    9.436577e-32, 9.436609e-32, 9.436603e-32, 9.436575e-32, 9.436607e-32, 
    9.436537e-32, 9.436585e-32, 9.436497e-32, 9.436544e-32, 9.436494e-32, 
    9.436503e-32, 9.436488e-32, 9.436474e-32, 9.436458e-32, 9.436427e-32, 
    9.436434e-32, 9.436407e-32, 9.436675e-32, 9.436659e-32, 9.43666e-32, 
    9.436644e-32, 9.436631e-32, 9.436604e-32, 9.436561e-32, 9.436577e-32, 
    9.436547e-32, 9.436541e-32, 9.436587e-32, 9.436559e-32, 9.436648e-32, 
    9.436634e-32, 9.436642e-32, 9.436674e-32, 9.436574e-32, 9.436625e-32, 
    9.43653e-32, 9.436558e-32, 9.436477e-32, 9.436517e-32, 9.436438e-32, 
    9.436404e-32, 9.436372e-32, 9.436335e-32, 9.43665e-32, 9.436661e-32, 
    9.436641e-32, 9.436614e-32, 9.436589e-32, 9.436556e-32, 9.436552e-32, 
    9.436547e-32, 9.43653e-32, 9.436517e-32, 9.436544e-32, 9.436513e-32, 
    9.43663e-32, 9.436569e-32, 9.436665e-32, 9.436636e-32, 9.436616e-32, 
    9.436625e-32, 9.436579e-32, 9.436568e-32, 9.436524e-32, 9.436547e-32, 
    9.436412e-32, 9.436472e-32, 9.436307e-32, 9.436353e-32, 9.436665e-32, 
    9.43665e-32, 9.436599e-32, 9.436624e-32, 9.436554e-32, 9.436537e-32, 
    9.436522e-32, 9.436505e-32, 9.436503e-32, 9.436492e-32, 9.43651e-32, 
    9.436493e-32, 9.436556e-32, 9.436528e-32, 9.436605e-32, 9.436586e-32, 
    9.436595e-32, 9.436604e-32, 9.436575e-32, 9.436544e-32, 9.436543e-32, 
    9.436533e-32, 9.436505e-32, 9.436554e-32, 9.436404e-32, 9.436497e-32, 
    9.436634e-32, 9.436606e-32, 9.436602e-32, 9.436612e-32, 9.436538e-32, 
    9.436565e-32, 9.436493e-32, 9.436512e-32, 9.43648e-32, 9.436496e-32, 
    9.436498e-32, 9.436519e-32, 9.436532e-32, 9.436564e-32, 9.43659e-32, 
    9.436611e-32, 9.436607e-32, 9.436584e-32, 9.436542e-32, 9.436503e-32, 
    9.436511e-32, 9.436482e-32, 9.436559e-32, 9.436527e-32, 9.436539e-32, 
    9.436507e-32, 9.436578e-32, 9.436518e-32, 9.436593e-32, 9.436586e-32, 
    9.436566e-32, 9.436525e-32, 9.436515e-32, 9.436506e-32, 9.436512e-32, 
    9.436541e-32, 9.436546e-32, 9.436567e-32, 9.436572e-32, 9.436588e-32, 
    9.436601e-32, 9.436589e-32, 9.436577e-32, 9.436541e-32, 9.436509e-32, 
    9.436474e-32, 9.436466e-32, 9.436425e-32, 9.436458e-32, 9.436404e-32, 
    9.43645e-32, 9.43637e-32, 9.436514e-32, 9.436451e-32, 9.436565e-32, 
    9.436552e-32, 9.436531e-32, 9.43648e-32, 9.436507e-32, 9.436475e-32, 
    9.436546e-32, 9.436582e-32, 9.436592e-32, 9.43661e-32, 9.436592e-32, 
    9.436593e-32, 9.436576e-32, 9.436581e-32, 9.43654e-32, 9.436562e-32, 
    9.436498e-32, 9.436475e-32, 9.43641e-32, 9.43637e-32, 9.43633e-32, 
    9.436312e-32, 9.436306e-32, 9.436304e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.031324e-14, 4.042231e-14, 4.040113e-14, 4.048902e-14, 4.044029e-14, 
    4.049781e-14, 4.033538e-14, 4.042663e-14, 4.036839e-14, 4.032309e-14, 
    4.065933e-14, 4.049294e-14, 4.083204e-14, 4.07261e-14, 4.099203e-14, 
    4.081554e-14, 4.102759e-14, 4.098698e-14, 4.110926e-14, 4.107425e-14, 
    4.123041e-14, 4.112541e-14, 4.131132e-14, 4.120536e-14, 4.122193e-14, 
    4.112195e-14, 4.052648e-14, 4.063862e-14, 4.051983e-14, 4.053583e-14, 
    4.052866e-14, 4.044128e-14, 4.03972e-14, 4.030492e-14, 4.032169e-14, 
    4.038947e-14, 4.054302e-14, 4.049095e-14, 4.062221e-14, 4.061925e-14, 
    4.076517e-14, 4.06994e-14, 4.094436e-14, 4.087482e-14, 4.107571e-14, 
    4.102521e-14, 4.107333e-14, 4.105875e-14, 4.107352e-14, 4.099946e-14, 
    4.103119e-14, 4.096601e-14, 4.071172e-14, 4.078651e-14, 4.056326e-14, 
    4.042873e-14, 4.033938e-14, 4.02759e-14, 4.028487e-14, 4.030198e-14, 
    4.038987e-14, 4.047247e-14, 4.053536e-14, 4.057741e-14, 4.061882e-14, 
    4.074399e-14, 4.081026e-14, 4.09584e-14, 4.093171e-14, 4.097695e-14, 
    4.102019e-14, 4.109271e-14, 4.108078e-14, 4.111271e-14, 4.097578e-14, 
    4.106679e-14, 4.091652e-14, 4.095762e-14, 4.062995e-14, 4.0505e-14, 
    4.045174e-14, 4.04052e-14, 4.029177e-14, 4.037011e-14, 4.033923e-14, 
    4.04127e-14, 4.045934e-14, 4.043628e-14, 4.057856e-14, 4.052326e-14, 
    4.081418e-14, 4.068898e-14, 4.101515e-14, 4.093719e-14, 4.103383e-14, 
    4.098454e-14, 4.106897e-14, 4.099298e-14, 4.11246e-14, 4.115322e-14, 
    4.113366e-14, 4.120883e-14, 4.098876e-14, 4.107332e-14, 4.043562e-14, 
    4.043939e-14, 4.045692e-14, 4.037983e-14, 4.037512e-14, 4.030446e-14, 
    4.036734e-14, 4.03941e-14, 4.046205e-14, 4.050219e-14, 4.054035e-14, 
    4.06242e-14, 4.071775e-14, 4.084845e-14, 4.094225e-14, 4.100508e-14, 
    4.096656e-14, 4.100057e-14, 4.096255e-14, 4.094473e-14, 4.114249e-14, 
    4.103148e-14, 4.119802e-14, 4.118882e-14, 4.111346e-14, 4.118985e-14, 
    4.044203e-14, 4.042038e-14, 4.034516e-14, 4.040403e-14, 4.029677e-14, 
    4.035681e-14, 4.03913e-14, 4.052439e-14, 4.055364e-14, 4.058071e-14, 
    4.063419e-14, 4.070277e-14, 4.082296e-14, 4.092741e-14, 4.102271e-14, 
    4.101573e-14, 4.101819e-14, 4.103945e-14, 4.098675e-14, 4.10481e-14, 
    4.105839e-14, 4.103149e-14, 4.118758e-14, 4.114301e-14, 4.118862e-14, 
    4.115961e-14, 4.042742e-14, 4.046384e-14, 4.044416e-14, 4.048116e-14, 
    4.045509e-14, 4.057095e-14, 4.060565e-14, 4.076796e-14, 4.070141e-14, 
    4.080734e-14, 4.071219e-14, 4.072905e-14, 4.081074e-14, 4.071734e-14, 
    4.092165e-14, 4.078313e-14, 4.104028e-14, 4.090209e-14, 4.104893e-14, 
    4.10223e-14, 4.106641e-14, 4.110588e-14, 4.115554e-14, 4.124707e-14, 
    4.122589e-14, 4.13024e-14, 4.051813e-14, 4.056532e-14, 4.056119e-14, 
    4.061056e-14, 4.064706e-14, 4.072615e-14, 4.085284e-14, 4.080522e-14, 
    4.089265e-14, 4.091018e-14, 4.077737e-14, 4.085891e-14, 4.05969e-14, 
    4.063925e-14, 4.061405e-14, 4.052184e-14, 4.081617e-14, 4.06652e-14, 
    4.094379e-14, 4.086217e-14, 4.110025e-14, 4.098188e-14, 4.121422e-14, 
    4.131331e-14, 4.14066e-14, 4.151537e-14, 4.059108e-14, 4.055903e-14, 
    4.061644e-14, 4.069577e-14, 4.076939e-14, 4.086714e-14, 4.087715e-14, 
    4.089545e-14, 4.094283e-14, 4.098265e-14, 4.090121e-14, 4.099264e-14, 
    4.064902e-14, 4.082927e-14, 4.054688e-14, 4.063197e-14, 4.069111e-14, 
    4.066519e-14, 4.079978e-14, 4.083147e-14, 4.096011e-14, 4.089366e-14, 
    4.128884e-14, 4.111418e-14, 4.159819e-14, 4.146316e-14, 4.054782e-14, 
    4.059098e-14, 4.074103e-14, 4.066967e-14, 4.087368e-14, 4.092382e-14, 
    4.096457e-14, 4.101662e-14, 4.102225e-14, 4.105308e-14, 4.100255e-14, 
    4.105109e-14, 4.086735e-14, 4.09495e-14, 4.072392e-14, 4.077886e-14, 
    4.07536e-14, 4.072586e-14, 4.081143e-14, 4.090249e-14, 4.090447e-14, 
    4.093362e-14, 4.101571e-14, 4.087451e-14, 4.131129e-14, 4.104168e-14, 
    4.063803e-14, 4.072103e-14, 4.073292e-14, 4.070077e-14, 4.09188e-14, 
    4.083985e-14, 4.105233e-14, 4.099495e-14, 4.108897e-14, 4.104226e-14, 
    4.103538e-14, 4.097536e-14, 4.093797e-14, 4.084346e-14, 4.07665e-14, 
    4.070544e-14, 4.071965e-14, 4.07867e-14, 4.090806e-14, 4.102274e-14, 
    4.099762e-14, 4.108182e-14, 4.08589e-14, 4.09524e-14, 4.091627e-14, 
    4.101049e-14, 4.080395e-14, 4.097974e-14, 4.075895e-14, 4.077833e-14, 
    4.083828e-14, 4.095872e-14, 4.09854e-14, 4.101382e-14, 4.09963e-14, 
    4.091115e-14, 4.08972e-14, 4.083683e-14, 4.082014e-14, 4.077412e-14, 
    4.073598e-14, 4.077082e-14, 4.080738e-14, 4.09112e-14, 4.100463e-14, 
    4.110643e-14, 4.113135e-14, 4.125004e-14, 4.115338e-14, 4.131278e-14, 
    4.117719e-14, 4.141183e-14, 4.098997e-14, 4.117328e-14, 4.084102e-14, 
    4.087688e-14, 4.094164e-14, 4.109016e-14, 4.101005e-14, 4.110375e-14, 
    4.089666e-14, 4.078899e-14, 4.076117e-14, 4.070915e-14, 4.076236e-14, 
    4.075803e-14, 4.080892e-14, 4.079257e-14, 4.091465e-14, 4.084909e-14, 
    4.10352e-14, 4.110302e-14, 4.129437e-14, 4.141147e-14, 4.153058e-14, 
    4.15831e-14, 4.159909e-14, 4.160576e-14 ;

 LITR1N_vr =
  5.557589e-05, 5.557568e-05, 5.557572e-05, 5.557555e-05, 5.557565e-05, 
    5.557554e-05, 5.557585e-05, 5.557567e-05, 5.557579e-05, 5.557587e-05, 
    5.557522e-05, 5.557554e-05, 5.557489e-05, 5.557509e-05, 5.557458e-05, 
    5.557492e-05, 5.557451e-05, 5.557459e-05, 5.557435e-05, 5.557442e-05, 
    5.557411e-05, 5.557432e-05, 5.557396e-05, 5.557416e-05, 5.557413e-05, 
    5.557432e-05, 5.557548e-05, 5.557526e-05, 5.557549e-05, 5.557546e-05, 
    5.557547e-05, 5.557565e-05, 5.557573e-05, 5.557591e-05, 5.557588e-05, 
    5.557575e-05, 5.557545e-05, 5.557555e-05, 5.55753e-05, 5.55753e-05, 
    5.557502e-05, 5.557514e-05, 5.557467e-05, 5.55748e-05, 5.557442e-05, 
    5.557451e-05, 5.557442e-05, 5.557445e-05, 5.557442e-05, 5.557456e-05, 
    5.55745e-05, 5.557463e-05, 5.557512e-05, 5.557498e-05, 5.557541e-05, 
    5.557567e-05, 5.557584e-05, 5.557597e-05, 5.557595e-05, 5.557591e-05, 
    5.557574e-05, 5.557558e-05, 5.557546e-05, 5.557538e-05, 5.55753e-05, 
    5.557506e-05, 5.557493e-05, 5.557464e-05, 5.55747e-05, 5.557461e-05, 
    5.557452e-05, 5.557438e-05, 5.55744e-05, 5.557434e-05, 5.557461e-05, 
    5.557443e-05, 5.557472e-05, 5.557464e-05, 5.557528e-05, 5.557552e-05, 
    5.557562e-05, 5.557571e-05, 5.557594e-05, 5.557578e-05, 5.557584e-05, 
    5.55757e-05, 5.557561e-05, 5.557566e-05, 5.557538e-05, 5.557549e-05, 
    5.557492e-05, 5.557516e-05, 5.557453e-05, 5.557468e-05, 5.55745e-05, 
    5.557459e-05, 5.557443e-05, 5.557458e-05, 5.557432e-05, 5.557427e-05, 
    5.55743e-05, 5.557416e-05, 5.557458e-05, 5.557442e-05, 5.557566e-05, 
    5.557565e-05, 5.557562e-05, 5.557577e-05, 5.557577e-05, 5.557591e-05, 
    5.557579e-05, 5.557574e-05, 5.557561e-05, 5.557553e-05, 5.557545e-05, 
    5.557529e-05, 5.557511e-05, 5.557486e-05, 5.557467e-05, 5.557455e-05, 
    5.557463e-05, 5.557456e-05, 5.557463e-05, 5.557467e-05, 5.557428e-05, 
    5.55745e-05, 5.557418e-05, 5.55742e-05, 5.557434e-05, 5.557419e-05, 
    5.557565e-05, 5.557569e-05, 5.557583e-05, 5.557572e-05, 5.557593e-05, 
    5.557581e-05, 5.557574e-05, 5.557549e-05, 5.557543e-05, 5.557538e-05, 
    5.557527e-05, 5.557514e-05, 5.557491e-05, 5.55747e-05, 5.557452e-05, 
    5.557453e-05, 5.557453e-05, 5.557448e-05, 5.557459e-05, 5.557447e-05, 
    5.557445e-05, 5.55745e-05, 5.55742e-05, 5.557428e-05, 5.55742e-05, 
    5.557425e-05, 5.557567e-05, 5.55756e-05, 5.557564e-05, 5.557557e-05, 
    5.557562e-05, 5.557539e-05, 5.557532e-05, 5.557501e-05, 5.557514e-05, 
    5.557494e-05, 5.557512e-05, 5.557509e-05, 5.557493e-05, 5.557511e-05, 
    5.557471e-05, 5.557498e-05, 5.557448e-05, 5.557475e-05, 5.557447e-05, 
    5.557452e-05, 5.557443e-05, 5.557436e-05, 5.557426e-05, 5.557408e-05, 
    5.557412e-05, 5.557398e-05, 5.55755e-05, 5.55754e-05, 5.557541e-05, 
    5.557532e-05, 5.557524e-05, 5.557509e-05, 5.557485e-05, 5.557494e-05, 
    5.557477e-05, 5.557474e-05, 5.557499e-05, 5.557483e-05, 5.557534e-05, 
    5.557526e-05, 5.557531e-05, 5.557549e-05, 5.557492e-05, 5.557521e-05, 
    5.557467e-05, 5.557483e-05, 5.557437e-05, 5.55746e-05, 5.557415e-05, 
    5.557395e-05, 5.557378e-05, 5.557356e-05, 5.557535e-05, 5.557542e-05, 
    5.557531e-05, 5.557515e-05, 5.557501e-05, 5.557482e-05, 5.55748e-05, 
    5.557476e-05, 5.557467e-05, 5.557459e-05, 5.557475e-05, 5.557458e-05, 
    5.557524e-05, 5.557489e-05, 5.557544e-05, 5.557527e-05, 5.557516e-05, 
    5.557521e-05, 5.557495e-05, 5.557489e-05, 5.557464e-05, 5.557477e-05, 
    5.5574e-05, 5.557434e-05, 5.55734e-05, 5.557367e-05, 5.557544e-05, 
    5.557535e-05, 5.557506e-05, 5.55752e-05, 5.557481e-05, 5.557471e-05, 
    5.557463e-05, 5.557453e-05, 5.557452e-05, 5.557446e-05, 5.557456e-05, 
    5.557446e-05, 5.557482e-05, 5.557466e-05, 5.55751e-05, 5.557499e-05, 
    5.557504e-05, 5.557509e-05, 5.557493e-05, 5.557475e-05, 5.557475e-05, 
    5.557469e-05, 5.557453e-05, 5.55748e-05, 5.557396e-05, 5.557448e-05, 
    5.557526e-05, 5.55751e-05, 5.557508e-05, 5.557514e-05, 5.557472e-05, 
    5.557487e-05, 5.557446e-05, 5.557457e-05, 5.557439e-05, 5.557448e-05, 
    5.557449e-05, 5.557461e-05, 5.557468e-05, 5.557487e-05, 5.557502e-05, 
    5.557513e-05, 5.557511e-05, 5.557498e-05, 5.557474e-05, 5.557452e-05, 
    5.557456e-05, 5.55744e-05, 5.557483e-05, 5.557466e-05, 5.557472e-05, 
    5.557454e-05, 5.557494e-05, 5.55746e-05, 5.557503e-05, 5.557499e-05, 
    5.557487e-05, 5.557464e-05, 5.557459e-05, 5.557454e-05, 5.557457e-05, 
    5.557474e-05, 5.557476e-05, 5.557488e-05, 5.557491e-05, 5.5575e-05, 
    5.557507e-05, 5.5575e-05, 5.557494e-05, 5.557474e-05, 5.557455e-05, 
    5.557436e-05, 5.557431e-05, 5.557408e-05, 5.557427e-05, 5.557396e-05, 
    5.557422e-05, 5.557376e-05, 5.557458e-05, 5.557423e-05, 5.557487e-05, 
    5.55748e-05, 5.557467e-05, 5.557439e-05, 5.557454e-05, 5.557436e-05, 
    5.557476e-05, 5.557497e-05, 5.557502e-05, 5.557512e-05, 5.557502e-05, 
    5.557503e-05, 5.557493e-05, 5.557496e-05, 5.557473e-05, 5.557486e-05, 
    5.557449e-05, 5.557436e-05, 5.557399e-05, 5.557376e-05, 5.557354e-05, 
    5.557343e-05, 5.55734e-05, 5.557339e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  6.986438e-13, 7.005341e-13, 7.001669e-13, 7.016901e-13, 7.008456e-13, 
    7.018426e-13, 6.990275e-13, 7.006089e-13, 6.995997e-13, 6.988145e-13, 
    7.046417e-13, 7.017581e-13, 7.076347e-13, 7.057989e-13, 7.104075e-13, 
    7.073488e-13, 7.110239e-13, 7.1032e-13, 7.124392e-13, 7.118323e-13, 
    7.145386e-13, 7.127191e-13, 7.15941e-13, 7.141047e-13, 7.143918e-13, 
    7.12659e-13, 7.023394e-13, 7.042827e-13, 7.02224e-13, 7.025014e-13, 
    7.023771e-13, 7.008628e-13, 7.000988e-13, 6.984997e-13, 6.987903e-13, 
    6.999649e-13, 7.026261e-13, 7.017236e-13, 7.039984e-13, 7.039471e-13, 
    7.064759e-13, 7.053362e-13, 7.095814e-13, 7.083762e-13, 7.118577e-13, 
    7.109826e-13, 7.118165e-13, 7.115637e-13, 7.118198e-13, 7.105362e-13, 
    7.110862e-13, 7.099566e-13, 7.055496e-13, 7.068458e-13, 7.029767e-13, 
    7.006453e-13, 6.990968e-13, 6.979967e-13, 6.981523e-13, 6.984486e-13, 
    6.999718e-13, 7.014033e-13, 7.024933e-13, 7.032219e-13, 7.039397e-13, 
    7.061089e-13, 7.072573e-13, 7.098247e-13, 7.093621e-13, 7.101461e-13, 
    7.108955e-13, 7.121523e-13, 7.119456e-13, 7.12499e-13, 7.101258e-13, 
    7.117032e-13, 7.090988e-13, 7.098112e-13, 7.041326e-13, 7.019672e-13, 
    7.010441e-13, 7.002374e-13, 6.982718e-13, 6.996293e-13, 6.990943e-13, 
    7.003674e-13, 7.011757e-13, 7.007761e-13, 7.032419e-13, 7.022836e-13, 
    7.073254e-13, 7.051554e-13, 7.108081e-13, 7.094571e-13, 7.111319e-13, 
    7.102776e-13, 7.117409e-13, 7.10424e-13, 7.12705e-13, 7.13201e-13, 
    7.128621e-13, 7.141647e-13, 7.103509e-13, 7.118163e-13, 7.007648e-13, 
    7.0083e-13, 7.011338e-13, 6.997978e-13, 6.997162e-13, 6.984917e-13, 
    6.995815e-13, 7.000452e-13, 7.012227e-13, 7.019185e-13, 7.025798e-13, 
    7.04033e-13, 7.056541e-13, 7.079192e-13, 7.095447e-13, 7.106336e-13, 
    7.099662e-13, 7.105555e-13, 7.098966e-13, 7.095878e-13, 7.130151e-13, 
    7.110912e-13, 7.139774e-13, 7.138179e-13, 7.12512e-13, 7.138359e-13, 
    7.008758e-13, 7.005006e-13, 6.99197e-13, 7.002173e-13, 6.983583e-13, 
    6.993988e-13, 6.999967e-13, 7.023031e-13, 7.0281e-13, 7.032792e-13, 
    7.042061e-13, 7.053945e-13, 7.074774e-13, 7.092876e-13, 7.109392e-13, 
    7.108183e-13, 7.108608e-13, 7.112294e-13, 7.103161e-13, 7.113793e-13, 
    7.115575e-13, 7.110912e-13, 7.137965e-13, 7.130241e-13, 7.138145e-13, 
    7.133117e-13, 7.006227e-13, 7.012538e-13, 7.009127e-13, 7.01554e-13, 
    7.011021e-13, 7.031099e-13, 7.037115e-13, 7.065243e-13, 7.05371e-13, 
    7.072068e-13, 7.055577e-13, 7.058499e-13, 7.072657e-13, 7.05647e-13, 
    7.091878e-13, 7.067872e-13, 7.112437e-13, 7.088487e-13, 7.113937e-13, 
    7.109321e-13, 7.116965e-13, 7.123806e-13, 7.132412e-13, 7.148274e-13, 
    7.144603e-13, 7.157864e-13, 7.021946e-13, 7.030124e-13, 7.029408e-13, 
    7.037965e-13, 7.04429e-13, 7.057996e-13, 7.079953e-13, 7.071701e-13, 
    7.086852e-13, 7.089891e-13, 7.066874e-13, 7.081005e-13, 7.035598e-13, 
    7.042937e-13, 7.038571e-13, 7.022589e-13, 7.073597e-13, 7.047435e-13, 
    7.095715e-13, 7.081569e-13, 7.12283e-13, 7.102316e-13, 7.142581e-13, 
    7.159755e-13, 7.175922e-13, 7.194772e-13, 7.034589e-13, 7.029034e-13, 
    7.038984e-13, 7.052732e-13, 7.06549e-13, 7.082432e-13, 7.084167e-13, 
    7.087337e-13, 7.095548e-13, 7.10245e-13, 7.088335e-13, 7.104181e-13, 
    7.044631e-13, 7.075868e-13, 7.02693e-13, 7.041675e-13, 7.051924e-13, 
    7.047433e-13, 7.070758e-13, 7.07625e-13, 7.098544e-13, 7.087027e-13, 
    7.155514e-13, 7.125244e-13, 7.209125e-13, 7.185723e-13, 7.027092e-13, 
    7.034573e-13, 7.060576e-13, 7.048209e-13, 7.083564e-13, 7.092255e-13, 
    7.099316e-13, 7.108336e-13, 7.109313e-13, 7.114655e-13, 7.105899e-13, 
    7.114311e-13, 7.082468e-13, 7.096703e-13, 7.057611e-13, 7.067132e-13, 
    7.062754e-13, 7.057947e-13, 7.072777e-13, 7.088557e-13, 7.0889e-13, 
    7.093952e-13, 7.108178e-13, 7.083708e-13, 7.159404e-13, 7.11268e-13, 
    7.042725e-13, 7.057109e-13, 7.05917e-13, 7.053599e-13, 7.091383e-13, 
    7.077701e-13, 7.114526e-13, 7.104581e-13, 7.120874e-13, 7.112779e-13, 
    7.111588e-13, 7.101187e-13, 7.094706e-13, 7.078328e-13, 7.064989e-13, 
    7.054409e-13, 7.05687e-13, 7.068491e-13, 7.089523e-13, 7.109398e-13, 
    7.105045e-13, 7.119636e-13, 7.081003e-13, 7.097207e-13, 7.090946e-13, 
    7.107274e-13, 7.07148e-13, 7.101945e-13, 7.063681e-13, 7.067041e-13, 
    7.077429e-13, 7.098301e-13, 7.102927e-13, 7.107852e-13, 7.104814e-13, 
    7.090058e-13, 7.087642e-13, 7.077179e-13, 7.074286e-13, 7.06631e-13, 
    7.059701e-13, 7.065738e-13, 7.072074e-13, 7.090067e-13, 7.106258e-13, 
    7.123902e-13, 7.128219e-13, 7.148789e-13, 7.132037e-13, 7.159663e-13, 
    7.136164e-13, 7.176828e-13, 7.103719e-13, 7.135487e-13, 7.077904e-13, 
    7.084119e-13, 7.095343e-13, 7.121082e-13, 7.107198e-13, 7.123437e-13, 
    7.087547e-13, 7.068888e-13, 7.064066e-13, 7.05505e-13, 7.064272e-13, 
    7.063522e-13, 7.072341e-13, 7.069508e-13, 7.090664e-13, 7.079304e-13, 
    7.111556e-13, 7.123311e-13, 7.156472e-13, 7.176765e-13, 7.197408e-13, 
    7.20651e-13, 7.20928e-13, 7.210438e-13 ;

 LITR2C =
  1.939601e-05, 1.939599e-05, 1.939599e-05, 1.939597e-05, 1.939598e-05, 
    1.939597e-05, 1.9396e-05, 1.939598e-05, 1.939599e-05, 1.9396e-05, 
    1.939594e-05, 1.939597e-05, 1.939591e-05, 1.939593e-05, 1.939588e-05, 
    1.939591e-05, 1.939588e-05, 1.939588e-05, 1.939586e-05, 1.939587e-05, 
    1.939584e-05, 1.939586e-05, 1.939583e-05, 1.939585e-05, 1.939584e-05, 
    1.939586e-05, 1.939597e-05, 1.939595e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939598e-05, 1.939599e-05, 1.939601e-05, 1.9396e-05, 
    1.939599e-05, 1.939596e-05, 1.939597e-05, 1.939595e-05, 1.939595e-05, 
    1.939592e-05, 1.939594e-05, 1.939589e-05, 1.93959e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939588e-05, 
    1.939588e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 1.939596e-05, 
    1.939598e-05, 1.9396e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 
    1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 
    1.939593e-05, 1.939592e-05, 1.939589e-05, 1.939589e-05, 1.939589e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939586e-05, 1.939589e-05, 
    1.939587e-05, 1.93959e-05, 1.939589e-05, 1.939595e-05, 1.939597e-05, 
    1.939598e-05, 1.939599e-05, 1.939601e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 
    1.939591e-05, 1.939594e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 1.939585e-05, 
    1.939586e-05, 1.939584e-05, 1.939588e-05, 1.939587e-05, 1.939598e-05, 
    1.939598e-05, 1.939598e-05, 1.939599e-05, 1.939599e-05, 1.939601e-05, 
    1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 
    1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939588e-05, 
    1.939589e-05, 1.939588e-05, 1.939589e-05, 1.939589e-05, 1.939586e-05, 
    1.939588e-05, 1.939585e-05, 1.939585e-05, 1.939586e-05, 1.939585e-05, 
    1.939598e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 1.939601e-05, 
    1.9396e-05, 1.939599e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939588e-05, 
    1.939588e-05, 1.939588e-05, 1.939587e-05, 1.939588e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939585e-05, 1.939586e-05, 1.939585e-05, 
    1.939585e-05, 1.939598e-05, 1.939598e-05, 1.939598e-05, 1.939597e-05, 
    1.939598e-05, 1.939596e-05, 1.939595e-05, 1.939592e-05, 1.939593e-05, 
    1.939592e-05, 1.939593e-05, 1.939593e-05, 1.939592e-05, 1.939593e-05, 
    1.93959e-05, 1.939592e-05, 1.939587e-05, 1.93959e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939586e-05, 1.939585e-05, 1.939584e-05, 
    1.939584e-05, 1.939583e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939595e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939592e-05, 
    1.93959e-05, 1.93959e-05, 1.939592e-05, 1.939591e-05, 1.939595e-05, 
    1.939595e-05, 1.939595e-05, 1.939597e-05, 1.939591e-05, 1.939594e-05, 
    1.939589e-05, 1.939591e-05, 1.939586e-05, 1.939589e-05, 1.939584e-05, 
    1.939583e-05, 1.939581e-05, 1.939579e-05, 1.939595e-05, 1.939596e-05, 
    1.939595e-05, 1.939594e-05, 1.939592e-05, 1.939591e-05, 1.93959e-05, 
    1.93959e-05, 1.939589e-05, 1.939589e-05, 1.93959e-05, 1.939588e-05, 
    1.939594e-05, 1.939591e-05, 1.939596e-05, 1.939595e-05, 1.939594e-05, 
    1.939594e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939583e-05, 1.939586e-05, 1.939577e-05, 1.93958e-05, 1.939596e-05, 
    1.939595e-05, 1.939593e-05, 1.939594e-05, 1.93959e-05, 1.939589e-05, 
    1.939589e-05, 1.939588e-05, 1.939588e-05, 1.939587e-05, 1.939588e-05, 
    1.939587e-05, 1.939591e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.93959e-05, 
    1.939589e-05, 1.939588e-05, 1.93959e-05, 1.939583e-05, 1.939587e-05, 
    1.939595e-05, 1.939593e-05, 1.939593e-05, 1.939593e-05, 1.93959e-05, 
    1.939591e-05, 1.939587e-05, 1.939588e-05, 1.939587e-05, 1.939587e-05, 
    1.939588e-05, 1.939589e-05, 1.939589e-05, 1.939591e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.939588e-05, 
    1.939588e-05, 1.939587e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939588e-05, 1.939592e-05, 1.939589e-05, 1.939593e-05, 1.939592e-05, 
    1.939591e-05, 1.939589e-05, 1.939588e-05, 1.939588e-05, 1.939588e-05, 
    1.93959e-05, 1.93959e-05, 1.939591e-05, 1.939591e-05, 1.939592e-05, 
    1.939593e-05, 1.939592e-05, 1.939592e-05, 1.93959e-05, 1.939588e-05, 
    1.939586e-05, 1.939586e-05, 1.939584e-05, 1.939585e-05, 1.939583e-05, 
    1.939585e-05, 1.939581e-05, 1.939588e-05, 1.939585e-05, 1.939591e-05, 
    1.93959e-05, 1.939589e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 
    1.93959e-05, 1.939592e-05, 1.939592e-05, 1.939593e-05, 1.939592e-05, 
    1.939593e-05, 1.939592e-05, 1.939592e-05, 1.93959e-05, 1.939591e-05, 
    1.939588e-05, 1.939586e-05, 1.939583e-05, 1.939581e-05, 1.939579e-05, 
    1.939578e-05, 1.939577e-05, 1.939577e-05 ;

 LITR2C_TO_SOIL1C =
  1.063863e-13, 1.066744e-13, 1.066185e-13, 1.068506e-13, 1.067219e-13, 
    1.068739e-13, 1.064448e-13, 1.066858e-13, 1.06532e-13, 1.064123e-13, 
    1.073005e-13, 1.06861e-13, 1.077567e-13, 1.074769e-13, 1.081794e-13, 
    1.077131e-13, 1.082733e-13, 1.08166e-13, 1.084891e-13, 1.083966e-13, 
    1.088091e-13, 1.085317e-13, 1.090228e-13, 1.087429e-13, 1.087867e-13, 
    1.085226e-13, 1.069496e-13, 1.072458e-13, 1.06932e-13, 1.069743e-13, 
    1.069553e-13, 1.067245e-13, 1.066081e-13, 1.063643e-13, 1.064086e-13, 
    1.065877e-13, 1.069933e-13, 1.068557e-13, 1.072025e-13, 1.071946e-13, 
    1.075801e-13, 1.074064e-13, 1.080535e-13, 1.078698e-13, 1.084004e-13, 
    1.08267e-13, 1.083941e-13, 1.083556e-13, 1.083946e-13, 1.08199e-13, 
    1.082828e-13, 1.081106e-13, 1.074389e-13, 1.076365e-13, 1.070467e-13, 
    1.066914e-13, 1.064553e-13, 1.062877e-13, 1.063114e-13, 1.063565e-13, 
    1.065887e-13, 1.068069e-13, 1.069731e-13, 1.070841e-13, 1.071935e-13, 
    1.075242e-13, 1.076992e-13, 1.080905e-13, 1.0802e-13, 1.081395e-13, 
    1.082538e-13, 1.084453e-13, 1.084138e-13, 1.084982e-13, 1.081364e-13, 
    1.083769e-13, 1.079799e-13, 1.080885e-13, 1.072229e-13, 1.068929e-13, 
    1.067522e-13, 1.066292e-13, 1.063296e-13, 1.065365e-13, 1.06455e-13, 
    1.06649e-13, 1.067722e-13, 1.067113e-13, 1.070872e-13, 1.069411e-13, 
    1.077096e-13, 1.073788e-13, 1.082404e-13, 1.080345e-13, 1.082898e-13, 
    1.081596e-13, 1.083826e-13, 1.081819e-13, 1.085296e-13, 1.086052e-13, 
    1.085535e-13, 1.087521e-13, 1.081707e-13, 1.083941e-13, 1.067096e-13, 
    1.067195e-13, 1.067658e-13, 1.065622e-13, 1.065498e-13, 1.063631e-13, 
    1.065292e-13, 1.065999e-13, 1.067794e-13, 1.068854e-13, 1.069862e-13, 
    1.072077e-13, 1.074548e-13, 1.078001e-13, 1.080479e-13, 1.082138e-13, 
    1.081121e-13, 1.082019e-13, 1.081015e-13, 1.080544e-13, 1.085768e-13, 
    1.082836e-13, 1.087235e-13, 1.086992e-13, 1.085002e-13, 1.08702e-13, 
    1.067265e-13, 1.066693e-13, 1.064706e-13, 1.066261e-13, 1.063428e-13, 
    1.065014e-13, 1.065925e-13, 1.069441e-13, 1.070213e-13, 1.070928e-13, 
    1.072341e-13, 1.074153e-13, 1.077327e-13, 1.080087e-13, 1.082604e-13, 
    1.08242e-13, 1.082485e-13, 1.083047e-13, 1.081654e-13, 1.083275e-13, 
    1.083547e-13, 1.082836e-13, 1.08696e-13, 1.085782e-13, 1.086987e-13, 
    1.086221e-13, 1.066879e-13, 1.067841e-13, 1.067321e-13, 1.068299e-13, 
    1.06761e-13, 1.07067e-13, 1.071587e-13, 1.075875e-13, 1.074117e-13, 
    1.076915e-13, 1.074401e-13, 1.074847e-13, 1.077005e-13, 1.074538e-13, 
    1.079935e-13, 1.076276e-13, 1.083068e-13, 1.079418e-13, 1.083297e-13, 
    1.082593e-13, 1.083759e-13, 1.084801e-13, 1.086113e-13, 1.088531e-13, 
    1.087971e-13, 1.089993e-13, 1.069275e-13, 1.070522e-13, 1.070413e-13, 
    1.071717e-13, 1.072681e-13, 1.07477e-13, 1.078117e-13, 1.076859e-13, 
    1.079168e-13, 1.079632e-13, 1.076123e-13, 1.078277e-13, 1.071356e-13, 
    1.072475e-13, 1.071809e-13, 1.069373e-13, 1.077148e-13, 1.07316e-13, 
    1.080519e-13, 1.078363e-13, 1.084653e-13, 1.081526e-13, 1.087663e-13, 
    1.090281e-13, 1.092745e-13, 1.095619e-13, 1.071202e-13, 1.070356e-13, 
    1.071872e-13, 1.073968e-13, 1.075912e-13, 1.078495e-13, 1.078759e-13, 
    1.079242e-13, 1.080494e-13, 1.081546e-13, 1.079395e-13, 1.08181e-13, 
    1.072733e-13, 1.077494e-13, 1.070035e-13, 1.072282e-13, 1.073845e-13, 
    1.07316e-13, 1.076715e-13, 1.077552e-13, 1.080951e-13, 1.079195e-13, 
    1.089634e-13, 1.085021e-13, 1.097807e-13, 1.094239e-13, 1.07006e-13, 
    1.0712e-13, 1.075163e-13, 1.073278e-13, 1.078667e-13, 1.079992e-13, 
    1.081068e-13, 1.082443e-13, 1.082592e-13, 1.083407e-13, 1.082072e-13, 
    1.083354e-13, 1.0785e-13, 1.08067e-13, 1.074711e-13, 1.076163e-13, 
    1.075495e-13, 1.074763e-13, 1.077023e-13, 1.079428e-13, 1.079481e-13, 
    1.080251e-13, 1.082419e-13, 1.078689e-13, 1.090227e-13, 1.083105e-13, 
    1.072443e-13, 1.074635e-13, 1.074949e-13, 1.0741e-13, 1.079859e-13, 
    1.077774e-13, 1.083387e-13, 1.081871e-13, 1.084354e-13, 1.083121e-13, 
    1.082939e-13, 1.081353e-13, 1.080366e-13, 1.077869e-13, 1.075836e-13, 
    1.074223e-13, 1.074598e-13, 1.07637e-13, 1.079576e-13, 1.082605e-13, 
    1.081942e-13, 1.084166e-13, 1.078277e-13, 1.080747e-13, 1.079793e-13, 
    1.082281e-13, 1.076825e-13, 1.081469e-13, 1.075637e-13, 1.076149e-13, 
    1.077732e-13, 1.080914e-13, 1.081619e-13, 1.082369e-13, 1.081907e-13, 
    1.079657e-13, 1.079289e-13, 1.077694e-13, 1.077253e-13, 1.076037e-13, 
    1.07503e-13, 1.07595e-13, 1.076916e-13, 1.079659e-13, 1.082127e-13, 
    1.084816e-13, 1.085474e-13, 1.088609e-13, 1.086056e-13, 1.090267e-13, 
    1.086685e-13, 1.092883e-13, 1.081739e-13, 1.086582e-13, 1.077805e-13, 
    1.078752e-13, 1.080463e-13, 1.084386e-13, 1.08227e-13, 1.084745e-13, 
    1.079275e-13, 1.07643e-13, 1.075695e-13, 1.074321e-13, 1.075727e-13, 
    1.075612e-13, 1.076957e-13, 1.076525e-13, 1.07975e-13, 1.078018e-13, 
    1.082934e-13, 1.084726e-13, 1.089781e-13, 1.092874e-13, 1.096021e-13, 
    1.097408e-13, 1.09783e-13, 1.098007e-13 ;

 LITR2C_vr =
  0.001107532, 0.001107531, 0.001107531, 0.00110753, 0.001107531, 0.00110753, 
    0.001107532, 0.001107531, 0.001107531, 0.001107532, 0.001107528, 
    0.00110753, 0.001107527, 0.001107528, 0.001107525, 0.001107527, 
    0.001107525, 0.001107525, 0.001107524, 0.001107524, 0.001107523, 
    0.001107524, 0.001107522, 0.001107523, 0.001107523, 0.001107524, 
    0.00110753, 0.001107529, 0.00110753, 0.00110753, 0.00110753, 0.001107531, 
    0.001107531, 0.001107532, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.001107527, 0.001107528, 
    0.001107525, 0.001107526, 0.001107524, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107525, 0.001107525, 
    0.001107528, 0.001107527, 0.001107529, 0.001107531, 0.001107532, 
    0.001107532, 0.001107532, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107527, 
    0.001107525, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107529, 0.00110753, 0.001107531, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.00110753, 
    0.001107531, 0.001107529, 0.00110753, 0.001107527, 0.001107528, 
    0.001107525, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107525, 0.001107524, 0.001107523, 0.001107524, 0.001107523, 
    0.001107525, 0.001107524, 0.001107531, 0.001107531, 0.00110753, 
    0.001107531, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.00110753, 0.00110753, 0.00110753, 0.001107529, 0.001107528, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107525, 
    0.001107525, 0.001107525, 0.001107523, 0.001107525, 0.001107523, 
    0.001107523, 0.001107524, 0.001107523, 0.001107531, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.00110753, 0.00110753, 0.001107529, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107525, 0.001107525, 
    0.001107524, 0.001107525, 0.001107524, 0.001107524, 0.001107525, 
    0.001107523, 0.001107523, 0.001107523, 0.001107523, 0.001107531, 
    0.00110753, 0.001107531, 0.00110753, 0.00110753, 0.001107529, 
    0.001107529, 0.001107527, 0.001107528, 0.001107527, 0.001107528, 
    0.001107528, 0.001107527, 0.001107528, 0.001107526, 0.001107527, 
    0.001107524, 0.001107526, 0.001107524, 0.001107525, 0.001107524, 
    0.001107524, 0.001107523, 0.001107522, 0.001107523, 0.001107522, 
    0.00110753, 0.001107529, 0.001107529, 0.001107529, 0.001107529, 
    0.001107528, 0.001107526, 0.001107527, 0.001107526, 0.001107526, 
    0.001107527, 0.001107526, 0.001107529, 0.001107529, 0.001107529, 
    0.00110753, 0.001107527, 0.001107528, 0.001107526, 0.001107526, 
    0.001107524, 0.001107525, 0.001107523, 0.001107522, 0.001107521, 
    0.00110752, 0.001107529, 0.001107529, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107526, 
    0.001107525, 0.001107526, 0.001107525, 0.001107528, 0.001107527, 
    0.00110753, 0.001107529, 0.001107528, 0.001107528, 0.001107527, 
    0.001107527, 0.001107525, 0.001107526, 0.001107522, 0.001107524, 
    0.001107519, 0.00110752, 0.00110753, 0.001107529, 0.001107528, 
    0.001107528, 0.001107526, 0.001107526, 0.001107525, 0.001107525, 
    0.001107525, 0.001107524, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107528, 0.001107527, 0.001107527, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107526, 0.001107522, 0.001107524, 0.001107529, 0.001107528, 
    0.001107528, 0.001107528, 0.001107526, 0.001107527, 0.001107524, 
    0.001107525, 0.001107524, 0.001107524, 0.001107524, 0.001107525, 
    0.001107526, 0.001107526, 0.001107527, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107526, 0.001107525, 0.001107526, 0.001107525, 0.001107527, 
    0.001107525, 0.001107527, 0.001107527, 0.001107527, 0.001107525, 
    0.001107525, 0.001107525, 0.001107525, 0.001107526, 0.001107526, 
    0.001107527, 0.001107527, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107526, 0.001107525, 0.001107524, 0.001107524, 
    0.001107522, 0.001107523, 0.001107522, 0.001107523, 0.001107521, 
    0.001107525, 0.001107523, 0.001107527, 0.001107526, 0.001107526, 
    0.001107524, 0.001107525, 0.001107524, 0.001107526, 0.001107527, 
    0.001107527, 0.001107528, 0.001107527, 0.001107527, 0.001107527, 
    0.001107527, 0.001107526, 0.001107526, 0.001107524, 0.001107524, 
    0.001107522, 0.001107521, 0.001107519, 0.001107519, 0.001107519, 
    0.001107519,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684264e-07, 2.684262e-07, 2.684262e-07, 2.68426e-07, 2.684261e-07, 
    2.68426e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 2.684264e-07, 
    2.684256e-07, 2.68426e-07, 2.684252e-07, 2.684254e-07, 2.684248e-07, 
    2.684252e-07, 2.684247e-07, 2.684248e-07, 2.684245e-07, 2.684246e-07, 
    2.684242e-07, 2.684244e-07, 2.68424e-07, 2.684242e-07, 2.684242e-07, 
    2.684244e-07, 2.684259e-07, 2.684257e-07, 2.684259e-07, 2.684259e-07, 
    2.684259e-07, 2.684261e-07, 2.684262e-07, 2.684265e-07, 2.684264e-07, 
    2.684262e-07, 2.684259e-07, 2.68426e-07, 2.684257e-07, 2.684257e-07, 
    2.684253e-07, 2.684255e-07, 2.684249e-07, 2.684251e-07, 2.684245e-07, 
    2.684247e-07, 2.684246e-07, 2.684246e-07, 2.684246e-07, 2.684247e-07, 
    2.684247e-07, 2.684248e-07, 2.684255e-07, 2.684253e-07, 2.684258e-07, 
    2.684262e-07, 2.684264e-07, 2.684265e-07, 2.684265e-07, 2.684265e-07, 
    2.684262e-07, 2.68426e-07, 2.684259e-07, 2.684258e-07, 2.684257e-07, 
    2.684254e-07, 2.684252e-07, 2.684249e-07, 2.684249e-07, 2.684248e-07, 
    2.684247e-07, 2.684245e-07, 2.684245e-07, 2.684245e-07, 2.684248e-07, 
    2.684246e-07, 2.684249e-07, 2.684249e-07, 2.684257e-07, 2.68426e-07, 
    2.684261e-07, 2.684262e-07, 2.684265e-07, 2.684263e-07, 2.684264e-07, 
    2.684262e-07, 2.684261e-07, 2.684261e-07, 2.684258e-07, 2.684259e-07, 
    2.684252e-07, 2.684255e-07, 2.684247e-07, 2.684249e-07, 2.684247e-07, 
    2.684248e-07, 2.684246e-07, 2.684248e-07, 2.684244e-07, 2.684244e-07, 
    2.684244e-07, 2.684242e-07, 2.684248e-07, 2.684246e-07, 2.684261e-07, 
    2.684261e-07, 2.684261e-07, 2.684263e-07, 2.684263e-07, 2.684265e-07, 
    2.684263e-07, 2.684262e-07, 2.684261e-07, 2.68426e-07, 2.684259e-07, 
    2.684257e-07, 2.684255e-07, 2.684251e-07, 2.684249e-07, 2.684247e-07, 
    2.684248e-07, 2.684247e-07, 2.684248e-07, 2.684249e-07, 2.684244e-07, 
    2.684247e-07, 2.684243e-07, 2.684243e-07, 2.684245e-07, 2.684243e-07, 
    2.684261e-07, 2.684262e-07, 2.684264e-07, 2.684262e-07, 2.684265e-07, 
    2.684263e-07, 2.684262e-07, 2.684259e-07, 2.684259e-07, 2.684258e-07, 
    2.684257e-07, 2.684255e-07, 2.684252e-07, 2.684249e-07, 2.684247e-07, 
    2.684247e-07, 2.684247e-07, 2.684247e-07, 2.684248e-07, 2.684246e-07, 
    2.684246e-07, 2.684247e-07, 2.684243e-07, 2.684244e-07, 2.684243e-07, 
    2.684243e-07, 2.684262e-07, 2.684261e-07, 2.684261e-07, 2.68426e-07, 
    2.684261e-07, 2.684258e-07, 2.684257e-07, 2.684253e-07, 2.684255e-07, 
    2.684252e-07, 2.684255e-07, 2.684254e-07, 2.684252e-07, 2.684255e-07, 
    2.684249e-07, 2.684253e-07, 2.684247e-07, 2.68425e-07, 2.684246e-07, 
    2.684247e-07, 2.684246e-07, 2.684245e-07, 2.684244e-07, 2.684241e-07, 
    2.684242e-07, 2.68424e-07, 2.684259e-07, 2.684258e-07, 2.684258e-07, 
    2.684257e-07, 2.684256e-07, 2.684254e-07, 2.684251e-07, 2.684252e-07, 
    2.68425e-07, 2.68425e-07, 2.684253e-07, 2.684251e-07, 2.684257e-07, 
    2.684257e-07, 2.684257e-07, 2.684259e-07, 2.684252e-07, 2.684256e-07, 
    2.684249e-07, 2.684251e-07, 2.684245e-07, 2.684248e-07, 2.684242e-07, 
    2.68424e-07, 2.684237e-07, 2.684235e-07, 2.684258e-07, 2.684259e-07, 
    2.684257e-07, 2.684255e-07, 2.684253e-07, 2.684251e-07, 2.684251e-07, 
    2.68425e-07, 2.684249e-07, 2.684248e-07, 2.68425e-07, 2.684248e-07, 
    2.684256e-07, 2.684252e-07, 2.684259e-07, 2.684257e-07, 2.684255e-07, 
    2.684256e-07, 2.684253e-07, 2.684252e-07, 2.684249e-07, 2.68425e-07, 
    2.68424e-07, 2.684245e-07, 2.684233e-07, 2.684236e-07, 2.684259e-07, 
    2.684258e-07, 2.684254e-07, 2.684256e-07, 2.684251e-07, 2.684249e-07, 
    2.684248e-07, 2.684247e-07, 2.684247e-07, 2.684246e-07, 2.684247e-07, 
    2.684246e-07, 2.684251e-07, 2.684249e-07, 2.684254e-07, 2.684253e-07, 
    2.684254e-07, 2.684254e-07, 2.684252e-07, 2.68425e-07, 2.68425e-07, 
    2.684249e-07, 2.684247e-07, 2.684251e-07, 2.68424e-07, 2.684246e-07, 
    2.684257e-07, 2.684254e-07, 2.684254e-07, 2.684255e-07, 2.684249e-07, 
    2.684251e-07, 2.684246e-07, 2.684248e-07, 2.684245e-07, 2.684246e-07, 
    2.684247e-07, 2.684248e-07, 2.684249e-07, 2.684251e-07, 2.684253e-07, 
    2.684255e-07, 2.684255e-07, 2.684253e-07, 2.68425e-07, 2.684247e-07, 
    2.684247e-07, 2.684245e-07, 2.684251e-07, 2.684249e-07, 2.684249e-07, 
    2.684247e-07, 2.684252e-07, 2.684248e-07, 2.684253e-07, 2.684253e-07, 
    2.684251e-07, 2.684249e-07, 2.684248e-07, 2.684247e-07, 2.684247e-07, 
    2.68425e-07, 2.68425e-07, 2.684251e-07, 2.684252e-07, 2.684253e-07, 
    2.684254e-07, 2.684253e-07, 2.684252e-07, 2.68425e-07, 2.684247e-07, 
    2.684245e-07, 2.684244e-07, 2.684241e-07, 2.684244e-07, 2.68424e-07, 
    2.684243e-07, 2.684237e-07, 2.684248e-07, 2.684243e-07, 2.684251e-07, 
    2.684251e-07, 2.684249e-07, 2.684245e-07, 2.684247e-07, 2.684245e-07, 
    2.68425e-07, 2.684253e-07, 2.684253e-07, 2.684255e-07, 2.684253e-07, 
    2.684253e-07, 2.684252e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684247e-07, 2.684245e-07, 2.68424e-07, 2.684237e-07, 2.684234e-07, 
    2.684233e-07, 2.684233e-07, 2.684232e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  1.642107e-25, 7.597807e-26, -1.715634e-25, -4.901811e-26, -2.205815e-26, 
    -1.02938e-25, -7.352717e-26, -1.176435e-25, -4.901811e-26, -1.56858e-25, 
    -9.803622e-27, 1.323489e-25, 7.352717e-27, -6.617445e-26, -2.769523e-25, 
    1.715634e-26, 2.450905e-26, 1.053889e-25, -2.132288e-25, 5.882173e-26, 
    -1.960724e-26, -1.960724e-26, 4.901811e-26, -1.053889e-25, 2.671487e-25, 
    -5.637083e-26, 1.54407e-25, -1.715634e-26, 9.068351e-26, -1.470543e-26, 
    -2.205815e-26, -2.941087e-26, -7.107626e-26, -5.146902e-26, 
    -1.666616e-25, -2.303851e-25, 2.205815e-26, -1.176435e-25, -1.102908e-25, 
    -2.156797e-25, -1.936215e-25, 9.313441e-26, 3.921449e-26, 2.941087e-26, 
    -5.637083e-26, -1.02938e-25, 4.901811e-27, -1.54407e-25, 6.617445e-26, 
    1.446034e-25, 5.882173e-26, -1.715634e-26, 1.29898e-25, -1.960724e-25, 
    2.230324e-25, -8.333079e-26, -1.347998e-25, -7.842898e-26, 6.372354e-26, 
    1.200944e-25, 4.901811e-26, 5.637083e-26, -7.107626e-26, 4.65672e-26, 
    1.078398e-25, -1.176435e-25, -2.230324e-25, 1.715634e-26, 6.862535e-26, 
    7.352717e-27, -1.347998e-25, 6.862535e-26, -8.333079e-26, 4.41163e-26, 
    -2.450905e-26, 3.186177e-26, -8.578169e-26, -1.421525e-25, 2.450905e-26, 
    -1.225453e-25, -8.333079e-26, -2.450905e-26, -1.470543e-25, 
    -1.151926e-25, 1.960724e-26, 1.740143e-25, -7.107626e-26, 7.597807e-26, 
    -1.887197e-25, -4.41163e-26, -3.921449e-26, -4.901811e-27, 1.54407e-25, 
    -1.372507e-25, 3.357741e-25, -1.715634e-26, 4.65672e-26, 1.323489e-25, 
    2.59796e-25, -1.078398e-25, 1.225453e-26, -2.450905e-26, -1.862688e-25, 
    -1.200944e-25, 3.676358e-26, 1.960724e-26, 6.617445e-26, 0, 9.803622e-26, 
    -1.176435e-25, 3.921449e-26, -1.249962e-25, -1.127417e-25, -5.882173e-26, 
    9.313441e-26, 6.617445e-26, 2.59796e-25, 7.352717e-27, -7.352717e-27, 
    -1.470543e-26, -9.803622e-26, -1.715634e-26, -4.65672e-26, -8.333079e-26, 
    1.225453e-25, 2.401887e-25, -2.32836e-25, -4.901811e-27, -2.08327e-25, 
    -9.803622e-27, 2.450906e-27, 1.838179e-25, 9.558531e-26, 1.127417e-25, 
    9.558531e-26, -1.691125e-25, 7.352717e-26, -4.901811e-26, -9.068351e-26, 
    -1.176435e-25, -6.127264e-26, 1.446034e-25, 3.676358e-26, -1.960724e-26, 
    5.882173e-26, -1.078398e-25, 5.391992e-26, 2.181306e-25, -2.450906e-27, 
    1.225453e-26, 8.333079e-26, -1.397016e-25, -1.666616e-25, 3.186177e-26, 
    6.372354e-26, 4.41163e-26, -7.842898e-26, 5.391992e-26, 1.838179e-25, 
    -1.372507e-25, -4.142031e-25, -7.352717e-27, -1.02938e-25, 1.225453e-25, 
    1.397016e-25, -1.887197e-25, -9.068351e-26, -4.166539e-26, -1.960724e-26, 
    6.127264e-26, 6.617445e-26, -9.313441e-26, -1.715634e-26, 5.391992e-26, 
    -3.749886e-25, 1.372507e-25, 1.372507e-25, -8.333079e-26, -1.02938e-25, 
    1.642107e-25, -1.347998e-25, -4.901811e-26, -1.960724e-25, 3.921449e-26, 
    2.450905e-26, 4.901811e-27, 1.053889e-25, -1.617598e-25, -7.352717e-27, 
    4.166539e-26, 8.333079e-26, -1.200944e-25, -1.936215e-25, 1.176435e-25, 
    -1.691125e-25, 7.597807e-26, -2.32836e-25, 1.470543e-26, -2.450905e-26, 
    3.186177e-26, 1.397016e-25, -2.132288e-25, -1.397016e-25, 1.372507e-25, 
    1.519561e-25, -2.32836e-25, -1.053889e-25, 1.397016e-25, -5.146902e-26, 
    -1.372507e-25, 1.715634e-25, 1.789161e-25, -6.372354e-26, 2.034252e-25, 
    -4.166539e-26, 2.941087e-26, 2.450905e-26, 1.56858e-25, 7.842898e-26, 
    -4.901811e-27, 1.887197e-25, -8.333079e-26, -7.107626e-26, -4.901811e-27, 
    -5.882173e-26, 1.470543e-26, -9.803622e-27, 1.838179e-25, 2.205815e-26, 
    -5.146902e-26, -1.617598e-25, -5.637083e-26, -7.597807e-26, -8.82326e-26, 
    7.842898e-26, -2.377378e-25, 1.446034e-25, 1.789161e-25, 1.715634e-25, 
    1.519561e-25, 2.450906e-27, -5.391992e-26, -1.053889e-25, -1.54407e-25, 
    -7.352717e-26, -1.372507e-25, 5.391992e-26, 6.372354e-26, -5.637083e-26, 
    3.186177e-26, 1.225453e-25, -2.941087e-25, -1.274471e-25, 1.54407e-25, 
    -6.127264e-26, -1.078398e-25, -2.941087e-25, 1.29898e-25, -1.911706e-25, 
    7.597807e-26, 3.431268e-26, -7.107626e-26, 4.591775e-41, 1.56858e-25, 
    -1.004871e-25, -1.519561e-25, 1.81367e-25, 2.401887e-25, -8.82326e-26, 
    1.225453e-26, -1.102908e-25, 1.56858e-25, -1.004871e-25, 6.617445e-26, 
    -2.352869e-25, 1.200944e-25, -2.205815e-26, -1.691125e-25, 4.41163e-26, 
    -3.676358e-26, 5.882173e-26, 1.397016e-25, -1.225453e-25, -1.56858e-25, 
    -8.087988e-26, -3.088141e-25, -4.901811e-26, -5.882173e-26, 
    -6.372354e-26, -1.225453e-25, 1.960724e-26, 1.446034e-25, 1.470543e-26, 
    2.352869e-25, -1.446034e-25, -7.597807e-26, 9.803622e-27, 4.65672e-26, 
    -1.764652e-25, 8.333079e-26, -8.087988e-26, -3.921449e-26, -6.127264e-26, 
    -1.176435e-25, 1.176435e-25, -3.210686e-25, 9.313441e-26, -4.65672e-26, 
    1.397016e-25, -8.333079e-26, 5.882173e-26, -1.200944e-25, 7.107626e-26, 
    -2.450905e-26, 1.225453e-25, 5.882173e-26, -6.862535e-26, -1.053889e-25, 
    -2.450906e-27, -1.225453e-26, 1.397016e-25, 3.210686e-25, 1.053889e-25, 
    5.391992e-26, -1.225453e-26, -1.862688e-25, -4.166539e-26, -1.960724e-26, 
    8.087988e-26, -5.882173e-26, 7.107626e-26, 2.475414e-25, 1.225453e-25, 
    -2.205815e-26, -1.764652e-25, 1.495052e-25, 1.887197e-25, 7.352717e-26,
  2.676251e-32, 2.676248e-32, 2.676249e-32, 2.676246e-32, 2.676247e-32, 
    2.676246e-32, 2.67625e-32, 2.676248e-32, 2.676249e-32, 2.67625e-32, 
    2.676242e-32, 2.676246e-32, 2.676238e-32, 2.67624e-32, 2.676234e-32, 
    2.676238e-32, 2.676233e-32, 2.676234e-32, 2.676231e-32, 2.676232e-32, 
    2.676228e-32, 2.67623e-32, 2.676226e-32, 2.676229e-32, 2.676228e-32, 
    2.676231e-32, 2.676245e-32, 2.676243e-32, 2.676246e-32, 2.676245e-32, 
    2.676245e-32, 2.676247e-32, 2.676249e-32, 2.676251e-32, 2.676251e-32, 
    2.676249e-32, 2.676245e-32, 2.676246e-32, 2.676243e-32, 2.676243e-32, 
    2.676239e-32, 2.676241e-32, 2.676235e-32, 2.676237e-32, 2.676232e-32, 
    2.676233e-32, 2.676232e-32, 2.676232e-32, 2.676232e-32, 2.676234e-32, 
    2.676233e-32, 2.676234e-32, 2.676241e-32, 2.676239e-32, 2.676244e-32, 
    2.676248e-32, 2.67625e-32, 2.676252e-32, 2.676252e-32, 2.676251e-32, 
    2.676249e-32, 2.676247e-32, 2.676245e-32, 2.676244e-32, 2.676243e-32, 
    2.67624e-32, 2.676238e-32, 2.676235e-32, 2.676235e-32, 2.676234e-32, 
    2.676233e-32, 2.676231e-32, 2.676232e-32, 2.676231e-32, 2.676234e-32, 
    2.676232e-32, 2.676236e-32, 2.676235e-32, 2.676243e-32, 2.676246e-32, 
    2.676247e-32, 2.676248e-32, 2.676251e-32, 2.676249e-32, 2.67625e-32, 
    2.676248e-32, 2.676247e-32, 2.676248e-32, 2.676244e-32, 2.676245e-32, 
    2.676238e-32, 2.676241e-32, 2.676233e-32, 2.676235e-32, 2.676233e-32, 
    2.676234e-32, 2.676232e-32, 2.676234e-32, 2.67623e-32, 2.67623e-32, 
    2.67623e-32, 2.676228e-32, 2.676234e-32, 2.676232e-32, 2.676248e-32, 
    2.676248e-32, 2.676247e-32, 2.676249e-32, 2.676249e-32, 2.676251e-32, 
    2.676249e-32, 2.676249e-32, 2.676247e-32, 2.676246e-32, 2.676245e-32, 
    2.676243e-32, 2.676241e-32, 2.676237e-32, 2.676235e-32, 2.676234e-32, 
    2.676234e-32, 2.676234e-32, 2.676234e-32, 2.676235e-32, 2.67623e-32, 
    2.676233e-32, 2.676229e-32, 2.676229e-32, 2.676231e-32, 2.676229e-32, 
    2.676247e-32, 2.676248e-32, 2.67625e-32, 2.676249e-32, 2.676251e-32, 
    2.67625e-32, 2.676249e-32, 2.676245e-32, 2.676245e-32, 2.676244e-32, 
    2.676243e-32, 2.676241e-32, 2.676238e-32, 2.676235e-32, 2.676233e-32, 
    2.676233e-32, 2.676233e-32, 2.676233e-32, 2.676234e-32, 2.676232e-32, 
    2.676232e-32, 2.676233e-32, 2.676229e-32, 2.67623e-32, 2.676229e-32, 
    2.676229e-32, 2.676248e-32, 2.676247e-32, 2.676247e-32, 2.676247e-32, 
    2.676247e-32, 2.676244e-32, 2.676243e-32, 2.676239e-32, 2.676241e-32, 
    2.676238e-32, 2.676241e-32, 2.67624e-32, 2.676238e-32, 2.676241e-32, 
    2.676236e-32, 2.676239e-32, 2.676233e-32, 2.676236e-32, 2.676232e-32, 
    2.676233e-32, 2.676232e-32, 2.676231e-32, 2.67623e-32, 2.676227e-32, 
    2.676228e-32, 2.676226e-32, 2.676246e-32, 2.676244e-32, 2.676244e-32, 
    2.676243e-32, 2.676242e-32, 2.67624e-32, 2.676237e-32, 2.676239e-32, 
    2.676236e-32, 2.676236e-32, 2.676239e-32, 2.676237e-32, 2.676244e-32, 
    2.676243e-32, 2.676243e-32, 2.676246e-32, 2.676238e-32, 2.676242e-32, 
    2.676235e-32, 2.676237e-32, 2.676231e-32, 2.676234e-32, 2.676228e-32, 
    2.676226e-32, 2.676224e-32, 2.676221e-32, 2.676244e-32, 2.676244e-32, 
    2.676243e-32, 2.676241e-32, 2.676239e-32, 2.676237e-32, 2.676237e-32, 
    2.676236e-32, 2.676235e-32, 2.676234e-32, 2.676236e-32, 2.676234e-32, 
    2.676242e-32, 2.676238e-32, 2.676245e-32, 2.676243e-32, 2.676241e-32, 
    2.676242e-32, 2.676239e-32, 2.676238e-32, 2.676234e-32, 2.676236e-32, 
    2.676227e-32, 2.676231e-32, 2.676219e-32, 2.676222e-32, 2.676245e-32, 
    2.676244e-32, 2.67624e-32, 2.676242e-32, 2.676237e-32, 2.676235e-32, 
    2.676234e-32, 2.676233e-32, 2.676233e-32, 2.676232e-32, 2.676234e-32, 
    2.676232e-32, 2.676237e-32, 2.676235e-32, 2.67624e-32, 2.676239e-32, 
    2.67624e-32, 2.67624e-32, 2.676238e-32, 2.676236e-32, 2.676236e-32, 
    2.676235e-32, 2.676233e-32, 2.676237e-32, 2.676226e-32, 2.676232e-32, 
    2.676243e-32, 2.676241e-32, 2.67624e-32, 2.676241e-32, 2.676236e-32, 
    2.676238e-32, 2.676232e-32, 2.676234e-32, 2.676231e-32, 2.676232e-32, 
    2.676233e-32, 2.676234e-32, 2.676235e-32, 2.676237e-32, 2.676239e-32, 
    2.676241e-32, 2.676241e-32, 2.676239e-32, 2.676236e-32, 2.676233e-32, 
    2.676234e-32, 2.676232e-32, 2.676237e-32, 2.676235e-32, 2.676236e-32, 
    2.676233e-32, 2.676239e-32, 2.676234e-32, 2.676239e-32, 2.676239e-32, 
    2.676238e-32, 2.676234e-32, 2.676234e-32, 2.676233e-32, 2.676234e-32, 
    2.676236e-32, 2.676236e-32, 2.676238e-32, 2.676238e-32, 2.676239e-32, 
    2.67624e-32, 2.676239e-32, 2.676238e-32, 2.676236e-32, 2.676234e-32, 
    2.676231e-32, 2.67623e-32, 2.676227e-32, 2.67623e-32, 2.676226e-32, 
    2.676229e-32, 2.676223e-32, 2.676234e-32, 2.676229e-32, 2.676237e-32, 
    2.676237e-32, 2.676235e-32, 2.676231e-32, 2.676233e-32, 2.676231e-32, 
    2.676236e-32, 2.676239e-32, 2.676239e-32, 2.676241e-32, 2.676239e-32, 
    2.67624e-32, 2.676238e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676233e-32, 2.676231e-32, 2.676226e-32, 2.676223e-32, 2.67622e-32, 
    2.676219e-32, 2.676219e-32, 2.676219e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  2.944617e-15, 2.952591e-15, 2.951042e-15, 2.957468e-15, 2.953905e-15, 
    2.958111e-15, 2.946235e-15, 2.952907e-15, 2.948649e-15, 2.945336e-15, 
    2.969921e-15, 2.957755e-15, 2.982548e-15, 2.974803e-15, 2.994246e-15, 
    2.981342e-15, 2.996847e-15, 2.993877e-15, 3.002818e-15, 3.000258e-15, 
    3.011675e-15, 3.003999e-15, 3.017592e-15, 3.009844e-15, 3.011056e-15, 
    3.003745e-15, 2.960208e-15, 2.968406e-15, 2.959721e-15, 2.960891e-15, 
    2.960367e-15, 2.953978e-15, 2.950755e-15, 2.944009e-15, 2.945234e-15, 
    2.95019e-15, 2.961417e-15, 2.95761e-15, 2.967207e-15, 2.96699e-15, 
    2.977659e-15, 2.972851e-15, 2.990761e-15, 2.985676e-15, 3.000365e-15, 
    2.996673e-15, 3.000191e-15, 2.999124e-15, 3.000204e-15, 2.994789e-15, 
    2.99711e-15, 2.992344e-15, 2.973751e-15, 2.97922e-15, 2.962896e-15, 
    2.953061e-15, 2.946528e-15, 2.941886e-15, 2.942543e-15, 2.943793e-15, 
    2.950219e-15, 2.956258e-15, 2.960857e-15, 2.963931e-15, 2.966959e-15, 
    2.976111e-15, 2.980956e-15, 2.991787e-15, 2.989836e-15, 2.993143e-15, 
    2.996305e-15, 3.001608e-15, 3.000735e-15, 3.00307e-15, 2.993058e-15, 
    2.999713e-15, 2.988725e-15, 2.99173e-15, 2.967773e-15, 2.958637e-15, 
    2.954743e-15, 2.95134e-15, 2.943047e-15, 2.948774e-15, 2.946517e-15, 
    2.951888e-15, 2.955298e-15, 2.953612e-15, 2.964015e-15, 2.959972e-15, 
    2.981243e-15, 2.972088e-15, 2.995936e-15, 2.990237e-15, 2.997303e-15, 
    2.993698e-15, 2.999872e-15, 2.994316e-15, 3.003939e-15, 3.006032e-15, 
    3.004602e-15, 3.010098e-15, 2.994008e-15, 3.00019e-15, 2.953565e-15, 
    2.95384e-15, 2.955121e-15, 2.949485e-15, 2.949141e-15, 2.943975e-15, 
    2.948572e-15, 2.950529e-15, 2.955497e-15, 2.958432e-15, 2.961222e-15, 
    2.967353e-15, 2.974192e-15, 2.983748e-15, 2.990606e-15, 2.9952e-15, 
    2.992384e-15, 2.99487e-15, 2.992091e-15, 2.990788e-15, 3.005247e-15, 
    2.997131e-15, 3.009308e-15, 3.008635e-15, 3.003125e-15, 3.00871e-15, 
    2.954033e-15, 2.95245e-15, 2.94695e-15, 2.951255e-15, 2.943412e-15, 
    2.947802e-15, 2.950324e-15, 2.960054e-15, 2.962193e-15, 2.964173e-15, 
    2.968083e-15, 2.973097e-15, 2.981884e-15, 2.989521e-15, 2.99649e-15, 
    2.995979e-15, 2.996159e-15, 2.997714e-15, 2.99386e-15, 2.998346e-15, 
    2.999098e-15, 2.997131e-15, 3.008544e-15, 3.005286e-15, 3.00862e-15, 
    3.006499e-15, 2.952965e-15, 2.955628e-15, 2.954189e-15, 2.956894e-15, 
    2.954988e-15, 2.963458e-15, 2.965996e-15, 2.977863e-15, 2.972998e-15, 
    2.980742e-15, 2.973786e-15, 2.975018e-15, 2.980991e-15, 2.974162e-15, 
    2.9891e-15, 2.978972e-15, 2.997774e-15, 2.98767e-15, 2.998407e-15, 
    2.996459e-15, 2.999684e-15, 3.00257e-15, 3.006201e-15, 3.012894e-15, 
    3.011345e-15, 3.01694e-15, 2.959597e-15, 2.963047e-15, 2.962745e-15, 
    2.966355e-15, 2.969023e-15, 2.974806e-15, 2.984069e-15, 2.980588e-15, 
    2.98698e-15, 2.988262e-15, 2.978551e-15, 2.984513e-15, 2.965356e-15, 
    2.968453e-15, 2.966611e-15, 2.959868e-15, 2.981388e-15, 2.97035e-15, 
    2.990719e-15, 2.984751e-15, 3.002159e-15, 2.993504e-15, 3.010492e-15, 
    3.017737e-15, 3.024558e-15, 3.032512e-15, 2.964931e-15, 2.962587e-15, 
    2.966785e-15, 2.972585e-15, 2.977968e-15, 2.985115e-15, 2.985847e-15, 
    2.987185e-15, 2.990649e-15, 2.993561e-15, 2.987606e-15, 2.994291e-15, 
    2.969167e-15, 2.982346e-15, 2.961699e-15, 2.96792e-15, 2.972244e-15, 
    2.970349e-15, 2.98019e-15, 2.982507e-15, 2.991912e-15, 2.987054e-15, 
    3.015948e-15, 3.003177e-15, 3.038567e-15, 3.028694e-15, 2.961768e-15, 
    2.964924e-15, 2.975894e-15, 2.970677e-15, 2.985593e-15, 2.989259e-15, 
    2.992238e-15, 2.996044e-15, 2.996456e-15, 2.99871e-15, 2.995016e-15, 
    2.998565e-15, 2.98513e-15, 2.991136e-15, 2.974643e-15, 2.97866e-15, 
    2.976813e-15, 2.974785e-15, 2.981042e-15, 2.987699e-15, 2.987844e-15, 
    2.989975e-15, 2.995977e-15, 2.985653e-15, 3.01759e-15, 2.997877e-15, 
    2.968363e-15, 2.974432e-15, 2.975301e-15, 2.972951e-15, 2.988892e-15, 
    2.983119e-15, 2.998655e-15, 2.99446e-15, 3.001334e-15, 2.997919e-15, 
    2.997416e-15, 2.993028e-15, 2.990293e-15, 2.983383e-15, 2.977756e-15, 
    2.973292e-15, 2.974331e-15, 2.979233e-15, 2.988107e-15, 2.996492e-15, 
    2.994655e-15, 3.000812e-15, 2.984512e-15, 2.991349e-15, 2.988707e-15, 
    2.995596e-15, 2.980494e-15, 2.993348e-15, 2.977204e-15, 2.978622e-15, 
    2.983005e-15, 2.99181e-15, 2.993762e-15, 2.99584e-15, 2.994558e-15, 
    2.988332e-15, 2.987313e-15, 2.982899e-15, 2.981678e-15, 2.978313e-15, 
    2.975525e-15, 2.978072e-15, 2.980745e-15, 2.988336e-15, 2.995167e-15, 
    3.002611e-15, 3.004433e-15, 3.013111e-15, 3.006043e-15, 3.017699e-15, 
    3.007785e-15, 3.024941e-15, 2.994096e-15, 3.007499e-15, 2.983205e-15, 
    2.985827e-15, 2.990562e-15, 3.001421e-15, 2.995564e-15, 3.002415e-15, 
    2.987273e-15, 2.979401e-15, 2.977366e-15, 2.973563e-15, 2.977453e-15, 
    2.977137e-15, 2.980858e-15, 2.979662e-15, 2.988588e-15, 2.983795e-15, 
    2.997402e-15, 3.002362e-15, 3.016353e-15, 3.024914e-15, 3.033624e-15, 
    3.037464e-15, 3.038632e-15, 3.039121e-15 ;

 LITR2N_vr =
  1.532743e-05, 1.532741e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 
    1.53274e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 1.532743e-05, 
    1.532738e-05, 1.53274e-05, 1.532735e-05, 1.532737e-05, 1.532733e-05, 
    1.532736e-05, 1.532733e-05, 1.532733e-05, 1.532731e-05, 1.532732e-05, 
    1.53273e-05, 1.532731e-05, 1.532729e-05, 1.53273e-05, 1.53273e-05, 
    1.532731e-05, 1.53274e-05, 1.532738e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532737e-05, 1.532734e-05, 1.532735e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532733e-05, 
    1.532733e-05, 1.532734e-05, 1.532737e-05, 1.532736e-05, 1.532739e-05, 
    1.532741e-05, 1.532742e-05, 1.532743e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 
    1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532731e-05, 1.532733e-05, 
    1.532732e-05, 1.532734e-05, 1.532734e-05, 1.532738e-05, 1.53274e-05, 
    1.532741e-05, 1.532741e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 
    1.532736e-05, 1.532737e-05, 1.532733e-05, 1.532734e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532731e-05, 1.532731e-05, 
    1.532731e-05, 1.53273e-05, 1.532733e-05, 1.532732e-05, 1.532741e-05, 
    1.532741e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532734e-05, 1.532733e-05, 
    1.532734e-05, 1.532733e-05, 1.532734e-05, 1.532734e-05, 1.532731e-05, 
    1.532733e-05, 1.53273e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.532741e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532743e-05, 
    1.532742e-05, 1.532742e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.532731e-05, 1.532741e-05, 1.532741e-05, 1.532741e-05, 1.53274e-05, 
    1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532736e-05, 1.532737e-05, 
    1.532736e-05, 1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532737e-05, 
    1.532734e-05, 1.532736e-05, 1.532732e-05, 1.532734e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 
    1.53273e-05, 1.532729e-05, 1.53274e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532736e-05, 
    1.532734e-05, 1.532734e-05, 1.532736e-05, 1.532735e-05, 1.532739e-05, 
    1.532738e-05, 1.532738e-05, 1.53274e-05, 1.532736e-05, 1.532738e-05, 
    1.532734e-05, 1.532735e-05, 1.532732e-05, 1.532733e-05, 1.53273e-05, 
    1.532729e-05, 1.532727e-05, 1.532726e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532735e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532733e-05, 1.532734e-05, 1.532733e-05, 
    1.532738e-05, 1.532735e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 
    1.532738e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 
    1.532729e-05, 1.532731e-05, 1.532724e-05, 1.532726e-05, 1.532739e-05, 
    1.532739e-05, 1.532737e-05, 1.532738e-05, 1.532735e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532733e-05, 
    1.532732e-05, 1.532735e-05, 1.532734e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532735e-05, 1.532729e-05, 1.532732e-05, 
    1.532738e-05, 1.532737e-05, 1.532737e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.532734e-05, 1.532735e-05, 1.532736e-05, 
    1.532737e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532733e-05, 1.532732e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532736e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532733e-05, 
    1.532734e-05, 1.532734e-05, 1.532735e-05, 1.532736e-05, 1.532736e-05, 
    1.532737e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532733e-05, 
    1.532732e-05, 1.532731e-05, 1.532729e-05, 1.532731e-05, 1.532729e-05, 
    1.53273e-05, 1.532727e-05, 1.532733e-05, 1.53273e-05, 1.532735e-05, 
    1.532735e-05, 1.532734e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532734e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532732e-05, 1.532732e-05, 1.532729e-05, 1.532727e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532724e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.063863e-13, 1.066744e-13, 1.066185e-13, 1.068506e-13, 1.067219e-13, 
    1.068739e-13, 1.064448e-13, 1.066858e-13, 1.06532e-13, 1.064123e-13, 
    1.073005e-13, 1.06861e-13, 1.077567e-13, 1.074769e-13, 1.081794e-13, 
    1.077131e-13, 1.082733e-13, 1.08166e-13, 1.084891e-13, 1.083966e-13, 
    1.088091e-13, 1.085317e-13, 1.090228e-13, 1.087429e-13, 1.087867e-13, 
    1.085226e-13, 1.069496e-13, 1.072458e-13, 1.06932e-13, 1.069743e-13, 
    1.069553e-13, 1.067245e-13, 1.066081e-13, 1.063643e-13, 1.064086e-13, 
    1.065877e-13, 1.069933e-13, 1.068557e-13, 1.072025e-13, 1.071946e-13, 
    1.075801e-13, 1.074064e-13, 1.080535e-13, 1.078698e-13, 1.084004e-13, 
    1.08267e-13, 1.083941e-13, 1.083556e-13, 1.083946e-13, 1.08199e-13, 
    1.082828e-13, 1.081106e-13, 1.074389e-13, 1.076365e-13, 1.070467e-13, 
    1.066914e-13, 1.064553e-13, 1.062877e-13, 1.063114e-13, 1.063565e-13, 
    1.065887e-13, 1.068069e-13, 1.069731e-13, 1.070841e-13, 1.071935e-13, 
    1.075242e-13, 1.076992e-13, 1.080905e-13, 1.0802e-13, 1.081395e-13, 
    1.082538e-13, 1.084453e-13, 1.084138e-13, 1.084982e-13, 1.081364e-13, 
    1.083769e-13, 1.079799e-13, 1.080885e-13, 1.072229e-13, 1.068929e-13, 
    1.067522e-13, 1.066292e-13, 1.063296e-13, 1.065365e-13, 1.06455e-13, 
    1.06649e-13, 1.067722e-13, 1.067113e-13, 1.070872e-13, 1.069411e-13, 
    1.077096e-13, 1.073788e-13, 1.082404e-13, 1.080345e-13, 1.082898e-13, 
    1.081596e-13, 1.083826e-13, 1.081819e-13, 1.085296e-13, 1.086052e-13, 
    1.085535e-13, 1.087521e-13, 1.081707e-13, 1.083941e-13, 1.067096e-13, 
    1.067195e-13, 1.067658e-13, 1.065622e-13, 1.065498e-13, 1.063631e-13, 
    1.065292e-13, 1.065999e-13, 1.067794e-13, 1.068854e-13, 1.069862e-13, 
    1.072077e-13, 1.074548e-13, 1.078001e-13, 1.080479e-13, 1.082138e-13, 
    1.081121e-13, 1.082019e-13, 1.081015e-13, 1.080544e-13, 1.085768e-13, 
    1.082836e-13, 1.087235e-13, 1.086992e-13, 1.085002e-13, 1.08702e-13, 
    1.067265e-13, 1.066693e-13, 1.064706e-13, 1.066261e-13, 1.063428e-13, 
    1.065014e-13, 1.065925e-13, 1.069441e-13, 1.070213e-13, 1.070928e-13, 
    1.072341e-13, 1.074153e-13, 1.077327e-13, 1.080087e-13, 1.082604e-13, 
    1.08242e-13, 1.082485e-13, 1.083047e-13, 1.081654e-13, 1.083275e-13, 
    1.083547e-13, 1.082836e-13, 1.08696e-13, 1.085782e-13, 1.086987e-13, 
    1.086221e-13, 1.066879e-13, 1.067841e-13, 1.067321e-13, 1.068299e-13, 
    1.06761e-13, 1.07067e-13, 1.071587e-13, 1.075875e-13, 1.074117e-13, 
    1.076915e-13, 1.074401e-13, 1.074847e-13, 1.077005e-13, 1.074538e-13, 
    1.079935e-13, 1.076276e-13, 1.083068e-13, 1.079418e-13, 1.083297e-13, 
    1.082593e-13, 1.083759e-13, 1.084801e-13, 1.086113e-13, 1.088531e-13, 
    1.087971e-13, 1.089993e-13, 1.069275e-13, 1.070522e-13, 1.070413e-13, 
    1.071717e-13, 1.072681e-13, 1.07477e-13, 1.078117e-13, 1.076859e-13, 
    1.079168e-13, 1.079632e-13, 1.076123e-13, 1.078277e-13, 1.071356e-13, 
    1.072475e-13, 1.071809e-13, 1.069373e-13, 1.077148e-13, 1.07316e-13, 
    1.080519e-13, 1.078363e-13, 1.084653e-13, 1.081526e-13, 1.087663e-13, 
    1.090281e-13, 1.092745e-13, 1.095619e-13, 1.071202e-13, 1.070356e-13, 
    1.071872e-13, 1.073968e-13, 1.075912e-13, 1.078495e-13, 1.078759e-13, 
    1.079242e-13, 1.080494e-13, 1.081546e-13, 1.079395e-13, 1.08181e-13, 
    1.072733e-13, 1.077494e-13, 1.070035e-13, 1.072282e-13, 1.073845e-13, 
    1.07316e-13, 1.076715e-13, 1.077552e-13, 1.080951e-13, 1.079195e-13, 
    1.089634e-13, 1.085021e-13, 1.097807e-13, 1.094239e-13, 1.07006e-13, 
    1.0712e-13, 1.075163e-13, 1.073278e-13, 1.078667e-13, 1.079992e-13, 
    1.081068e-13, 1.082443e-13, 1.082592e-13, 1.083407e-13, 1.082072e-13, 
    1.083354e-13, 1.0785e-13, 1.08067e-13, 1.074711e-13, 1.076163e-13, 
    1.075495e-13, 1.074763e-13, 1.077023e-13, 1.079428e-13, 1.079481e-13, 
    1.080251e-13, 1.082419e-13, 1.078689e-13, 1.090227e-13, 1.083105e-13, 
    1.072443e-13, 1.074635e-13, 1.074949e-13, 1.0741e-13, 1.079859e-13, 
    1.077774e-13, 1.083387e-13, 1.081871e-13, 1.084354e-13, 1.083121e-13, 
    1.082939e-13, 1.081353e-13, 1.080366e-13, 1.077869e-13, 1.075836e-13, 
    1.074223e-13, 1.074598e-13, 1.07637e-13, 1.079576e-13, 1.082605e-13, 
    1.081942e-13, 1.084166e-13, 1.078277e-13, 1.080747e-13, 1.079793e-13, 
    1.082281e-13, 1.076825e-13, 1.081469e-13, 1.075637e-13, 1.076149e-13, 
    1.077732e-13, 1.080914e-13, 1.081619e-13, 1.082369e-13, 1.081907e-13, 
    1.079657e-13, 1.079289e-13, 1.077694e-13, 1.077253e-13, 1.076037e-13, 
    1.07503e-13, 1.07595e-13, 1.076916e-13, 1.079659e-13, 1.082127e-13, 
    1.084816e-13, 1.085474e-13, 1.088609e-13, 1.086056e-13, 1.090267e-13, 
    1.086685e-13, 1.092883e-13, 1.081739e-13, 1.086582e-13, 1.077805e-13, 
    1.078752e-13, 1.080463e-13, 1.084386e-13, 1.08227e-13, 1.084745e-13, 
    1.079275e-13, 1.07643e-13, 1.075695e-13, 1.074321e-13, 1.075727e-13, 
    1.075612e-13, 1.076957e-13, 1.076525e-13, 1.07975e-13, 1.078018e-13, 
    1.082934e-13, 1.084726e-13, 1.089781e-13, 1.092874e-13, 1.096021e-13, 
    1.097408e-13, 1.09783e-13, 1.098007e-13 ;

 LITR3C =
  9.697999e-06, 9.69799e-06, 9.697992e-06, 9.697984e-06, 9.697988e-06, 
    9.697983e-06, 9.697997e-06, 9.697989e-06, 9.697995e-06, 9.697998e-06, 
    9.697968e-06, 9.697984e-06, 9.697953e-06, 9.697963e-06, 9.697939e-06, 
    9.697955e-06, 9.697936e-06, 9.697939e-06, 9.697928e-06, 9.697931e-06, 
    9.697917e-06, 9.697927e-06, 9.69791e-06, 9.69792e-06, 9.697918e-06, 
    9.697927e-06, 9.69798e-06, 9.69797e-06, 9.697981e-06, 9.697979e-06, 
    9.69798e-06, 9.697988e-06, 9.697992e-06, 9.698e-06, 9.697999e-06, 
    9.697993e-06, 9.697979e-06, 9.697984e-06, 9.697972e-06, 9.697972e-06, 
    9.697959e-06, 9.697965e-06, 9.697943e-06, 9.697949e-06, 9.697931e-06, 
    9.697936e-06, 9.697932e-06, 9.697933e-06, 9.697932e-06, 9.697938e-06, 
    9.697936e-06, 9.697941e-06, 9.697964e-06, 9.697957e-06, 9.697977e-06, 
    9.697989e-06, 9.697997e-06, 9.698003e-06, 9.698002e-06, 9.698e-06, 
    9.697993e-06, 9.697986e-06, 9.697979e-06, 9.697976e-06, 9.697972e-06, 
    9.697961e-06, 9.697955e-06, 9.697942e-06, 9.697944e-06, 9.69794e-06, 
    9.697937e-06, 9.69793e-06, 9.697931e-06, 9.697928e-06, 9.69794e-06, 
    9.697932e-06, 9.697946e-06, 9.697942e-06, 9.697971e-06, 9.697982e-06, 
    9.697987e-06, 9.697991e-06, 9.698001e-06, 9.697995e-06, 9.697997e-06, 
    9.697991e-06, 9.697987e-06, 9.697988e-06, 9.697976e-06, 9.697981e-06, 
    9.697955e-06, 9.697966e-06, 9.697937e-06, 9.697944e-06, 9.697935e-06, 
    9.697939e-06, 9.697932e-06, 9.697938e-06, 9.697927e-06, 9.697925e-06, 
    9.697927e-06, 9.697919e-06, 9.697939e-06, 9.697932e-06, 9.697988e-06, 
    9.697988e-06, 9.697987e-06, 9.697994e-06, 9.697994e-06, 9.698e-06, 
    9.697995e-06, 9.697992e-06, 9.697987e-06, 9.697983e-06, 9.697979e-06, 
    9.697972e-06, 9.697964e-06, 9.697952e-06, 9.697943e-06, 9.697937e-06, 
    9.697941e-06, 9.697938e-06, 9.697941e-06, 9.697943e-06, 9.697926e-06, 
    9.697936e-06, 9.69792e-06, 9.697921e-06, 9.697928e-06, 9.697921e-06, 
    9.697988e-06, 9.69799e-06, 9.697997e-06, 9.697991e-06, 9.698001e-06, 
    9.697996e-06, 9.697993e-06, 9.697981e-06, 9.697978e-06, 9.697976e-06, 
    9.697971e-06, 9.697965e-06, 9.697954e-06, 9.697945e-06, 9.697937e-06, 
    9.697937e-06, 9.697937e-06, 9.697935e-06, 9.697939e-06, 9.697934e-06, 
    9.697933e-06, 9.697936e-06, 9.697921e-06, 9.697926e-06, 9.697921e-06, 
    9.697924e-06, 9.697989e-06, 9.697987e-06, 9.697987e-06, 9.697985e-06, 
    9.697987e-06, 9.697977e-06, 9.697974e-06, 9.697959e-06, 9.697965e-06, 
    9.697956e-06, 9.697964e-06, 9.697962e-06, 9.697955e-06, 9.697964e-06, 
    9.697945e-06, 9.697957e-06, 9.697935e-06, 9.697947e-06, 9.697934e-06, 
    9.697937e-06, 9.697932e-06, 9.697928e-06, 9.697924e-06, 9.697916e-06, 
    9.697918e-06, 9.697911e-06, 9.697981e-06, 9.697977e-06, 9.697977e-06, 
    9.697973e-06, 9.697969e-06, 9.697963e-06, 9.697951e-06, 9.697956e-06, 
    9.697947e-06, 9.697947e-06, 9.697958e-06, 9.697951e-06, 9.697974e-06, 
    9.69797e-06, 9.697973e-06, 9.697981e-06, 9.697955e-06, 9.697968e-06, 
    9.697943e-06, 9.69795e-06, 9.697929e-06, 9.69794e-06, 9.697919e-06, 
    9.69791e-06, 9.697902e-06, 9.697892e-06, 9.697975e-06, 9.697977e-06, 
    9.697973e-06, 9.697966e-06, 9.697958e-06, 9.69795e-06, 9.697949e-06, 
    9.697947e-06, 9.697943e-06, 9.697939e-06, 9.697947e-06, 9.697938e-06, 
    9.697969e-06, 9.697954e-06, 9.697978e-06, 9.697971e-06, 9.697966e-06, 
    9.697968e-06, 9.697956e-06, 9.697953e-06, 9.697942e-06, 9.697947e-06, 
    9.697912e-06, 9.697928e-06, 9.697885e-06, 9.697897e-06, 9.697978e-06, 
    9.697975e-06, 9.697961e-06, 9.697967e-06, 9.697949e-06, 9.697945e-06, 
    9.697941e-06, 9.697937e-06, 9.697937e-06, 9.697934e-06, 9.697937e-06, 
    9.697934e-06, 9.69795e-06, 9.697943e-06, 9.697963e-06, 9.697958e-06, 
    9.69796e-06, 9.697963e-06, 9.697955e-06, 9.697947e-06, 9.697947e-06, 
    9.697944e-06, 9.697937e-06, 9.697949e-06, 9.69791e-06, 9.697935e-06, 
    9.69797e-06, 9.697963e-06, 9.697962e-06, 9.697965e-06, 9.697946e-06, 
    9.697953e-06, 9.697934e-06, 9.697938e-06, 9.69793e-06, 9.697935e-06, 
    9.697935e-06, 9.69794e-06, 9.697944e-06, 9.697952e-06, 9.697959e-06, 
    9.697965e-06, 9.697963e-06, 9.697957e-06, 9.697947e-06, 9.697937e-06, 
    9.697938e-06, 9.697931e-06, 9.697951e-06, 9.697942e-06, 9.697946e-06, 
    9.697937e-06, 9.697956e-06, 9.69794e-06, 9.697959e-06, 9.697958e-06, 
    9.697953e-06, 9.697942e-06, 9.697939e-06, 9.697937e-06, 9.697938e-06, 
    9.697946e-06, 9.697947e-06, 9.697953e-06, 9.697954e-06, 9.697958e-06, 
    9.697962e-06, 9.697958e-06, 9.697956e-06, 9.697946e-06, 9.697937e-06, 
    9.697928e-06, 9.697927e-06, 9.697916e-06, 9.697925e-06, 9.69791e-06, 
    9.697922e-06, 9.697901e-06, 9.697939e-06, 9.697923e-06, 9.697952e-06, 
    9.697949e-06, 9.697943e-06, 9.69793e-06, 9.697937e-06, 9.697929e-06, 
    9.697947e-06, 9.697957e-06, 9.697959e-06, 9.697964e-06, 9.697959e-06, 
    9.69796e-06, 9.697956e-06, 9.697957e-06, 9.697946e-06, 9.697952e-06, 
    9.697935e-06, 9.697929e-06, 9.697912e-06, 9.697901e-06, 9.697891e-06, 
    9.697886e-06, 9.697885e-06, 9.697884e-06 ;

 LITR3C_TO_SOIL2C =
  5.319314e-14, 5.33372e-14, 5.330921e-14, 5.34253e-14, 5.336093e-14, 
    5.343692e-14, 5.322238e-14, 5.33429e-14, 5.326598e-14, 5.320614e-14, 
    5.365024e-14, 5.343048e-14, 5.387835e-14, 5.373844e-14, 5.408968e-14, 
    5.385656e-14, 5.413665e-14, 5.408301e-14, 5.424451e-14, 5.419827e-14, 
    5.440452e-14, 5.426585e-14, 5.45114e-14, 5.437145e-14, 5.439333e-14, 
    5.426127e-14, 5.347478e-14, 5.362289e-14, 5.346599e-14, 5.348713e-14, 
    5.347765e-14, 5.336225e-14, 5.330402e-14, 5.318215e-14, 5.320429e-14, 
    5.329382e-14, 5.349663e-14, 5.342785e-14, 5.360122e-14, 5.359731e-14, 
    5.379004e-14, 5.370317e-14, 5.402671e-14, 5.393486e-14, 5.42002e-14, 
    5.41335e-14, 5.419706e-14, 5.41778e-14, 5.419731e-14, 5.409948e-14, 
    5.41414e-14, 5.40553e-14, 5.371944e-14, 5.381822e-14, 5.352335e-14, 
    5.334567e-14, 5.322766e-14, 5.314382e-14, 5.315567e-14, 5.317826e-14, 
    5.329434e-14, 5.340344e-14, 5.348651e-14, 5.354204e-14, 5.359674e-14, 
    5.376206e-14, 5.384959e-14, 5.404526e-14, 5.401e-14, 5.406975e-14, 
    5.412687e-14, 5.422265e-14, 5.42069e-14, 5.424907e-14, 5.406821e-14, 
    5.418842e-14, 5.398994e-14, 5.404423e-14, 5.361145e-14, 5.344641e-14, 
    5.337607e-14, 5.331459e-14, 5.316478e-14, 5.326824e-14, 5.322746e-14, 
    5.33245e-14, 5.338609e-14, 5.335564e-14, 5.354356e-14, 5.347052e-14, 
    5.385477e-14, 5.36894e-14, 5.412021e-14, 5.401724e-14, 5.414488e-14, 
    5.407977e-14, 5.41913e-14, 5.409093e-14, 5.426478e-14, 5.430258e-14, 
    5.427674e-14, 5.437603e-14, 5.408536e-14, 5.419704e-14, 5.335478e-14, 
    5.335975e-14, 5.33829e-14, 5.328108e-14, 5.327486e-14, 5.318154e-14, 
    5.32646e-14, 5.329994e-14, 5.338968e-14, 5.34427e-14, 5.34931e-14, 
    5.360385e-14, 5.37274e-14, 5.390003e-14, 5.402392e-14, 5.410691e-14, 
    5.405604e-14, 5.410095e-14, 5.405073e-14, 5.40272e-14, 5.42884e-14, 
    5.414178e-14, 5.436175e-14, 5.434959e-14, 5.425006e-14, 5.435096e-14, 
    5.336323e-14, 5.333465e-14, 5.32353e-14, 5.331305e-14, 5.317138e-14, 
    5.325068e-14, 5.329624e-14, 5.347202e-14, 5.351065e-14, 5.35464e-14, 
    5.361704e-14, 5.370762e-14, 5.386636e-14, 5.400432e-14, 5.41302e-14, 
    5.412098e-14, 5.412423e-14, 5.415231e-14, 5.40827e-14, 5.416374e-14, 
    5.417732e-14, 5.414178e-14, 5.434796e-14, 5.42891e-14, 5.434933e-14, 
    5.431101e-14, 5.334395e-14, 5.339205e-14, 5.336605e-14, 5.341492e-14, 
    5.338048e-14, 5.353351e-14, 5.357935e-14, 5.379372e-14, 5.370583e-14, 
    5.384573e-14, 5.372006e-14, 5.374233e-14, 5.385022e-14, 5.372686e-14, 
    5.399672e-14, 5.381376e-14, 5.41534e-14, 5.397088e-14, 5.416483e-14, 
    5.412965e-14, 5.418791e-14, 5.424005e-14, 5.430564e-14, 5.442653e-14, 
    5.439855e-14, 5.449962e-14, 5.346375e-14, 5.352607e-14, 5.352061e-14, 
    5.358583e-14, 5.363403e-14, 5.373849e-14, 5.390583e-14, 5.384294e-14, 
    5.395841e-14, 5.398157e-14, 5.380615e-14, 5.391385e-14, 5.356779e-14, 
    5.362372e-14, 5.359045e-14, 5.346865e-14, 5.385739e-14, 5.365801e-14, 
    5.402596e-14, 5.391815e-14, 5.423261e-14, 5.407626e-14, 5.438314e-14, 
    5.451403e-14, 5.463725e-14, 5.478092e-14, 5.356011e-14, 5.351777e-14, 
    5.359359e-14, 5.369837e-14, 5.379561e-14, 5.392472e-14, 5.393794e-14, 
    5.396211e-14, 5.402469e-14, 5.407729e-14, 5.396972e-14, 5.409048e-14, 
    5.363663e-14, 5.38747e-14, 5.350173e-14, 5.36141e-14, 5.369221e-14, 
    5.365799e-14, 5.383576e-14, 5.387761e-14, 5.404752e-14, 5.395974e-14, 
    5.448171e-14, 5.425101e-14, 5.489031e-14, 5.471195e-14, 5.350296e-14, 
    5.355997e-14, 5.375815e-14, 5.36639e-14, 5.393336e-14, 5.399959e-14, 
    5.40534e-14, 5.412215e-14, 5.412959e-14, 5.417031e-14, 5.410358e-14, 
    5.416769e-14, 5.3925e-14, 5.403349e-14, 5.373555e-14, 5.380812e-14, 
    5.377475e-14, 5.373812e-14, 5.385114e-14, 5.39714e-14, 5.397402e-14, 
    5.401252e-14, 5.412095e-14, 5.393445e-14, 5.451136e-14, 5.415526e-14, 
    5.362211e-14, 5.373173e-14, 5.374744e-14, 5.370498e-14, 5.399295e-14, 
    5.388867e-14, 5.416932e-14, 5.409353e-14, 5.42177e-14, 5.415601e-14, 
    5.414693e-14, 5.406766e-14, 5.401827e-14, 5.389344e-14, 5.379179e-14, 
    5.371115e-14, 5.372991e-14, 5.381847e-14, 5.397877e-14, 5.413024e-14, 
    5.409706e-14, 5.420827e-14, 5.391383e-14, 5.403733e-14, 5.398961e-14, 
    5.411406e-14, 5.384125e-14, 5.407344e-14, 5.378182e-14, 5.380743e-14, 
    5.38866e-14, 5.404567e-14, 5.408092e-14, 5.411846e-14, 5.409531e-14, 
    5.398284e-14, 5.396443e-14, 5.388469e-14, 5.386264e-14, 5.380185e-14, 
    5.375148e-14, 5.379749e-14, 5.384578e-14, 5.398291e-14, 5.410631e-14, 
    5.424078e-14, 5.427369e-14, 5.443046e-14, 5.430278e-14, 5.451333e-14, 
    5.433424e-14, 5.464416e-14, 5.408696e-14, 5.432907e-14, 5.389022e-14, 
    5.393758e-14, 5.402312e-14, 5.421929e-14, 5.411347e-14, 5.423724e-14, 
    5.396371e-14, 5.38215e-14, 5.378475e-14, 5.371604e-14, 5.378632e-14, 
    5.378061e-14, 5.384782e-14, 5.382623e-14, 5.398746e-14, 5.390088e-14, 
    5.414669e-14, 5.423628e-14, 5.448901e-14, 5.464368e-14, 5.480101e-14, 
    5.487038e-14, 5.489149e-14, 5.490031e-14 ;

 LITR3C_vr =
  0.0005537658, 0.0005537652, 0.0005537653, 0.0005537649, 0.0005537652, 
    0.0005537649, 0.0005537657, 0.0005537652, 0.0005537655, 0.0005537657, 
    0.0005537641, 0.0005537649, 0.0005537631, 0.0005537637, 0.0005537623, 
    0.0005537632, 0.0005537621, 0.0005537624, 0.0005537617, 0.0005537619, 
    0.0005537611, 0.0005537617, 0.0005537607, 0.0005537613, 0.0005537611, 
    0.0005537617, 0.0005537647, 0.0005537641, 0.0005537648, 0.0005537646, 
    0.0005537647, 0.0005537652, 0.0005537654, 0.0005537659, 0.0005537657, 
    0.0005537654, 0.0005537646, 0.0005537649, 0.0005537642, 0.0005537642, 
    0.0005537635, 0.0005537638, 0.0005537626, 0.0005537629, 0.0005537619, 
    0.0005537621, 0.0005537619, 0.000553762, 0.0005537619, 0.0005537623, 
    0.0005537621, 0.0005537625, 0.0005537638, 0.0005537634, 0.0005537645, 
    0.0005537652, 0.0005537657, 0.000553766, 0.0005537659, 0.0005537659, 
    0.0005537654, 0.000553765, 0.0005537646, 0.0005537645, 0.0005537642, 
    0.0005537636, 0.0005537632, 0.0005537625, 0.0005537627, 0.0005537624, 
    0.0005537622, 0.0005537618, 0.0005537619, 0.0005537617, 0.0005537624, 
    0.000553762, 0.0005537627, 0.0005537625, 0.0005537642, 0.0005537648, 
    0.0005537651, 0.0005537653, 0.0005537659, 0.0005537655, 0.0005537657, 
    0.0005537653, 0.000553765, 0.0005537652, 0.0005537645, 0.0005537648, 
    0.0005537632, 0.0005537639, 0.0005537622, 0.0005537626, 0.0005537621, 
    0.0005537624, 0.000553762, 0.0005537623, 0.0005537617, 0.0005537615, 
    0.0005537616, 0.0005537612, 0.0005537624, 0.0005537619, 0.0005537652, 
    0.0005537652, 0.000553765, 0.0005537655, 0.0005537655, 0.0005537659, 
    0.0005537655, 0.0005537654, 0.000553765, 0.0005537648, 0.0005537646, 
    0.0005537642, 0.0005537637, 0.0005537631, 0.0005537626, 0.0005537622, 
    0.0005537625, 0.0005537623, 0.0005537625, 0.0005537626, 0.0005537616, 
    0.0005537621, 0.0005537613, 0.0005537613, 0.0005537617, 0.0005537613, 
    0.0005537652, 0.0005537653, 0.0005537656, 0.0005537653, 0.0005537659, 
    0.0005537656, 0.0005537654, 0.0005537647, 0.0005537646, 0.0005537645, 
    0.0005537642, 0.0005537638, 0.0005537632, 0.0005537627, 0.0005537622, 
    0.0005537622, 0.0005537622, 0.0005537621, 0.0005537624, 0.000553762, 
    0.000553762, 0.0005537621, 0.0005537613, 0.0005537616, 0.0005537613, 
    0.0005537615, 0.0005537652, 0.000553765, 0.0005537651, 0.0005537649, 
    0.0005537651, 0.0005537645, 0.0005537643, 0.0005537635, 0.0005537638, 
    0.0005537633, 0.0005537638, 0.0005537636, 0.0005537632, 0.0005537638, 
    0.0005537627, 0.0005537634, 0.0005537621, 0.0005537628, 0.000553762, 
    0.0005537622, 0.000553762, 0.0005537617, 0.0005537615, 0.000553761, 
    0.0005537611, 0.0005537607, 0.0005537648, 0.0005537645, 0.0005537645, 
    0.0005537643, 0.0005537641, 0.0005537637, 0.0005537631, 0.0005537633, 
    0.0005537628, 0.0005537628, 0.0005537634, 0.000553763, 0.0005537643, 
    0.0005537641, 0.0005537643, 0.0005537648, 0.0005537632, 0.000553764, 
    0.0005537626, 0.000553763, 0.0005537618, 0.0005537624, 0.0005537612, 
    0.0005537607, 0.0005537602, 0.0005537596, 0.0005537644, 0.0005537645, 
    0.0005537642, 0.0005537638, 0.0005537635, 0.0005537629, 0.0005537629, 
    0.0005537628, 0.0005537626, 0.0005537624, 0.0005537628, 0.0005537623, 
    0.0005537641, 0.0005537632, 0.0005537646, 0.0005537642, 0.0005537639, 
    0.000553764, 0.0005537633, 0.0005537631, 0.0005537625, 0.0005537628, 
    0.0005537608, 0.0005537617, 0.0005537592, 0.0005537599, 0.0005537646, 
    0.0005537644, 0.0005537636, 0.000553764, 0.0005537629, 0.0005537627, 
    0.0005537625, 0.0005537622, 0.0005537622, 0.000553762, 0.0005537622, 
    0.000553762, 0.0005537629, 0.0005537625, 0.0005537637, 0.0005537634, 
    0.0005537635, 0.0005537637, 0.0005537632, 0.0005537628, 0.0005537628, 
    0.0005537627, 0.0005537622, 0.0005537629, 0.0005537607, 0.0005537621, 
    0.0005537641, 0.0005537637, 0.0005537636, 0.0005537638, 0.0005537627, 
    0.0005537631, 0.000553762, 0.0005537623, 0.0005537618, 0.0005537621, 
    0.0005537621, 0.0005537624, 0.0005537626, 0.0005537631, 0.0005537635, 
    0.0005537638, 0.0005537637, 0.0005537634, 0.0005537628, 0.0005537622, 
    0.0005537623, 0.0005537619, 0.000553763, 0.0005537625, 0.0005537627, 
    0.0005537622, 0.0005537633, 0.0005537624, 0.0005537635, 0.0005537634, 
    0.0005537631, 0.0005537625, 0.0005537624, 0.0005537622, 0.0005537623, 
    0.0005537627, 0.0005537628, 0.0005537631, 0.0005537632, 0.0005537635, 
    0.0005537636, 0.0005537635, 0.0005537633, 0.0005537627, 0.0005537622, 
    0.0005537617, 0.0005537616, 0.000553761, 0.0005537615, 0.0005537607, 
    0.0005537614, 0.0005537602, 0.0005537624, 0.0005537614, 0.0005537631, 
    0.0005537629, 0.0005537626, 0.0005537618, 0.0005537622, 0.0005537618, 
    0.0005537628, 0.0005537634, 0.0005537635, 0.0005537638, 0.0005537635, 
    0.0005537635, 0.0005537632, 0.0005537634, 0.0005537627, 0.0005537631, 
    0.0005537621, 0.0005537618, 0.0005537608, 0.0005537602, 0.0005537596, 
    0.0005537593, 0.0005537592, 0.0005537592,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342132e-07, 1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 
    1.34213e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342128e-07, 1.34213e-07, 1.342126e-07, 1.342127e-07, 1.342124e-07, 
    1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 1.342123e-07, 
    1.342121e-07, 1.342122e-07, 1.34212e-07, 1.342121e-07, 1.342121e-07, 
    1.342122e-07, 1.34213e-07, 1.342128e-07, 1.34213e-07, 1.342129e-07, 
    1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342128e-07, 
    1.342127e-07, 1.342127e-07, 1.342124e-07, 1.342125e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 
    1.342123e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 1.342129e-07, 
    1.342131e-07, 1.342132e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 
    1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 1.342124e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342124e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342128e-07, 1.34213e-07, 
    1.342131e-07, 1.342131e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342131e-07, 1.342129e-07, 1.34213e-07, 
    1.342126e-07, 1.342128e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 1.342122e-07, 
    1.342122e-07, 1.342121e-07, 1.342124e-07, 1.342123e-07, 1.342131e-07, 
    1.342131e-07, 1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342124e-07, 1.342124e-07, 1.342124e-07, 1.342122e-07, 
    1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.342131e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.342122e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342129e-07, 1.342127e-07, 1.342127e-07, 
    1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 
    1.342125e-07, 1.342126e-07, 1.342123e-07, 1.342125e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342121e-07, 
    1.342121e-07, 1.34212e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342126e-07, 
    1.342125e-07, 1.342125e-07, 1.342126e-07, 1.342125e-07, 1.342129e-07, 
    1.342128e-07, 1.342128e-07, 1.34213e-07, 1.342126e-07, 1.342128e-07, 
    1.342124e-07, 1.342125e-07, 1.342122e-07, 1.342124e-07, 1.342121e-07, 
    1.34212e-07, 1.342119e-07, 1.342117e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342125e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342124e-07, 1.342125e-07, 1.342124e-07, 
    1.342128e-07, 1.342126e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342128e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 
    1.34212e-07, 1.342122e-07, 1.342116e-07, 1.342118e-07, 1.342129e-07, 
    1.342129e-07, 1.342127e-07, 1.342128e-07, 1.342125e-07, 1.342125e-07, 
    1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342124e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342124e-07, 1.342123e-07, 1.342125e-07, 1.34212e-07, 1.342123e-07, 
    1.342128e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 1.342125e-07, 
    1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 1.342123e-07, 
    1.342123e-07, 1.342124e-07, 1.342124e-07, 1.342126e-07, 1.342127e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342125e-07, 
    1.342124e-07, 1.342126e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 
    1.342125e-07, 1.342125e-07, 1.342126e-07, 1.342126e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342124e-07, 
    1.342122e-07, 1.342122e-07, 1.342121e-07, 1.342122e-07, 1.34212e-07, 
    1.342121e-07, 1.342119e-07, 1.342124e-07, 1.342122e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342122e-07, 
    1.342125e-07, 1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342126e-07, 1.342125e-07, 1.342126e-07, 
    1.342123e-07, 1.342122e-07, 1.34212e-07, 1.342119e-07, 1.342117e-07, 
    1.342116e-07, 1.342116e-07, 1.342116e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  4.043994e-26, 2.695996e-26, -2.32836e-26, -5.759628e-26, -4.289085e-26, 
    -7.842898e-26, 2.573451e-26, -1.311234e-25, -2.32836e-26, -3.921449e-26, 
    -5.514538e-26, 4.166539e-26, -9.435986e-26, 4.41163e-26, -7.352717e-27, 
    -4.901811e-26, 1.004871e-25, 2.450906e-27, -4.043994e-26, -4.289085e-26, 
    1.102908e-26, 9.558531e-26, 0, 2.450905e-26, -1.017126e-25, 3.676358e-26, 
    -2.08327e-26, 1.347998e-26, -1.041635e-25, -3.921449e-26, -7.352717e-26, 
    -3.676358e-27, -8.578169e-27, 4.901811e-26, 4.534175e-26, 1.593089e-25, 
    -9.068351e-26, 7.352717e-26, 7.230172e-26, -2.021997e-25, 3.553813e-26, 
    -4.534175e-26, -1.102908e-26, -6.4949e-26, -2.08327e-26, -3.921449e-26, 
    1.225453e-26, -2.450906e-27, -6.862535e-26, 4.779266e-26, 5.514538e-26, 
    -3.553813e-26, -6.862535e-26, 2.695996e-26, 3.676358e-27, 1.151926e-25, 
    2.205815e-26, -5.882173e-26, 7.352717e-27, 1.446034e-25, 2.32836e-26, 
    4.901811e-26, 1.225453e-27, -2.450906e-27, -4.41163e-26, -3.921449e-26, 
    1.752397e-25, -8.578169e-26, -6.372354e-26, -5.269447e-26, 1.960724e-26, 
    1.838179e-26, -1.715634e-26, -3.186177e-26, -1.838179e-26, 7.597807e-26, 
    3.676358e-26, 3.063632e-26, 1.102908e-25, 5.146902e-26, -2.573451e-26, 
    1.838179e-26, -9.068351e-26, 3.676358e-27, 4.043994e-26, 3.308722e-26, 
    -2.450905e-26, -8.945805e-26, 2.450905e-26, -3.431268e-26, 3.553813e-26, 
    9.803622e-27, -4.289085e-26, 7.352717e-26, 3.063632e-26, -7.352717e-26, 
    7.842898e-26, 3.308722e-26, -9.558531e-26, 1.225453e-25, -1.053889e-25, 
    6.4949e-26, 8.455624e-26, 6.617445e-26, -3.798904e-26, -7.720352e-26, 
    5.759628e-26, -1.838179e-26, 1.115162e-25, 5.514538e-26, -8.578169e-27, 
    -7.352717e-26, 3.553813e-26, 5.391992e-26, -8.333079e-26, 5.514538e-26, 
    -1.715634e-26, -1.066144e-25, 1.715634e-26, 1.225453e-27, 1.397016e-25, 
    -7.107626e-26, -4.65672e-26, -2.205815e-26, 2.450905e-26, -7.352717e-26, 
    2.450905e-26, -6.862535e-26, 4.901811e-27, -2.573451e-26, -2.450905e-26, 
    -9.435986e-26, -2.818541e-26, -6.372354e-26, -6.249809e-26, 
    -7.475262e-26, -1.519561e-25, -4.289085e-26, 2.573451e-26, 6.4949e-26, 
    -9.803622e-26, 4.65672e-26, -6.617445e-26, -1.225453e-27, -3.676358e-26, 
    -6.004719e-26, 2.08327e-26, -2.818541e-26, -3.186177e-26, 1.360253e-25, 
    1.102908e-25, -2.450906e-27, -6.127264e-26, -6.617445e-26, -5.759628e-26, 
    -4.901811e-27, -1.249962e-25, -1.960724e-26, -3.921449e-26, 6.127264e-26, 
    -4.41163e-26, -1.593089e-26, -3.063632e-26, -2.941087e-26, 9.803622e-27, 
    3.921449e-26, -2.941087e-26, -5.391992e-26, -6.249809e-26, 1.29898e-25, 
    -3.186177e-26, -1.262216e-25, -1.960724e-26, 1.237707e-25, -1.249962e-25, 
    -1.102908e-26, 7.352717e-27, 9.068351e-26, -8.087988e-26, 2.450905e-26, 
    2.450906e-27, -2.32836e-26, -1.041635e-25, -5.637083e-26, -2.32836e-26, 
    -4.289085e-26, 4.166539e-26, -6.372354e-26, 1.29898e-25, -3.798904e-26, 
    -5.024356e-26, -2.695996e-26, 6.4949e-26, -7.842898e-26, 1.593089e-26, 
    -5.637083e-26, 5.391992e-26, 5.759628e-26, 7.352717e-27, -1.066144e-25, 
    1.838179e-26, -4.901811e-27, 3.676358e-27, -1.838179e-26, -1.115162e-25, 
    2.818541e-26, 2.573451e-26, -1.078398e-25, 8.210533e-26, 9.803622e-26, 
    9.190896e-26, -3.676358e-27, -3.553813e-26, -2.450906e-27, 2.205815e-26, 
    4.901811e-27, 7.352717e-27, -1.225453e-27, 3.553813e-26, 1.347998e-26, 
    -2.365124e-25, -3.553813e-26, -8.087988e-26, 9.313441e-26, 5.024356e-26, 
    1.151926e-25, -1.960724e-26, -1.139671e-25, 3.676358e-26, -7.352717e-26, 
    1.470543e-25, -6.617445e-26, -2.450905e-26, 3.676358e-27, 2.32836e-26, 
    -5.269447e-26, -3.063632e-26, -4.779266e-26, 1.470543e-26, 6.127264e-27, 
    -4.534175e-26, 4.65672e-26, -2.205815e-26, -2.573451e-26, -1.225453e-26, 
    3.431268e-26, 5.637083e-26, 1.642107e-25, -5.024356e-26, -1.838179e-26, 
    -5.024356e-26, 1.053889e-25, -3.431268e-26, 6.127264e-27, -8.578169e-27, 
    5.637083e-26, 2.941087e-26, -1.593089e-26, -2.205815e-26, 4.65672e-26, 
    -5.759628e-26, 3.431268e-26, 6.127264e-26, -1.495052e-25, 5.637083e-26, 
    3.798904e-26, 3.798904e-26, 1.715634e-26, 1.715634e-26, 8.700715e-26, 
    1.715634e-26, 1.347998e-26, 2.818541e-26, -3.063632e-26, 1.593089e-26, 
    1.960724e-26, 9.435986e-26, -3.431268e-26, 8.82326e-26, -2.941087e-26, 
    -5.514538e-26, 6.73999e-26, -6.249809e-26, -9.803622e-26, 7.352717e-26, 
    1.838179e-26, 3.798904e-26, 2.818541e-26, -2.573451e-26, 1.838179e-25, 
    9.068351e-26, -7.230172e-26, -3.431268e-26, -1.102908e-26, -1.115162e-25, 
    1.225453e-26, -3.676358e-27, -7.352717e-26, 5.269447e-26, -6.127264e-26, 
    1.556325e-25, -6.127264e-27, 6.004719e-26, 7.352717e-27, 2.450906e-27, 
    -1.02938e-25, 9.803622e-27, 3.553813e-26, -7.475262e-26, 5.269447e-26, 
    3.921449e-26, 1.887197e-25, 1.102908e-26, -1.323489e-25, 7.352717e-26, 
    -6.249809e-26, 7.107626e-26, -7.230172e-26, -1.960724e-26, 6.73999e-26, 
    4.166539e-26, -4.166539e-26, 5.024356e-26, 6.617445e-26, -2.450905e-26, 
    -3.431268e-26, 4.65672e-26, 3.921449e-26, -9.803622e-26, 8.578169e-26, 
    -2.450905e-26, 4.043994e-26, -5.146902e-26, 6.004719e-26, 2.450906e-27, 
    -4.779266e-26, -8.210533e-26, -5.024356e-26,
  1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 
    1.338123e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338121e-32, 1.338123e-32, 1.338119e-32, 1.33812e-32, 1.338117e-32, 
    1.338119e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 1.338116e-32, 
    1.338114e-32, 1.338115e-32, 1.338113e-32, 1.338114e-32, 1.338114e-32, 
    1.338115e-32, 1.338123e-32, 1.338121e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338122e-32, 1.338123e-32, 1.338121e-32, 1.338121e-32, 
    1.33812e-32, 1.33812e-32, 1.338117e-32, 1.338118e-32, 1.338116e-32, 
    1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338117e-32, 
    1.338116e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 
    1.338124e-32, 1.338125e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 
    1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338117e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.338121e-32, 1.338123e-32, 
    1.338124e-32, 1.338124e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 
    1.338119e-32, 1.338121e-32, 1.338117e-32, 1.338118e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 1.338115e-32, 
    1.338115e-32, 1.338114e-32, 1.338117e-32, 1.338116e-32, 1.338124e-32, 
    1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 
    1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338115e-32, 
    1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338124e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338116e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338115e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 
    1.338124e-32, 1.338122e-32, 1.338122e-32, 1.33812e-32, 1.33812e-32, 
    1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.33812e-32, 
    1.338118e-32, 1.338119e-32, 1.338116e-32, 1.338118e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338114e-32, 
    1.338114e-32, 1.338113e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338119e-32, 
    1.338118e-32, 1.338118e-32, 1.338119e-32, 1.338119e-32, 1.338122e-32, 
    1.338121e-32, 1.338121e-32, 1.338123e-32, 1.338119e-32, 1.338121e-32, 
    1.338117e-32, 1.338118e-32, 1.338115e-32, 1.338117e-32, 1.338114e-32, 
    1.338113e-32, 1.338112e-32, 1.33811e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338117e-32, 
    1.338121e-32, 1.338119e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.338121e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338113e-32, 1.338115e-32, 1.338109e-32, 1.338111e-32, 1.338122e-32, 
    1.338122e-32, 1.33812e-32, 1.338121e-32, 1.338118e-32, 1.338118e-32, 
    1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338116e-32, 1.338117e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338118e-32, 1.338113e-32, 1.338116e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338118e-32, 
    1.338119e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.338118e-32, 1.338119e-32, 1.33812e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338117e-32, 1.338119e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 
    1.338118e-32, 1.338118e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 
    1.338115e-32, 1.338115e-32, 1.338114e-32, 1.338115e-32, 1.338113e-32, 
    1.338115e-32, 1.338112e-32, 1.338117e-32, 1.338115e-32, 1.338119e-32, 
    1.338118e-32, 1.338118e-32, 1.338116e-32, 1.338117e-32, 1.338115e-32, 
    1.338118e-32, 1.338119e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338118e-32, 1.338119e-32, 
    1.338116e-32, 1.338115e-32, 1.338113e-32, 1.338112e-32, 1.33811e-32, 
    1.338109e-32, 1.338109e-32, 1.338109e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.472308e-15, 1.476296e-15, 1.475521e-15, 1.478734e-15, 1.476953e-15, 
    1.479056e-15, 1.473118e-15, 1.476453e-15, 1.474324e-15, 1.472668e-15, 
    1.48496e-15, 1.478878e-15, 1.491274e-15, 1.487401e-15, 1.497123e-15, 
    1.490671e-15, 1.498423e-15, 1.496938e-15, 1.501409e-15, 1.500129e-15, 
    1.505838e-15, 1.501999e-15, 1.508796e-15, 1.504922e-15, 1.505528e-15, 
    1.501872e-15, 1.480104e-15, 1.484203e-15, 1.47986e-15, 1.480445e-15, 
    1.480183e-15, 1.476989e-15, 1.475377e-15, 1.472004e-15, 1.472617e-15, 
    1.475095e-15, 1.480708e-15, 1.478805e-15, 1.483603e-15, 1.483495e-15, 
    1.48883e-15, 1.486425e-15, 1.49538e-15, 1.492838e-15, 1.500182e-15, 
    1.498336e-15, 1.500095e-15, 1.499562e-15, 1.500102e-15, 1.497394e-15, 
    1.498555e-15, 1.496172e-15, 1.486875e-15, 1.48961e-15, 1.481448e-15, 
    1.47653e-15, 1.473264e-15, 1.470943e-15, 1.471271e-15, 1.471896e-15, 
    1.475109e-15, 1.478129e-15, 1.480428e-15, 1.481965e-15, 1.48348e-15, 
    1.488055e-15, 1.490478e-15, 1.495894e-15, 1.494918e-15, 1.496572e-15, 
    1.498153e-15, 1.500804e-15, 1.500368e-15, 1.501535e-15, 1.496529e-15, 
    1.499856e-15, 1.494362e-15, 1.495865e-15, 1.483886e-15, 1.479319e-15, 
    1.477371e-15, 1.47567e-15, 1.471523e-15, 1.474387e-15, 1.473258e-15, 
    1.475944e-15, 1.477649e-15, 1.476806e-15, 1.482007e-15, 1.479986e-15, 
    1.490621e-15, 1.486044e-15, 1.497968e-15, 1.495118e-15, 1.498651e-15, 
    1.496849e-15, 1.499936e-15, 1.497158e-15, 1.50197e-15, 1.503016e-15, 
    1.502301e-15, 1.505049e-15, 1.497004e-15, 1.500095e-15, 1.476782e-15, 
    1.47692e-15, 1.477561e-15, 1.474742e-15, 1.47457e-15, 1.471987e-15, 
    1.474286e-15, 1.475264e-15, 1.477748e-15, 1.479216e-15, 1.480611e-15, 
    1.483676e-15, 1.487096e-15, 1.491874e-15, 1.495303e-15, 1.4976e-15, 
    1.496192e-15, 1.497435e-15, 1.496045e-15, 1.495394e-15, 1.502624e-15, 
    1.498565e-15, 1.504654e-15, 1.504317e-15, 1.501563e-15, 1.504355e-15, 
    1.477016e-15, 1.476225e-15, 1.473475e-15, 1.475627e-15, 1.471706e-15, 
    1.473901e-15, 1.475162e-15, 1.480027e-15, 1.481096e-15, 1.482086e-15, 
    1.484041e-15, 1.486548e-15, 1.490942e-15, 1.494761e-15, 1.498245e-15, 
    1.49799e-15, 1.498079e-15, 1.498857e-15, 1.49693e-15, 1.499173e-15, 
    1.499549e-15, 1.498565e-15, 1.504272e-15, 1.502643e-15, 1.50431e-15, 
    1.503249e-15, 1.476482e-15, 1.477814e-15, 1.477094e-15, 1.478447e-15, 
    1.477494e-15, 1.481729e-15, 1.482998e-15, 1.488932e-15, 1.486499e-15, 
    1.490371e-15, 1.486893e-15, 1.487509e-15, 1.490495e-15, 1.487081e-15, 
    1.49455e-15, 1.489486e-15, 1.498887e-15, 1.493835e-15, 1.499203e-15, 
    1.49823e-15, 1.499842e-15, 1.501285e-15, 1.503101e-15, 1.506447e-15, 
    1.505672e-15, 1.50847e-15, 1.479798e-15, 1.481523e-15, 1.481372e-15, 
    1.483177e-15, 1.484512e-15, 1.487403e-15, 1.492035e-15, 1.490294e-15, 
    1.49349e-15, 1.494131e-15, 1.489275e-15, 1.492256e-15, 1.482678e-15, 
    1.484226e-15, 1.483305e-15, 1.479934e-15, 1.490694e-15, 1.485175e-15, 
    1.495359e-15, 1.492375e-15, 1.501079e-15, 1.496752e-15, 1.505246e-15, 
    1.508869e-15, 1.512279e-15, 1.516256e-15, 1.482465e-15, 1.481294e-15, 
    1.483392e-15, 1.486292e-15, 1.488984e-15, 1.492557e-15, 1.492923e-15, 
    1.493592e-15, 1.495324e-15, 1.49678e-15, 1.493803e-15, 1.497145e-15, 
    1.484584e-15, 1.491173e-15, 1.48085e-15, 1.48396e-15, 1.486122e-15, 
    1.485175e-15, 1.490095e-15, 1.491253e-15, 1.495956e-15, 1.493527e-15, 
    1.507974e-15, 1.501589e-15, 1.519284e-15, 1.514347e-15, 1.480884e-15, 
    1.482462e-15, 1.487947e-15, 1.485338e-15, 1.492796e-15, 1.49463e-15, 
    1.496119e-15, 1.498022e-15, 1.498228e-15, 1.499355e-15, 1.497508e-15, 
    1.499282e-15, 1.492565e-15, 1.495568e-15, 1.487322e-15, 1.48933e-15, 
    1.488406e-15, 1.487393e-15, 1.490521e-15, 1.49385e-15, 1.493922e-15, 
    1.494988e-15, 1.497989e-15, 1.492827e-15, 1.508795e-15, 1.498938e-15, 
    1.484182e-15, 1.487216e-15, 1.487651e-15, 1.486475e-15, 1.494446e-15, 
    1.49156e-15, 1.499328e-15, 1.49723e-15, 1.500667e-15, 1.498959e-15, 
    1.498708e-15, 1.496514e-15, 1.495147e-15, 1.491692e-15, 1.488878e-15, 
    1.486646e-15, 1.487165e-15, 1.489617e-15, 1.494053e-15, 1.498246e-15, 
    1.497328e-15, 1.500406e-15, 1.492256e-15, 1.495674e-15, 1.494354e-15, 
    1.497798e-15, 1.490247e-15, 1.496674e-15, 1.488602e-15, 1.489311e-15, 
    1.491502e-15, 1.495905e-15, 1.496881e-15, 1.49792e-15, 1.497279e-15, 
    1.494166e-15, 1.493656e-15, 1.491449e-15, 1.490839e-15, 1.489157e-15, 
    1.487763e-15, 1.489036e-15, 1.490372e-15, 1.494168e-15, 1.497584e-15, 
    1.501305e-15, 1.502216e-15, 1.506555e-15, 1.503022e-15, 1.508849e-15, 
    1.503892e-15, 1.51247e-15, 1.497048e-15, 1.503749e-15, 1.491602e-15, 
    1.492913e-15, 1.495281e-15, 1.500711e-15, 1.497782e-15, 1.501207e-15, 
    1.493637e-15, 1.4897e-15, 1.488683e-15, 1.486781e-15, 1.488727e-15, 
    1.488569e-15, 1.490429e-15, 1.489831e-15, 1.494294e-15, 1.491897e-15, 
    1.498701e-15, 1.501181e-15, 1.508176e-15, 1.512457e-15, 1.516812e-15, 
    1.518732e-15, 1.519316e-15, 1.51956e-15 ;

 LITR3N_vr =
  7.663713e-06, 7.663706e-06, 7.663707e-06, 7.663701e-06, 7.663704e-06, 
    7.663701e-06, 7.663712e-06, 7.663705e-06, 7.66371e-06, 7.663712e-06, 
    7.663689e-06, 7.663701e-06, 7.663677e-06, 7.663684e-06, 7.663665e-06, 
    7.663678e-06, 7.663662e-06, 7.663666e-06, 7.663657e-06, 7.66366e-06, 
    7.663649e-06, 7.663656e-06, 7.663642e-06, 7.663651e-06, 7.663649e-06, 
    7.663656e-06, 7.663698e-06, 7.663691e-06, 7.663699e-06, 7.663698e-06, 
    7.663698e-06, 7.663704e-06, 7.663708e-06, 7.663714e-06, 7.663712e-06, 
    7.663708e-06, 7.663697e-06, 7.663701e-06, 7.663692e-06, 7.663692e-06, 
    7.663682e-06, 7.663686e-06, 7.663669e-06, 7.663673e-06, 7.66366e-06, 
    7.663663e-06, 7.66366e-06, 7.663661e-06, 7.66366e-06, 7.663665e-06, 
    7.663662e-06, 7.663667e-06, 7.663685e-06, 7.66368e-06, 7.663696e-06, 
    7.663705e-06, 7.663712e-06, 7.663716e-06, 7.663715e-06, 7.663714e-06, 
    7.663708e-06, 7.663702e-06, 7.663698e-06, 7.663694e-06, 7.663692e-06, 
    7.663683e-06, 7.663678e-06, 7.663668e-06, 7.66367e-06, 7.663666e-06, 
    7.663663e-06, 7.663658e-06, 7.663659e-06, 7.663657e-06, 7.663666e-06, 
    7.66366e-06, 7.663671e-06, 7.663668e-06, 7.663691e-06, 7.6637e-06, 
    7.663703e-06, 7.663707e-06, 7.663715e-06, 7.66371e-06, 7.663712e-06, 
    7.663706e-06, 7.663703e-06, 7.663704e-06, 7.663694e-06, 7.663699e-06, 
    7.663678e-06, 7.663687e-06, 7.663663e-06, 7.663669e-06, 7.663662e-06, 
    7.663666e-06, 7.66366e-06, 7.663665e-06, 7.663656e-06, 7.663654e-06, 
    7.663655e-06, 7.66365e-06, 7.663665e-06, 7.66366e-06, 7.663705e-06, 
    7.663704e-06, 7.663703e-06, 7.663709e-06, 7.663709e-06, 7.663714e-06, 
    7.66371e-06, 7.663708e-06, 7.663702e-06, 7.6637e-06, 7.663697e-06, 
    7.663692e-06, 7.663685e-06, 7.663675e-06, 7.663669e-06, 7.663664e-06, 
    7.663667e-06, 7.663665e-06, 7.663667e-06, 7.663669e-06, 7.663654e-06, 
    7.663662e-06, 7.663651e-06, 7.663652e-06, 7.663657e-06, 7.663652e-06, 
    7.663704e-06, 7.663706e-06, 7.663712e-06, 7.663707e-06, 7.663714e-06, 
    7.663711e-06, 7.663708e-06, 7.663699e-06, 7.663696e-06, 7.663694e-06, 
    7.663691e-06, 7.663686e-06, 7.663677e-06, 7.66367e-06, 7.663663e-06, 
    7.663663e-06, 7.663663e-06, 7.663662e-06, 7.663666e-06, 7.663662e-06, 
    7.663661e-06, 7.663662e-06, 7.663652e-06, 7.663654e-06, 7.663652e-06, 
    7.663653e-06, 7.663705e-06, 7.663702e-06, 7.663704e-06, 7.663702e-06, 
    7.663703e-06, 7.663695e-06, 7.663692e-06, 7.663682e-06, 7.663686e-06, 
    7.663679e-06, 7.663685e-06, 7.663684e-06, 7.663678e-06, 7.663685e-06, 
    7.663671e-06, 7.66368e-06, 7.663662e-06, 7.663672e-06, 7.663662e-06, 
    7.663663e-06, 7.66366e-06, 7.663657e-06, 7.663653e-06, 7.663647e-06, 
    7.663649e-06, 7.663643e-06, 7.663699e-06, 7.663695e-06, 7.663696e-06, 
    7.663692e-06, 7.66369e-06, 7.663684e-06, 7.663675e-06, 7.663679e-06, 
    7.663672e-06, 7.663672e-06, 7.663681e-06, 7.663675e-06, 7.663693e-06, 
    7.663691e-06, 7.663692e-06, 7.663699e-06, 7.663678e-06, 7.663689e-06, 
    7.663669e-06, 7.663674e-06, 7.663658e-06, 7.663666e-06, 7.66365e-06, 
    7.663642e-06, 7.663636e-06, 7.663628e-06, 7.663693e-06, 7.663696e-06, 
    7.663692e-06, 7.663686e-06, 7.663682e-06, 7.663674e-06, 7.663673e-06, 
    7.663672e-06, 7.663669e-06, 7.663666e-06, 7.663672e-06, 7.663665e-06, 
    7.66369e-06, 7.663677e-06, 7.663697e-06, 7.663691e-06, 7.663687e-06, 
    7.663689e-06, 7.663679e-06, 7.663677e-06, 7.663668e-06, 7.663672e-06, 
    7.663644e-06, 7.663657e-06, 7.663622e-06, 7.663632e-06, 7.663697e-06, 
    7.663693e-06, 7.663683e-06, 7.663688e-06, 7.663673e-06, 7.663671e-06, 
    7.663667e-06, 7.663663e-06, 7.663663e-06, 7.663661e-06, 7.663664e-06, 
    7.663662e-06, 7.663674e-06, 7.663669e-06, 7.663684e-06, 7.663681e-06, 
    7.663682e-06, 7.663684e-06, 7.663678e-06, 7.663672e-06, 7.663672e-06, 
    7.66367e-06, 7.663663e-06, 7.663673e-06, 7.663642e-06, 7.663662e-06, 
    7.663691e-06, 7.663684e-06, 7.663683e-06, 7.663686e-06, 7.663671e-06, 
    7.663676e-06, 7.663662e-06, 7.663665e-06, 7.663659e-06, 7.663662e-06, 
    7.663662e-06, 7.663667e-06, 7.663669e-06, 7.663676e-06, 7.663682e-06, 
    7.663686e-06, 7.663684e-06, 7.66368e-06, 7.663672e-06, 7.663663e-06, 
    7.663665e-06, 7.663659e-06, 7.663675e-06, 7.663668e-06, 7.663671e-06, 
    7.663664e-06, 7.663679e-06, 7.663666e-06, 7.663682e-06, 7.663681e-06, 
    7.663676e-06, 7.663668e-06, 7.663666e-06, 7.663664e-06, 7.663665e-06, 
    7.663671e-06, 7.663672e-06, 7.663676e-06, 7.663678e-06, 7.663681e-06, 
    7.663683e-06, 7.663681e-06, 7.663679e-06, 7.663671e-06, 7.663664e-06, 
    7.663657e-06, 7.663655e-06, 7.663647e-06, 7.663654e-06, 7.663642e-06, 
    7.663652e-06, 7.663636e-06, 7.663665e-06, 7.663652e-06, 7.663676e-06, 
    7.663673e-06, 7.663669e-06, 7.663659e-06, 7.663664e-06, 7.663658e-06, 
    7.663672e-06, 7.66368e-06, 7.663682e-06, 7.663685e-06, 7.663682e-06, 
    7.663682e-06, 7.663678e-06, 7.66368e-06, 7.663671e-06, 7.663675e-06, 
    7.663662e-06, 7.663658e-06, 7.663644e-06, 7.663636e-06, 7.663627e-06, 
    7.663623e-06, 7.663622e-06, 7.663622e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.319314e-14, 5.33372e-14, 5.330921e-14, 5.34253e-14, 5.336093e-14, 
    5.343692e-14, 5.322238e-14, 5.33429e-14, 5.326598e-14, 5.320614e-14, 
    5.365024e-14, 5.343048e-14, 5.387835e-14, 5.373844e-14, 5.408968e-14, 
    5.385656e-14, 5.413665e-14, 5.408301e-14, 5.424451e-14, 5.419827e-14, 
    5.440452e-14, 5.426585e-14, 5.45114e-14, 5.437145e-14, 5.439333e-14, 
    5.426127e-14, 5.347478e-14, 5.362289e-14, 5.346599e-14, 5.348713e-14, 
    5.347765e-14, 5.336225e-14, 5.330402e-14, 5.318215e-14, 5.320429e-14, 
    5.329382e-14, 5.349663e-14, 5.342785e-14, 5.360122e-14, 5.359731e-14, 
    5.379004e-14, 5.370317e-14, 5.402671e-14, 5.393486e-14, 5.42002e-14, 
    5.41335e-14, 5.419706e-14, 5.41778e-14, 5.419731e-14, 5.409948e-14, 
    5.41414e-14, 5.40553e-14, 5.371944e-14, 5.381822e-14, 5.352335e-14, 
    5.334567e-14, 5.322766e-14, 5.314382e-14, 5.315567e-14, 5.317826e-14, 
    5.329434e-14, 5.340344e-14, 5.348651e-14, 5.354204e-14, 5.359674e-14, 
    5.376206e-14, 5.384959e-14, 5.404526e-14, 5.401e-14, 5.406975e-14, 
    5.412687e-14, 5.422265e-14, 5.42069e-14, 5.424907e-14, 5.406821e-14, 
    5.418842e-14, 5.398994e-14, 5.404423e-14, 5.361145e-14, 5.344641e-14, 
    5.337607e-14, 5.331459e-14, 5.316478e-14, 5.326824e-14, 5.322746e-14, 
    5.33245e-14, 5.338609e-14, 5.335564e-14, 5.354356e-14, 5.347052e-14, 
    5.385477e-14, 5.36894e-14, 5.412021e-14, 5.401724e-14, 5.414488e-14, 
    5.407977e-14, 5.41913e-14, 5.409093e-14, 5.426478e-14, 5.430258e-14, 
    5.427674e-14, 5.437603e-14, 5.408536e-14, 5.419704e-14, 5.335478e-14, 
    5.335975e-14, 5.33829e-14, 5.328108e-14, 5.327486e-14, 5.318154e-14, 
    5.32646e-14, 5.329994e-14, 5.338968e-14, 5.34427e-14, 5.34931e-14, 
    5.360385e-14, 5.37274e-14, 5.390003e-14, 5.402392e-14, 5.410691e-14, 
    5.405604e-14, 5.410095e-14, 5.405073e-14, 5.40272e-14, 5.42884e-14, 
    5.414178e-14, 5.436175e-14, 5.434959e-14, 5.425006e-14, 5.435096e-14, 
    5.336323e-14, 5.333465e-14, 5.32353e-14, 5.331305e-14, 5.317138e-14, 
    5.325068e-14, 5.329624e-14, 5.347202e-14, 5.351065e-14, 5.35464e-14, 
    5.361704e-14, 5.370762e-14, 5.386636e-14, 5.400432e-14, 5.41302e-14, 
    5.412098e-14, 5.412423e-14, 5.415231e-14, 5.40827e-14, 5.416374e-14, 
    5.417732e-14, 5.414178e-14, 5.434796e-14, 5.42891e-14, 5.434933e-14, 
    5.431101e-14, 5.334395e-14, 5.339205e-14, 5.336605e-14, 5.341492e-14, 
    5.338048e-14, 5.353351e-14, 5.357935e-14, 5.379372e-14, 5.370583e-14, 
    5.384573e-14, 5.372006e-14, 5.374233e-14, 5.385022e-14, 5.372686e-14, 
    5.399672e-14, 5.381376e-14, 5.41534e-14, 5.397088e-14, 5.416483e-14, 
    5.412965e-14, 5.418791e-14, 5.424005e-14, 5.430564e-14, 5.442653e-14, 
    5.439855e-14, 5.449962e-14, 5.346375e-14, 5.352607e-14, 5.352061e-14, 
    5.358583e-14, 5.363403e-14, 5.373849e-14, 5.390583e-14, 5.384294e-14, 
    5.395841e-14, 5.398157e-14, 5.380615e-14, 5.391385e-14, 5.356779e-14, 
    5.362372e-14, 5.359045e-14, 5.346865e-14, 5.385739e-14, 5.365801e-14, 
    5.402596e-14, 5.391815e-14, 5.423261e-14, 5.407626e-14, 5.438314e-14, 
    5.451403e-14, 5.463725e-14, 5.478092e-14, 5.356011e-14, 5.351777e-14, 
    5.359359e-14, 5.369837e-14, 5.379561e-14, 5.392472e-14, 5.393794e-14, 
    5.396211e-14, 5.402469e-14, 5.407729e-14, 5.396972e-14, 5.409048e-14, 
    5.363663e-14, 5.38747e-14, 5.350173e-14, 5.36141e-14, 5.369221e-14, 
    5.365799e-14, 5.383576e-14, 5.387761e-14, 5.404752e-14, 5.395974e-14, 
    5.448171e-14, 5.425101e-14, 5.489031e-14, 5.471195e-14, 5.350296e-14, 
    5.355997e-14, 5.375815e-14, 5.36639e-14, 5.393336e-14, 5.399959e-14, 
    5.40534e-14, 5.412215e-14, 5.412959e-14, 5.417031e-14, 5.410358e-14, 
    5.416769e-14, 5.3925e-14, 5.403349e-14, 5.373555e-14, 5.380812e-14, 
    5.377475e-14, 5.373812e-14, 5.385114e-14, 5.39714e-14, 5.397402e-14, 
    5.401252e-14, 5.412095e-14, 5.393445e-14, 5.451136e-14, 5.415526e-14, 
    5.362211e-14, 5.373173e-14, 5.374744e-14, 5.370498e-14, 5.399295e-14, 
    5.388867e-14, 5.416932e-14, 5.409353e-14, 5.42177e-14, 5.415601e-14, 
    5.414693e-14, 5.406766e-14, 5.401827e-14, 5.389344e-14, 5.379179e-14, 
    5.371115e-14, 5.372991e-14, 5.381847e-14, 5.397877e-14, 5.413024e-14, 
    5.409706e-14, 5.420827e-14, 5.391383e-14, 5.403733e-14, 5.398961e-14, 
    5.411406e-14, 5.384125e-14, 5.407344e-14, 5.378182e-14, 5.380743e-14, 
    5.38866e-14, 5.404567e-14, 5.408092e-14, 5.411846e-14, 5.409531e-14, 
    5.398284e-14, 5.396443e-14, 5.388469e-14, 5.386264e-14, 5.380185e-14, 
    5.375148e-14, 5.379749e-14, 5.384578e-14, 5.398291e-14, 5.410631e-14, 
    5.424078e-14, 5.427369e-14, 5.443046e-14, 5.430278e-14, 5.451333e-14, 
    5.433424e-14, 5.464416e-14, 5.408696e-14, 5.432907e-14, 5.389022e-14, 
    5.393758e-14, 5.402312e-14, 5.421929e-14, 5.411347e-14, 5.423724e-14, 
    5.396371e-14, 5.38215e-14, 5.378475e-14, 5.371604e-14, 5.378632e-14, 
    5.378061e-14, 5.384782e-14, 5.382623e-14, 5.398746e-14, 5.390088e-14, 
    5.414669e-14, 5.423628e-14, 5.448901e-14, 5.464368e-14, 5.480101e-14, 
    5.487038e-14, 5.489149e-14, 5.490031e-14 ;

 LITTERC =
  5.976207e-05, 5.976193e-05, 5.976195e-05, 5.976183e-05, 5.97619e-05, 
    5.976182e-05, 5.976204e-05, 5.976192e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976183e-05, 5.976138e-05, 5.976152e-05, 5.976116e-05, 
    5.97614e-05, 5.976111e-05, 5.976117e-05, 5.976101e-05, 5.976105e-05, 
    5.976085e-05, 5.976098e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976178e-05, 5.976163e-05, 5.976179e-05, 5.976177e-05, 
    5.976178e-05, 5.97619e-05, 5.976196e-05, 5.976208e-05, 5.976206e-05, 
    5.976197e-05, 5.976176e-05, 5.976183e-05, 5.976166e-05, 5.976166e-05, 
    5.976147e-05, 5.976155e-05, 5.976123e-05, 5.976132e-05, 5.976105e-05, 
    5.976112e-05, 5.976105e-05, 5.976107e-05, 5.976105e-05, 5.976115e-05, 
    5.976111e-05, 5.97612e-05, 5.976154e-05, 5.976144e-05, 5.976174e-05, 
    5.976191e-05, 5.976203e-05, 5.976212e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976177e-05, 5.976172e-05, 5.976166e-05, 
    5.976149e-05, 5.976141e-05, 5.976121e-05, 5.976124e-05, 5.976118e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.9761e-05, 5.976118e-05, 
    5.976106e-05, 5.976126e-05, 5.976121e-05, 5.976165e-05, 5.976181e-05, 
    5.976189e-05, 5.976195e-05, 5.97621e-05, 5.976199e-05, 5.976203e-05, 
    5.976194e-05, 5.976187e-05, 5.976191e-05, 5.976171e-05, 5.976179e-05, 
    5.97614e-05, 5.976157e-05, 5.976113e-05, 5.976123e-05, 5.976111e-05, 
    5.976117e-05, 5.976106e-05, 5.976116e-05, 5.976098e-05, 5.976095e-05, 
    5.976097e-05, 5.976087e-05, 5.976117e-05, 5.976105e-05, 5.976191e-05, 
    5.97619e-05, 5.976188e-05, 5.976198e-05, 5.976199e-05, 5.976208e-05, 
    5.9762e-05, 5.976196e-05, 5.976187e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976153e-05, 5.976135e-05, 5.976123e-05, 5.976114e-05, 
    5.97612e-05, 5.976115e-05, 5.97612e-05, 5.976123e-05, 5.976096e-05, 
    5.976111e-05, 5.976089e-05, 5.97609e-05, 5.9761e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976171e-05, 
    5.976164e-05, 5.976155e-05, 5.976139e-05, 5.976125e-05, 5.976112e-05, 
    5.976113e-05, 5.976113e-05, 5.97611e-05, 5.976117e-05, 5.976109e-05, 
    5.976107e-05, 5.976111e-05, 5.97609e-05, 5.976096e-05, 5.97609e-05, 
    5.976094e-05, 5.976192e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976188e-05, 5.976173e-05, 5.976168e-05, 5.976146e-05, 5.976155e-05, 
    5.976141e-05, 5.976154e-05, 5.976151e-05, 5.976141e-05, 5.976153e-05, 
    5.976126e-05, 5.976144e-05, 5.97611e-05, 5.976128e-05, 5.976109e-05, 
    5.976112e-05, 5.976106e-05, 5.976101e-05, 5.976094e-05, 5.976082e-05, 
    5.976085e-05, 5.976075e-05, 5.97618e-05, 5.976173e-05, 5.976174e-05, 
    5.976167e-05, 5.976162e-05, 5.976152e-05, 5.976135e-05, 5.976141e-05, 
    5.97613e-05, 5.976127e-05, 5.976145e-05, 5.976134e-05, 5.976169e-05, 
    5.976163e-05, 5.976167e-05, 5.976179e-05, 5.97614e-05, 5.97616e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976073e-05, 5.976061e-05, 5.976046e-05, 5.97617e-05, 5.976174e-05, 
    5.976166e-05, 5.976156e-05, 5.976146e-05, 5.976133e-05, 5.976131e-05, 
    5.976129e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976116e-05, 
    5.976162e-05, 5.976138e-05, 5.976176e-05, 5.976165e-05, 5.976157e-05, 
    5.97616e-05, 5.976142e-05, 5.976138e-05, 5.976121e-05, 5.976129e-05, 
    5.976076e-05, 5.9761e-05, 5.976035e-05, 5.976053e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.976159e-05, 5.976132e-05, 5.976125e-05, 
    5.97612e-05, 5.976113e-05, 5.976112e-05, 5.976108e-05, 5.976115e-05, 
    5.976109e-05, 5.976133e-05, 5.976122e-05, 5.976152e-05, 5.976145e-05, 
    5.976148e-05, 5.976152e-05, 5.976141e-05, 5.976128e-05, 5.976128e-05, 
    5.976124e-05, 5.976113e-05, 5.976132e-05, 5.976074e-05, 5.97611e-05, 
    5.976163e-05, 5.976153e-05, 5.976151e-05, 5.976155e-05, 5.976126e-05, 
    5.976137e-05, 5.976108e-05, 5.976116e-05, 5.976103e-05, 5.97611e-05, 
    5.97611e-05, 5.976118e-05, 5.976123e-05, 5.976136e-05, 5.976146e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976127e-05, 5.976112e-05, 
    5.976115e-05, 5.976104e-05, 5.976134e-05, 5.976122e-05, 5.976126e-05, 
    5.976114e-05, 5.976141e-05, 5.976118e-05, 5.976147e-05, 5.976145e-05, 
    5.976137e-05, 5.976121e-05, 5.976117e-05, 5.976113e-05, 5.976116e-05, 
    5.976127e-05, 5.976129e-05, 5.976137e-05, 5.976139e-05, 5.976145e-05, 
    5.97615e-05, 5.976146e-05, 5.976141e-05, 5.976127e-05, 5.976115e-05, 
    5.976101e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976073e-05, 
    5.976091e-05, 5.97606e-05, 5.976117e-05, 5.976092e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976103e-05, 5.976114e-05, 5.976101e-05, 
    5.976129e-05, 5.976143e-05, 5.976147e-05, 5.976154e-05, 5.976147e-05, 
    5.976147e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976135e-05, 
    5.97611e-05, 5.976101e-05, 5.976076e-05, 5.97606e-05, 5.976044e-05, 
    5.976037e-05, 5.976035e-05, 5.976034e-05 ;

 LITTERC_HR =
  8.582233e-13, 8.605457e-13, 8.600946e-13, 8.61966e-13, 8.609284e-13, 
    8.621533e-13, 8.586947e-13, 8.606376e-13, 8.593977e-13, 8.58433e-13, 
    8.655925e-13, 8.620496e-13, 8.692698e-13, 8.670143e-13, 8.726766e-13, 
    8.689185e-13, 8.734338e-13, 8.725691e-13, 8.751727e-13, 8.744272e-13, 
    8.777522e-13, 8.755167e-13, 8.794752e-13, 8.77219e-13, 8.775718e-13, 
    8.754428e-13, 8.627638e-13, 8.651514e-13, 8.62622e-13, 8.629628e-13, 
    8.628101e-13, 8.609495e-13, 8.600109e-13, 8.580462e-13, 8.584032e-13, 
    8.598464e-13, 8.631159e-13, 8.620071e-13, 8.648021e-13, 8.647391e-13, 
    8.678461e-13, 8.664457e-13, 8.716615e-13, 8.701809e-13, 8.744583e-13, 
    8.733831e-13, 8.744077e-13, 8.740972e-13, 8.744117e-13, 8.728347e-13, 
    8.735105e-13, 8.721225e-13, 8.667079e-13, 8.683005e-13, 8.635468e-13, 
    8.606823e-13, 8.587798e-13, 8.574282e-13, 8.576193e-13, 8.579834e-13, 
    8.598548e-13, 8.616137e-13, 8.629528e-13, 8.638481e-13, 8.6473e-13, 
    8.673951e-13, 8.688061e-13, 8.719605e-13, 8.713922e-13, 8.723554e-13, 
    8.732762e-13, 8.748203e-13, 8.745663e-13, 8.752462e-13, 8.723305e-13, 
    8.742684e-13, 8.710687e-13, 8.719439e-13, 8.64967e-13, 8.623064e-13, 
    8.611724e-13, 8.601812e-13, 8.577662e-13, 8.594341e-13, 8.587766e-13, 
    8.60341e-13, 8.613341e-13, 8.60843e-13, 8.638726e-13, 8.626952e-13, 
    8.688898e-13, 8.662237e-13, 8.731688e-13, 8.715089e-13, 8.735666e-13, 
    8.72517e-13, 8.743149e-13, 8.726968e-13, 8.754994e-13, 8.761088e-13, 
    8.756923e-13, 8.772928e-13, 8.726071e-13, 8.744074e-13, 8.608291e-13, 
    8.609092e-13, 8.612826e-13, 8.596411e-13, 8.595408e-13, 8.580363e-13, 
    8.593753e-13, 8.59945e-13, 8.613918e-13, 8.622466e-13, 8.630591e-13, 
    8.648445e-13, 8.668363e-13, 8.696193e-13, 8.716165e-13, 8.729544e-13, 
    8.721343e-13, 8.728583e-13, 8.720488e-13, 8.716694e-13, 8.758803e-13, 
    8.735166e-13, 8.770627e-13, 8.768667e-13, 8.752623e-13, 8.768888e-13, 
    8.609655e-13, 8.605046e-13, 8.58903e-13, 8.601565e-13, 8.578724e-13, 
    8.591509e-13, 8.598855e-13, 8.627192e-13, 8.63342e-13, 8.639184e-13, 
    8.650572e-13, 8.665174e-13, 8.690765e-13, 8.713006e-13, 8.733298e-13, 
    8.731813e-13, 8.732336e-13, 8.736864e-13, 8.725642e-13, 8.738706e-13, 
    8.740895e-13, 8.735166e-13, 8.768404e-13, 8.758914e-13, 8.768625e-13, 
    8.762447e-13, 8.606545e-13, 8.6143e-13, 8.61011e-13, 8.617988e-13, 
    8.612435e-13, 8.637105e-13, 8.644496e-13, 8.679055e-13, 8.664885e-13, 
    8.68744e-13, 8.667179e-13, 8.670769e-13, 8.688164e-13, 8.668277e-13, 
    8.71178e-13, 8.682285e-13, 8.73704e-13, 8.707614e-13, 8.738882e-13, 
    8.733211e-13, 8.742602e-13, 8.751007e-13, 8.761581e-13, 8.78107e-13, 
    8.77656e-13, 8.792853e-13, 8.625859e-13, 8.635906e-13, 8.635026e-13, 
    8.64554e-13, 8.653311e-13, 8.670152e-13, 8.697128e-13, 8.686989e-13, 
    8.705605e-13, 8.709338e-13, 8.681058e-13, 8.698421e-13, 8.642631e-13, 
    8.651649e-13, 8.646285e-13, 8.626649e-13, 8.689319e-13, 8.657175e-13, 
    8.716494e-13, 8.699114e-13, 8.749808e-13, 8.724604e-13, 8.774076e-13, 
    8.795176e-13, 8.81504e-13, 8.8382e-13, 8.641393e-13, 8.634568e-13, 
    8.646792e-13, 8.663683e-13, 8.679359e-13, 8.700174e-13, 8.702305e-13, 
    8.706201e-13, 8.716289e-13, 8.724769e-13, 8.707427e-13, 8.726895e-13, 
    8.65373e-13, 8.692109e-13, 8.631982e-13, 8.650098e-13, 8.66269e-13, 
    8.657173e-13, 8.685831e-13, 8.692578e-13, 8.719969e-13, 8.705819e-13, 
    8.789965e-13, 8.752774e-13, 8.855835e-13, 8.827082e-13, 8.632181e-13, 
    8.641372e-13, 8.673321e-13, 8.658126e-13, 8.701565e-13, 8.712243e-13, 
    8.720918e-13, 8.732001e-13, 8.733201e-13, 8.739765e-13, 8.729007e-13, 
    8.739342e-13, 8.700218e-13, 8.717709e-13, 8.669677e-13, 8.681375e-13, 
    8.675997e-13, 8.670091e-13, 8.688312e-13, 8.707699e-13, 8.708122e-13, 
    8.714328e-13, 8.731807e-13, 8.701742e-13, 8.794746e-13, 8.737338e-13, 
    8.651389e-13, 8.669062e-13, 8.671594e-13, 8.664749e-13, 8.711172e-13, 
    8.694361e-13, 8.739606e-13, 8.727388e-13, 8.747405e-13, 8.73746e-13, 
    8.735996e-13, 8.723216e-13, 8.715254e-13, 8.695131e-13, 8.678743e-13, 
    8.665743e-13, 8.668767e-13, 8.683045e-13, 8.708886e-13, 8.733305e-13, 
    8.727957e-13, 8.745885e-13, 8.698418e-13, 8.718328e-13, 8.710635e-13, 
    8.730696e-13, 8.686718e-13, 8.724148e-13, 8.677136e-13, 8.681264e-13, 
    8.694028e-13, 8.719672e-13, 8.725355e-13, 8.731406e-13, 8.727674e-13, 
    8.709544e-13, 8.706574e-13, 8.69372e-13, 8.690165e-13, 8.680366e-13, 
    8.672246e-13, 8.679663e-13, 8.687447e-13, 8.709555e-13, 8.729448e-13, 
    8.751125e-13, 8.75643e-13, 8.781703e-13, 8.761121e-13, 8.795063e-13, 
    8.766191e-13, 8.816153e-13, 8.726327e-13, 8.765359e-13, 8.694611e-13, 
    8.702247e-13, 8.716036e-13, 8.747661e-13, 8.730603e-13, 8.750555e-13, 
    8.706459e-13, 8.683533e-13, 8.677608e-13, 8.666532e-13, 8.677861e-13, 
    8.67694e-13, 8.687776e-13, 8.684295e-13, 8.710288e-13, 8.69633e-13, 
    8.735957e-13, 8.750399e-13, 8.791143e-13, 8.816076e-13, 8.841439e-13, 
    8.852622e-13, 8.856025e-13, 8.857447e-13 ;

 LITTERC_LOSS =
  1.58942e-12, 1.593722e-12, 1.592886e-12, 1.596352e-12, 1.59443e-12, 
    1.596699e-12, 1.590293e-12, 1.593892e-12, 1.591595e-12, 1.589809e-12, 
    1.603068e-12, 1.596507e-12, 1.609879e-12, 1.605701e-12, 1.616188e-12, 
    1.609228e-12, 1.617591e-12, 1.615989e-12, 1.620811e-12, 1.61943e-12, 
    1.625588e-12, 1.621448e-12, 1.628779e-12, 1.624601e-12, 1.625254e-12, 
    1.621311e-12, 1.59783e-12, 1.602251e-12, 1.597567e-12, 1.598198e-12, 
    1.597915e-12, 1.59447e-12, 1.592731e-12, 1.589092e-12, 1.589754e-12, 
    1.592426e-12, 1.598482e-12, 1.596428e-12, 1.601604e-12, 1.601488e-12, 
    1.607242e-12, 1.604648e-12, 1.614308e-12, 1.611566e-12, 1.619488e-12, 
    1.617497e-12, 1.619394e-12, 1.618819e-12, 1.619402e-12, 1.616481e-12, 
    1.617733e-12, 1.615162e-12, 1.605134e-12, 1.608084e-12, 1.59928e-12, 
    1.593975e-12, 1.590451e-12, 1.587948e-12, 1.588302e-12, 1.588976e-12, 
    1.592442e-12, 1.595699e-12, 1.59818e-12, 1.599838e-12, 1.601471e-12, 
    1.606407e-12, 1.60902e-12, 1.614862e-12, 1.613809e-12, 1.615593e-12, 
    1.617299e-12, 1.620158e-12, 1.619688e-12, 1.620947e-12, 1.615547e-12, 
    1.619136e-12, 1.61321e-12, 1.614831e-12, 1.60191e-12, 1.596983e-12, 
    1.594882e-12, 1.593047e-12, 1.588574e-12, 1.591663e-12, 1.590445e-12, 
    1.593342e-12, 1.595182e-12, 1.594272e-12, 1.599883e-12, 1.597702e-12, 
    1.609175e-12, 1.604237e-12, 1.6171e-12, 1.614026e-12, 1.617837e-12, 
    1.615893e-12, 1.619222e-12, 1.616226e-12, 1.621416e-12, 1.622545e-12, 
    1.621773e-12, 1.624737e-12, 1.616059e-12, 1.619394e-12, 1.594247e-12, 
    1.594395e-12, 1.595086e-12, 1.592046e-12, 1.591861e-12, 1.589074e-12, 
    1.591554e-12, 1.592609e-12, 1.595289e-12, 1.596872e-12, 1.598376e-12, 
    1.601683e-12, 1.605372e-12, 1.610526e-12, 1.614225e-12, 1.616703e-12, 
    1.615184e-12, 1.616525e-12, 1.615025e-12, 1.614323e-12, 1.622121e-12, 
    1.617744e-12, 1.624311e-12, 1.623948e-12, 1.620977e-12, 1.623989e-12, 
    1.594499e-12, 1.593645e-12, 1.590679e-12, 1.593001e-12, 1.588771e-12, 
    1.591138e-12, 1.592499e-12, 1.597747e-12, 1.5989e-12, 1.599968e-12, 
    1.602077e-12, 1.604781e-12, 1.609521e-12, 1.61364e-12, 1.617398e-12, 
    1.617123e-12, 1.61722e-12, 1.618058e-12, 1.61598e-12, 1.618399e-12, 
    1.618805e-12, 1.617744e-12, 1.6239e-12, 1.622142e-12, 1.623941e-12, 
    1.622796e-12, 1.593923e-12, 1.595359e-12, 1.594583e-12, 1.596042e-12, 
    1.595014e-12, 1.599583e-12, 1.600952e-12, 1.607352e-12, 1.604728e-12, 
    1.608905e-12, 1.605153e-12, 1.605817e-12, 1.609039e-12, 1.605356e-12, 
    1.613413e-12, 1.60795e-12, 1.618091e-12, 1.612641e-12, 1.618432e-12, 
    1.617382e-12, 1.619121e-12, 1.620678e-12, 1.622636e-12, 1.626245e-12, 
    1.62541e-12, 1.628428e-12, 1.5975e-12, 1.599361e-12, 1.599198e-12, 
    1.601145e-12, 1.602584e-12, 1.605703e-12, 1.610699e-12, 1.608821e-12, 
    1.612269e-12, 1.612961e-12, 1.607723e-12, 1.610939e-12, 1.600606e-12, 
    1.602276e-12, 1.601283e-12, 1.597646e-12, 1.609253e-12, 1.6033e-12, 
    1.614286e-12, 1.611067e-12, 1.620456e-12, 1.615788e-12, 1.62495e-12, 
    1.628858e-12, 1.632537e-12, 1.636826e-12, 1.600377e-12, 1.599113e-12, 
    1.601377e-12, 1.604505e-12, 1.607408e-12, 1.611263e-12, 1.611658e-12, 
    1.61238e-12, 1.614248e-12, 1.615818e-12, 1.612607e-12, 1.616212e-12, 
    1.602662e-12, 1.60977e-12, 1.598634e-12, 1.601989e-12, 1.604321e-12, 
    1.603299e-12, 1.608607e-12, 1.609857e-12, 1.614929e-12, 1.612309e-12, 
    1.627893e-12, 1.621005e-12, 1.640092e-12, 1.634767e-12, 1.598671e-12, 
    1.600373e-12, 1.60629e-12, 1.603476e-12, 1.611521e-12, 1.613498e-12, 
    1.615105e-12, 1.617158e-12, 1.61738e-12, 1.618596e-12, 1.616603e-12, 
    1.618517e-12, 1.611271e-12, 1.614511e-12, 1.605615e-12, 1.607782e-12, 
    1.606786e-12, 1.605692e-12, 1.609066e-12, 1.612657e-12, 1.612735e-12, 
    1.613885e-12, 1.617122e-12, 1.611554e-12, 1.628778e-12, 1.618146e-12, 
    1.602228e-12, 1.605501e-12, 1.60597e-12, 1.604703e-12, 1.6133e-12, 
    1.610187e-12, 1.618566e-12, 1.616303e-12, 1.620011e-12, 1.618169e-12, 
    1.617898e-12, 1.615531e-12, 1.614056e-12, 1.610329e-12, 1.607294e-12, 
    1.604887e-12, 1.605447e-12, 1.608091e-12, 1.612877e-12, 1.617399e-12, 
    1.616409e-12, 1.619729e-12, 1.610938e-12, 1.614625e-12, 1.613201e-12, 
    1.616916e-12, 1.608771e-12, 1.615703e-12, 1.606997e-12, 1.607761e-12, 
    1.610125e-12, 1.614874e-12, 1.615927e-12, 1.617048e-12, 1.616356e-12, 
    1.612999e-12, 1.612449e-12, 1.610068e-12, 1.60941e-12, 1.607595e-12, 
    1.606091e-12, 1.607465e-12, 1.608906e-12, 1.613001e-12, 1.616685e-12, 
    1.6207e-12, 1.621682e-12, 1.626363e-12, 1.622551e-12, 1.628837e-12, 
    1.62349e-12, 1.632743e-12, 1.616107e-12, 1.623336e-12, 1.610233e-12, 
    1.611647e-12, 1.614201e-12, 1.620058e-12, 1.616899e-12, 1.620594e-12, 
    1.612427e-12, 1.608181e-12, 1.607084e-12, 1.605033e-12, 1.607131e-12, 
    1.60696e-12, 1.608967e-12, 1.608323e-12, 1.613136e-12, 1.610551e-12, 
    1.61789e-12, 1.620565e-12, 1.628111e-12, 1.632729e-12, 1.637426e-12, 
    1.639497e-12, 1.640127e-12, 1.640391e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  3.916361e-18, 3.914928e-18, 3.915199e-18, 3.914059e-18, 3.914681e-18, 
    3.913942e-18, 3.916058e-18, 3.914881e-18, 3.915625e-18, 3.916215e-18, 
    3.911885e-18, 3.914005e-18, 3.909574e-18, 3.910941e-18, 3.907476e-18, 
    3.909802e-18, 3.907003e-18, 3.907516e-18, 3.905907e-18, 3.906365e-18, 
    3.904367e-18, 3.905694e-18, 3.90329e-18, 3.904669e-18, 3.904464e-18, 
    3.905743e-18, 3.913552e-18, 3.912157e-18, 3.91364e-18, 3.91344e-18, 
    3.913524e-18, 3.914678e-18, 3.915278e-18, 3.916452e-18, 3.916234e-18, 
    3.915361e-18, 3.913349e-18, 3.914014e-18, 3.912288e-18, 3.912326e-18, 
    3.910426e-18, 3.911282e-18, 3.908075e-18, 3.908979e-18, 3.906346e-18, 
    3.907011e-18, 3.906382e-18, 3.906569e-18, 3.906379e-18, 3.907354e-18, 
    3.906938e-18, 3.907787e-18, 3.911127e-18, 3.910153e-18, 3.913076e-18, 
    3.914879e-18, 3.916012e-18, 3.916836e-18, 3.91672e-18, 3.916503e-18, 
    3.915356e-18, 3.914257e-18, 3.913427e-18, 3.912877e-18, 3.912331e-18, 
    3.910753e-18, 3.909859e-18, 3.907905e-18, 3.908234e-18, 3.907659e-18, 
    3.907076e-18, 3.906131e-18, 3.906283e-18, 3.905872e-18, 3.907657e-18, 
    3.906479e-18, 3.908428e-18, 3.907897e-18, 3.912276e-18, 3.91383e-18, 
    3.914571e-18, 3.91515e-18, 3.916632e-18, 3.915614e-18, 3.916017e-18, 
    3.915038e-18, 3.91443e-18, 3.914727e-18, 3.912862e-18, 3.91359e-18, 
    3.909806e-18, 3.911433e-18, 3.907145e-18, 3.908165e-18, 3.906897e-18, 
    3.907539e-18, 3.906446e-18, 3.907429e-18, 3.905712e-18, 3.905348e-18, 
    3.905599e-18, 3.904608e-18, 3.907486e-18, 3.906391e-18, 3.914739e-18, 
    3.914692e-18, 3.914458e-18, 3.915488e-18, 3.915546e-18, 3.916463e-18, 
    3.915639e-18, 3.915295e-18, 3.914387e-18, 3.913868e-18, 3.913368e-18, 
    3.91227e-18, 3.91106e-18, 3.909345e-18, 3.9081e-18, 3.90727e-18, 
    3.907773e-18, 3.90733e-18, 3.907829e-18, 3.908058e-18, 3.905491e-18, 
    3.906939e-18, 3.90475e-18, 3.904868e-18, 3.905865e-18, 3.904855e-18, 
    3.914657e-18, 3.914935e-18, 3.915933e-18, 3.915152e-18, 3.916562e-18, 
    3.915784e-18, 3.915343e-18, 3.913595e-18, 3.913189e-18, 3.912842e-18, 
    3.912135e-18, 3.911239e-18, 3.909676e-18, 3.908303e-18, 3.907039e-18, 
    3.90713e-18, 3.907098e-18, 3.906826e-18, 3.907514e-18, 3.906712e-18, 
    3.906586e-18, 3.906929e-18, 3.904884e-18, 3.905467e-18, 3.904871e-18, 
    3.905247e-18, 3.914842e-18, 3.914369e-18, 3.914626e-18, 3.914148e-18, 
    3.914492e-18, 3.91299e-18, 3.91254e-18, 3.910412e-18, 3.911262e-18, 
    3.909885e-18, 3.911115e-18, 3.910902e-18, 3.909878e-18, 3.911042e-18, 
    3.908397e-18, 3.910224e-18, 3.906815e-18, 3.908673e-18, 3.906701e-18, 
    3.907045e-18, 3.906466e-18, 3.905959e-18, 3.905304e-18, 3.904124e-18, 
    3.904393e-18, 3.903393e-18, 3.913656e-18, 3.913052e-18, 3.913088e-18, 
    3.912444e-18, 3.911972e-18, 3.910929e-18, 3.909277e-18, 3.909892e-18, 
    3.908744e-18, 3.90852e-18, 3.910254e-18, 3.909205e-18, 3.912635e-18, 
    3.912098e-18, 3.912405e-18, 3.913619e-18, 3.909774e-18, 3.911755e-18, 
    3.908083e-18, 3.90915e-18, 3.906034e-18, 3.9076e-18, 3.904546e-18, 
    3.903288e-18, 3.902026e-18, 3.900645e-18, 3.912704e-18, 3.913116e-18, 
    3.912363e-18, 3.911354e-18, 3.910369e-18, 3.909088e-18, 3.908948e-18, 
    3.908714e-18, 3.908085e-18, 3.907565e-18, 3.908656e-18, 3.907433e-18, 
    3.912008e-18, 3.909594e-18, 3.913288e-18, 3.912197e-18, 3.911405e-18, 
    3.911735e-18, 3.909958e-18, 3.909546e-18, 3.907878e-18, 3.90873e-18, 
    3.903613e-18, 3.905876e-18, 3.89954e-18, 3.901317e-18, 3.913264e-18, 
    3.912697e-18, 3.910751e-18, 3.911674e-18, 3.908994e-18, 3.908343e-18, 
    3.907799e-18, 3.907133e-18, 3.907048e-18, 3.906651e-18, 3.907303e-18, 
    3.90667e-18, 3.909086e-18, 3.908003e-18, 3.910953e-18, 3.910244e-18, 
    3.910564e-18, 3.910928e-18, 3.909807e-18, 3.908643e-18, 3.908591e-18, 
    3.908222e-18, 3.907234e-18, 3.908982e-18, 3.903372e-18, 3.90688e-18, 
    3.912081e-18, 3.911029e-18, 3.910844e-18, 3.911258e-18, 3.908409e-18, 
    3.909444e-18, 3.906657e-18, 3.907403e-18, 3.906173e-18, 3.906786e-18, 
    3.906878e-18, 3.90766e-18, 3.908155e-18, 3.909402e-18, 3.910409e-18, 
    3.911194e-18, 3.91101e-18, 3.910146e-18, 3.908565e-18, 3.907053e-18, 
    3.907387e-18, 3.906267e-18, 3.909189e-18, 3.907976e-18, 3.908454e-18, 
    3.907205e-18, 3.909914e-18, 3.90769e-18, 3.910493e-18, 3.910242e-18, 
    3.909464e-18, 3.907913e-18, 3.907529e-18, 3.907169e-18, 3.907385e-18, 
    3.90852e-18, 3.908694e-18, 3.909476e-18, 3.909706e-18, 3.910295e-18, 
    3.910795e-18, 3.910345e-18, 3.909878e-18, 3.908509e-18, 3.907291e-18, 
    3.905956e-18, 3.905619e-18, 3.904131e-18, 3.90538e-18, 3.903358e-18, 
    3.905133e-18, 3.902033e-18, 3.90752e-18, 3.905131e-18, 3.909419e-18, 
    3.90895e-18, 3.90813e-18, 3.906195e-18, 3.90721e-18, 3.906009e-18, 
    3.908698e-18, 3.91013e-18, 3.910467e-18, 3.911151e-18, 3.910451e-18, 
    3.910507e-18, 3.909839e-18, 3.910052e-18, 3.908463e-18, 3.909315e-18, 
    3.906888e-18, 3.906012e-18, 3.903507e-18, 3.901993e-18, 3.900409e-18, 
    3.899725e-18, 3.899515e-18, 3.899428e-18 ;

 MEG_acetic_acid =
  5.874542e-19, 5.872391e-19, 5.872799e-19, 5.871088e-19, 5.872021e-19, 
    5.870913e-19, 5.874087e-19, 5.872322e-19, 5.873438e-19, 5.874323e-19, 
    5.867827e-19, 5.871007e-19, 5.864361e-19, 5.866411e-19, 5.861214e-19, 
    5.864703e-19, 5.860504e-19, 5.861273e-19, 5.85886e-19, 5.859548e-19, 
    5.85655e-19, 5.858541e-19, 5.854934e-19, 5.857004e-19, 5.856696e-19, 
    5.858614e-19, 5.870327e-19, 5.868235e-19, 5.87046e-19, 5.87016e-19, 
    5.870286e-19, 5.872017e-19, 5.872917e-19, 5.874678e-19, 5.874351e-19, 
    5.873041e-19, 5.870024e-19, 5.87102e-19, 5.868431e-19, 5.868488e-19, 
    5.865639e-19, 5.866923e-19, 5.862112e-19, 5.863469e-19, 5.859519e-19, 
    5.860517e-19, 5.859572e-19, 5.859853e-19, 5.859569e-19, 5.861031e-19, 
    5.860407e-19, 5.86168e-19, 5.866691e-19, 5.86523e-19, 5.869614e-19, 
    5.872319e-19, 5.874017e-19, 5.875255e-19, 5.87508e-19, 5.874755e-19, 
    5.873035e-19, 5.871385e-19, 5.87014e-19, 5.869315e-19, 5.868497e-19, 
    5.866129e-19, 5.864788e-19, 5.861858e-19, 5.862351e-19, 5.861488e-19, 
    5.860614e-19, 5.859196e-19, 5.859424e-19, 5.858808e-19, 5.861486e-19, 
    5.859718e-19, 5.862642e-19, 5.861845e-19, 5.868413e-19, 5.870745e-19, 
    5.871857e-19, 5.872725e-19, 5.874948e-19, 5.873421e-19, 5.874026e-19, 
    5.872557e-19, 5.871644e-19, 5.87209e-19, 5.869293e-19, 5.870384e-19, 
    5.86471e-19, 5.86715e-19, 5.860716e-19, 5.862247e-19, 5.860345e-19, 
    5.861308e-19, 5.859668e-19, 5.861143e-19, 5.858567e-19, 5.858022e-19, 
    5.858398e-19, 5.856911e-19, 5.861229e-19, 5.859586e-19, 5.872109e-19, 
    5.872037e-19, 5.871687e-19, 5.873232e-19, 5.873319e-19, 5.874694e-19, 
    5.873457e-19, 5.872942e-19, 5.871581e-19, 5.870802e-19, 5.870053e-19, 
    5.868405e-19, 5.86659e-19, 5.864018e-19, 5.862149e-19, 5.860906e-19, 
    5.861659e-19, 5.860995e-19, 5.861743e-19, 5.862087e-19, 5.858236e-19, 
    5.860408e-19, 5.857125e-19, 5.857302e-19, 5.858798e-19, 5.857281e-19, 
    5.871985e-19, 5.872402e-19, 5.873898e-19, 5.872727e-19, 5.874842e-19, 
    5.873676e-19, 5.873015e-19, 5.870392e-19, 5.869783e-19, 5.869262e-19, 
    5.868201e-19, 5.866859e-19, 5.864514e-19, 5.862455e-19, 5.860558e-19, 
    5.860695e-19, 5.860648e-19, 5.860239e-19, 5.861271e-19, 5.860068e-19, 
    5.859879e-19, 5.860393e-19, 5.857326e-19, 5.8582e-19, 5.857306e-19, 
    5.857871e-19, 5.872263e-19, 5.871554e-19, 5.871939e-19, 5.871222e-19, 
    5.871738e-19, 5.869484e-19, 5.868809e-19, 5.865618e-19, 5.866892e-19, 
    5.864827e-19, 5.866671e-19, 5.866352e-19, 5.864818e-19, 5.866563e-19, 
    5.862595e-19, 5.865335e-19, 5.860223e-19, 5.86301e-19, 5.860051e-19, 
    5.860566e-19, 5.859699e-19, 5.858938e-19, 5.857956e-19, 5.856186e-19, 
    5.85659e-19, 5.855088e-19, 5.870484e-19, 5.869578e-19, 5.869632e-19, 
    5.868667e-19, 5.867958e-19, 5.866392e-19, 5.863915e-19, 5.864838e-19, 
    5.863116e-19, 5.86278e-19, 5.86538e-19, 5.863807e-19, 5.868952e-19, 
    5.868147e-19, 5.868607e-19, 5.870427e-19, 5.864661e-19, 5.867633e-19, 
    5.862124e-19, 5.863725e-19, 5.859051e-19, 5.861399e-19, 5.856818e-19, 
    5.854931e-19, 5.853039e-19, 5.850968e-19, 5.869056e-19, 5.869674e-19, 
    5.868544e-19, 5.86703e-19, 5.865553e-19, 5.863633e-19, 5.863422e-19, 
    5.86307e-19, 5.862127e-19, 5.861348e-19, 5.862984e-19, 5.86115e-19, 
    5.868012e-19, 5.864392e-19, 5.869932e-19, 5.868296e-19, 5.867108e-19, 
    5.867603e-19, 5.864936e-19, 5.864318e-19, 5.861816e-19, 5.863094e-19, 
    5.85542e-19, 5.858814e-19, 5.849309e-19, 5.851976e-19, 5.869896e-19, 
    5.869045e-19, 5.866127e-19, 5.867511e-19, 5.86349e-19, 5.862514e-19, 
    5.861698e-19, 5.860698e-19, 5.860572e-19, 5.859976e-19, 5.860955e-19, 
    5.860005e-19, 5.863628e-19, 5.862004e-19, 5.866429e-19, 5.865366e-19, 
    5.865846e-19, 5.866392e-19, 5.864711e-19, 5.862965e-19, 5.862886e-19, 
    5.862333e-19, 5.860851e-19, 5.863473e-19, 5.855058e-19, 5.86032e-19, 
    5.868121e-19, 5.866543e-19, 5.866266e-19, 5.866887e-19, 5.862614e-19, 
    5.864166e-19, 5.859985e-19, 5.861105e-19, 5.85926e-19, 5.86018e-19, 
    5.860317e-19, 5.86149e-19, 5.862233e-19, 5.864102e-19, 5.865613e-19, 
    5.866791e-19, 5.866514e-19, 5.865219e-19, 5.862848e-19, 5.860579e-19, 
    5.861081e-19, 5.8594e-19, 5.863783e-19, 5.861964e-19, 5.862681e-19, 
    5.860807e-19, 5.864871e-19, 5.861535e-19, 5.86574e-19, 5.865362e-19, 
    5.864196e-19, 5.861869e-19, 5.861293e-19, 5.860754e-19, 5.861078e-19, 
    5.86278e-19, 5.863041e-19, 5.864214e-19, 5.864559e-19, 5.865442e-19, 
    5.866192e-19, 5.865517e-19, 5.864816e-19, 5.862763e-19, 5.860936e-19, 
    5.858934e-19, 5.858428e-19, 5.856196e-19, 5.858069e-19, 5.855037e-19, 
    5.8577e-19, 5.85305e-19, 5.86128e-19, 5.857696e-19, 5.864129e-19, 
    5.863424e-19, 5.862195e-19, 5.859292e-19, 5.860815e-19, 5.859014e-19, 
    5.863048e-19, 5.865195e-19, 5.8657e-19, 5.866727e-19, 5.865676e-19, 
    5.86576e-19, 5.864758e-19, 5.865078e-19, 5.862694e-19, 5.863972e-19, 
    5.860332e-19, 5.859017e-19, 5.855261e-19, 5.852988e-19, 5.850613e-19, 
    5.849588e-19, 5.849272e-19, 5.849142e-19 ;

 MEG_acetone =
  1.220792e-16, 1.22056e-16, 1.220604e-16, 1.22042e-16, 1.22052e-16, 
    1.220401e-16, 1.220743e-16, 1.220553e-16, 1.220673e-16, 1.220769e-16, 
    1.220068e-16, 1.220411e-16, 1.219694e-16, 1.219916e-16, 1.219355e-16, 
    1.219731e-16, 1.219279e-16, 1.219362e-16, 1.219102e-16, 1.219176e-16, 
    1.218853e-16, 1.219068e-16, 1.218679e-16, 1.218902e-16, 1.218869e-16, 
    1.219075e-16, 1.220338e-16, 1.220112e-16, 1.220352e-16, 1.22032e-16, 
    1.220333e-16, 1.22052e-16, 1.220617e-16, 1.220807e-16, 1.220772e-16, 
    1.22063e-16, 1.220305e-16, 1.220412e-16, 1.220133e-16, 1.220139e-16, 
    1.219832e-16, 1.219971e-16, 1.219452e-16, 1.219598e-16, 1.219173e-16, 
    1.21928e-16, 1.219178e-16, 1.219209e-16, 1.219178e-16, 1.219335e-16, 
    1.219268e-16, 1.219406e-16, 1.219946e-16, 1.219788e-16, 1.220261e-16, 
    1.220552e-16, 1.220736e-16, 1.220869e-16, 1.22085e-16, 1.220815e-16, 
    1.22063e-16, 1.220452e-16, 1.220318e-16, 1.220229e-16, 1.22014e-16, 
    1.219885e-16, 1.219741e-16, 1.219425e-16, 1.219478e-16, 1.219385e-16, 
    1.219291e-16, 1.219138e-16, 1.219163e-16, 1.219096e-16, 1.219385e-16, 
    1.219194e-16, 1.219509e-16, 1.219423e-16, 1.220131e-16, 1.220383e-16, 
    1.220503e-16, 1.220596e-16, 1.220836e-16, 1.220671e-16, 1.220737e-16, 
    1.220578e-16, 1.22048e-16, 1.220528e-16, 1.220226e-16, 1.220344e-16, 
    1.219732e-16, 1.219995e-16, 1.219302e-16, 1.219467e-16, 1.219262e-16, 
    1.219365e-16, 1.219189e-16, 1.219348e-16, 1.21907e-16, 1.219012e-16, 
    1.219052e-16, 1.218892e-16, 1.219357e-16, 1.21918e-16, 1.22053e-16, 
    1.220522e-16, 1.220484e-16, 1.220651e-16, 1.22066e-16, 1.220809e-16, 
    1.220675e-16, 1.22062e-16, 1.220473e-16, 1.220389e-16, 1.220308e-16, 
    1.22013e-16, 1.219935e-16, 1.219657e-16, 1.219456e-16, 1.219322e-16, 
    1.219403e-16, 1.219332e-16, 1.219412e-16, 1.219449e-16, 1.219035e-16, 
    1.219268e-16, 1.218915e-16, 1.218934e-16, 1.219095e-16, 1.218932e-16, 
    1.220517e-16, 1.220562e-16, 1.220723e-16, 1.220597e-16, 1.220825e-16, 
    1.220699e-16, 1.220628e-16, 1.220345e-16, 1.220279e-16, 1.220223e-16, 
    1.220108e-16, 1.219964e-16, 1.219711e-16, 1.219489e-16, 1.219285e-16, 
    1.219299e-16, 1.219294e-16, 1.21925e-16, 1.219361e-16, 1.219232e-16, 
    1.219211e-16, 1.219267e-16, 1.218937e-16, 1.219031e-16, 1.218935e-16, 
    1.218995e-16, 1.220546e-16, 1.22047e-16, 1.220511e-16, 1.220434e-16, 
    1.22049e-16, 1.220247e-16, 1.220174e-16, 1.21983e-16, 1.219967e-16, 
    1.219745e-16, 1.219944e-16, 1.219909e-16, 1.219744e-16, 1.219932e-16, 
    1.219504e-16, 1.219799e-16, 1.219248e-16, 1.219549e-16, 1.21923e-16, 
    1.219286e-16, 1.219192e-16, 1.21911e-16, 1.219005e-16, 1.218814e-16, 
    1.218858e-16, 1.218696e-16, 1.220355e-16, 1.220257e-16, 1.220263e-16, 
    1.220159e-16, 1.220082e-16, 1.219914e-16, 1.219646e-16, 1.219746e-16, 
    1.21956e-16, 1.219524e-16, 1.219804e-16, 1.219635e-16, 1.220189e-16, 
    1.220103e-16, 1.220152e-16, 1.220349e-16, 1.219727e-16, 1.220047e-16, 
    1.219453e-16, 1.219626e-16, 1.219122e-16, 1.219375e-16, 1.218882e-16, 
    1.218679e-16, 1.218476e-16, 1.218253e-16, 1.220201e-16, 1.220267e-16, 
    1.220145e-16, 1.219982e-16, 1.219823e-16, 1.219616e-16, 1.219593e-16, 
    1.219555e-16, 1.219454e-16, 1.21937e-16, 1.219546e-16, 1.219348e-16, 
    1.220088e-16, 1.219698e-16, 1.220295e-16, 1.220119e-16, 1.219991e-16, 
    1.220044e-16, 1.219757e-16, 1.21969e-16, 1.21942e-16, 1.219558e-16, 
    1.218732e-16, 1.219097e-16, 1.218075e-16, 1.218361e-16, 1.220291e-16, 
    1.2202e-16, 1.219885e-16, 1.220034e-16, 1.219601e-16, 1.219496e-16, 
    1.219407e-16, 1.2193e-16, 1.219286e-16, 1.219222e-16, 1.219327e-16, 
    1.219225e-16, 1.219615e-16, 1.21944e-16, 1.219917e-16, 1.219803e-16, 
    1.219855e-16, 1.219914e-16, 1.219732e-16, 1.219544e-16, 1.219536e-16, 
    1.219476e-16, 1.219316e-16, 1.219599e-16, 1.218693e-16, 1.219259e-16, 
    1.2201e-16, 1.21993e-16, 1.2199e-16, 1.219967e-16, 1.219506e-16, 
    1.219673e-16, 1.219223e-16, 1.219343e-16, 1.219145e-16, 1.219244e-16, 
    1.219259e-16, 1.219385e-16, 1.219465e-16, 1.219667e-16, 1.219829e-16, 
    1.219957e-16, 1.219927e-16, 1.219787e-16, 1.219531e-16, 1.219287e-16, 
    1.219341e-16, 1.21916e-16, 1.219632e-16, 1.219436e-16, 1.219513e-16, 
    1.219311e-16, 1.219749e-16, 1.21939e-16, 1.219843e-16, 1.219802e-16, 
    1.219677e-16, 1.219426e-16, 1.219364e-16, 1.219306e-16, 1.219341e-16, 
    1.219524e-16, 1.219552e-16, 1.219679e-16, 1.219716e-16, 1.219811e-16, 
    1.219892e-16, 1.219819e-16, 1.219744e-16, 1.219522e-16, 1.219325e-16, 
    1.21911e-16, 1.219055e-16, 1.218815e-16, 1.219017e-16, 1.21869e-16, 
    1.218977e-16, 1.218477e-16, 1.219362e-16, 1.218976e-16, 1.219669e-16, 
    1.219594e-16, 1.219461e-16, 1.219148e-16, 1.219312e-16, 1.219118e-16, 
    1.219553e-16, 1.219784e-16, 1.219839e-16, 1.21995e-16, 1.219836e-16, 
    1.219845e-16, 1.219737e-16, 1.219772e-16, 1.219515e-16, 1.219653e-16, 
    1.21926e-16, 1.219119e-16, 1.218715e-16, 1.21847e-16, 1.218215e-16, 
    1.218105e-16, 1.218071e-16, 1.218057e-16 ;

 MEG_carene_3 =
  4.842127e-17, 4.84116e-17, 4.841343e-17, 4.840574e-17, 4.840993e-17, 
    4.840495e-17, 4.841923e-17, 4.841128e-17, 4.84163e-17, 4.842029e-17, 
    4.839107e-17, 4.840537e-17, 4.837549e-17, 4.838471e-17, 4.836135e-17, 
    4.837703e-17, 4.835816e-17, 4.836161e-17, 4.835078e-17, 4.835387e-17, 
    4.834041e-17, 4.834935e-17, 4.833316e-17, 4.834245e-17, 4.834106e-17, 
    4.834967e-17, 4.840231e-17, 4.83929e-17, 4.840291e-17, 4.840156e-17, 
    4.840213e-17, 4.840991e-17, 4.841396e-17, 4.842188e-17, 4.842041e-17, 
    4.841452e-17, 4.840095e-17, 4.840543e-17, 4.839379e-17, 4.839405e-17, 
    4.838124e-17, 4.838702e-17, 4.836538e-17, 4.837148e-17, 4.835374e-17, 
    4.835822e-17, 4.835398e-17, 4.835524e-17, 4.835396e-17, 4.836053e-17, 
    4.835772e-17, 4.836344e-17, 4.838597e-17, 4.83794e-17, 4.839911e-17, 
    4.841126e-17, 4.841891e-17, 4.842448e-17, 4.842369e-17, 4.842223e-17, 
    4.841449e-17, 4.840707e-17, 4.840147e-17, 4.839777e-17, 4.839409e-17, 
    4.838344e-17, 4.837741e-17, 4.836424e-17, 4.836646e-17, 4.836258e-17, 
    4.835866e-17, 4.835229e-17, 4.835331e-17, 4.835054e-17, 4.836257e-17, 
    4.835463e-17, 4.836777e-17, 4.836419e-17, 4.839371e-17, 4.840419e-17, 
    4.840919e-17, 4.84131e-17, 4.84231e-17, 4.841623e-17, 4.841895e-17, 
    4.841234e-17, 4.840824e-17, 4.841024e-17, 4.839766e-17, 4.840257e-17, 
    4.837706e-17, 4.838803e-17, 4.835911e-17, 4.836599e-17, 4.835745e-17, 
    4.836177e-17, 4.835441e-17, 4.836103e-17, 4.834946e-17, 4.834702e-17, 
    4.83487e-17, 4.834203e-17, 4.836142e-17, 4.835404e-17, 4.841033e-17, 
    4.841e-17, 4.840843e-17, 4.841537e-17, 4.841577e-17, 4.842196e-17, 
    4.841639e-17, 4.841407e-17, 4.840795e-17, 4.840445e-17, 4.840108e-17, 
    4.839368e-17, 4.838552e-17, 4.837395e-17, 4.836555e-17, 4.835996e-17, 
    4.836335e-17, 4.836036e-17, 4.836372e-17, 4.836527e-17, 4.834798e-17, 
    4.835773e-17, 4.834299e-17, 4.834378e-17, 4.83505e-17, 4.834369e-17, 
    4.840977e-17, 4.841165e-17, 4.841838e-17, 4.841311e-17, 4.842262e-17, 
    4.841737e-17, 4.84144e-17, 4.840261e-17, 4.839987e-17, 4.839753e-17, 
    4.839276e-17, 4.838672e-17, 4.837618e-17, 4.836692e-17, 4.83584e-17, 
    4.835902e-17, 4.835881e-17, 4.835697e-17, 4.83616e-17, 4.83562e-17, 
    4.835535e-17, 4.835766e-17, 4.83439e-17, 4.834781e-17, 4.83438e-17, 
    4.834634e-17, 4.841102e-17, 4.840783e-17, 4.840956e-17, 4.840634e-17, 
    4.840866e-17, 4.839853e-17, 4.839549e-17, 4.838115e-17, 4.838688e-17, 
    4.837759e-17, 4.838588e-17, 4.838445e-17, 4.837754e-17, 4.838539e-17, 
    4.836756e-17, 4.837987e-17, 4.83569e-17, 4.836942e-17, 4.835612e-17, 
    4.835844e-17, 4.835455e-17, 4.835113e-17, 4.834672e-17, 4.833878e-17, 
    4.834059e-17, 4.833385e-17, 4.840302e-17, 4.839895e-17, 4.839919e-17, 
    4.839485e-17, 4.839166e-17, 4.838463e-17, 4.837349e-17, 4.837764e-17, 
    4.83699e-17, 4.836839e-17, 4.838008e-17, 4.837301e-17, 4.839613e-17, 
    4.839251e-17, 4.839458e-17, 4.840276e-17, 4.837684e-17, 4.83902e-17, 
    4.836544e-17, 4.837264e-17, 4.835164e-17, 4.836218e-17, 4.834162e-17, 
    4.833315e-17, 4.832466e-17, 4.831538e-17, 4.83966e-17, 4.839938e-17, 
    4.83943e-17, 4.838749e-17, 4.838085e-17, 4.837222e-17, 4.837127e-17, 
    4.836969e-17, 4.836545e-17, 4.836195e-17, 4.83693e-17, 4.836106e-17, 
    4.83919e-17, 4.837563e-17, 4.840053e-17, 4.839318e-17, 4.838784e-17, 
    4.839007e-17, 4.837808e-17, 4.83753e-17, 4.836406e-17, 4.83698e-17, 
    4.833534e-17, 4.835057e-17, 4.830795e-17, 4.83199e-17, 4.840038e-17, 
    4.839655e-17, 4.838343e-17, 4.838965e-17, 4.837158e-17, 4.83672e-17, 
    4.836352e-17, 4.835903e-17, 4.835846e-17, 4.835579e-17, 4.836018e-17, 
    4.835592e-17, 4.83722e-17, 4.83649e-17, 4.838479e-17, 4.838001e-17, 
    4.838217e-17, 4.838463e-17, 4.837707e-17, 4.836922e-17, 4.836886e-17, 
    4.836638e-17, 4.835971e-17, 4.83715e-17, 4.833371e-17, 4.835733e-17, 
    4.83924e-17, 4.83853e-17, 4.838406e-17, 4.838685e-17, 4.836764e-17, 
    4.837462e-17, 4.835583e-17, 4.836086e-17, 4.835257e-17, 4.83567e-17, 
    4.835732e-17, 4.836259e-17, 4.836593e-17, 4.837433e-17, 4.838112e-17, 
    4.838642e-17, 4.838517e-17, 4.837935e-17, 4.836869e-17, 4.83585e-17, 
    4.836075e-17, 4.83532e-17, 4.83729e-17, 4.836472e-17, 4.836794e-17, 
    4.835952e-17, 4.837779e-17, 4.836279e-17, 4.838169e-17, 4.837999e-17, 
    4.837475e-17, 4.836429e-17, 4.83617e-17, 4.835928e-17, 4.836074e-17, 
    4.836839e-17, 4.836956e-17, 4.837484e-17, 4.837638e-17, 4.838035e-17, 
    4.838373e-17, 4.838069e-17, 4.837754e-17, 4.836831e-17, 4.83601e-17, 
    4.835111e-17, 4.834884e-17, 4.833882e-17, 4.834723e-17, 4.833362e-17, 
    4.834556e-17, 4.832471e-17, 4.836164e-17, 4.834555e-17, 4.837445e-17, 
    4.837129e-17, 4.836575e-17, 4.835272e-17, 4.835956e-17, 4.835147e-17, 
    4.836959e-17, 4.837924e-17, 4.838151e-17, 4.838613e-17, 4.838141e-17, 
    4.838178e-17, 4.837728e-17, 4.837871e-17, 4.8368e-17, 4.837374e-17, 
    4.835739e-17, 4.835148e-17, 4.833462e-17, 4.832444e-17, 4.83138e-17, 
    4.83092e-17, 4.830779e-17, 4.830721e-17 ;

 MEG_ethanol =
  3.916361e-18, 3.914928e-18, 3.915199e-18, 3.914059e-18, 3.914681e-18, 
    3.913942e-18, 3.916058e-18, 3.914881e-18, 3.915625e-18, 3.916215e-18, 
    3.911885e-18, 3.914005e-18, 3.909574e-18, 3.910941e-18, 3.907476e-18, 
    3.909802e-18, 3.907003e-18, 3.907516e-18, 3.905907e-18, 3.906365e-18, 
    3.904367e-18, 3.905694e-18, 3.90329e-18, 3.904669e-18, 3.904464e-18, 
    3.905743e-18, 3.913552e-18, 3.912157e-18, 3.91364e-18, 3.91344e-18, 
    3.913524e-18, 3.914678e-18, 3.915278e-18, 3.916452e-18, 3.916234e-18, 
    3.915361e-18, 3.913349e-18, 3.914014e-18, 3.912288e-18, 3.912326e-18, 
    3.910426e-18, 3.911282e-18, 3.908075e-18, 3.908979e-18, 3.906346e-18, 
    3.907011e-18, 3.906382e-18, 3.906569e-18, 3.906379e-18, 3.907354e-18, 
    3.906938e-18, 3.907787e-18, 3.911127e-18, 3.910153e-18, 3.913076e-18, 
    3.914879e-18, 3.916012e-18, 3.916836e-18, 3.91672e-18, 3.916503e-18, 
    3.915356e-18, 3.914257e-18, 3.913427e-18, 3.912877e-18, 3.912331e-18, 
    3.910753e-18, 3.909859e-18, 3.907905e-18, 3.908234e-18, 3.907659e-18, 
    3.907076e-18, 3.906131e-18, 3.906283e-18, 3.905872e-18, 3.907657e-18, 
    3.906479e-18, 3.908428e-18, 3.907897e-18, 3.912276e-18, 3.91383e-18, 
    3.914571e-18, 3.91515e-18, 3.916632e-18, 3.915614e-18, 3.916017e-18, 
    3.915038e-18, 3.91443e-18, 3.914727e-18, 3.912862e-18, 3.91359e-18, 
    3.909806e-18, 3.911433e-18, 3.907145e-18, 3.908165e-18, 3.906897e-18, 
    3.907539e-18, 3.906446e-18, 3.907429e-18, 3.905712e-18, 3.905348e-18, 
    3.905599e-18, 3.904608e-18, 3.907486e-18, 3.906391e-18, 3.914739e-18, 
    3.914692e-18, 3.914458e-18, 3.915488e-18, 3.915546e-18, 3.916463e-18, 
    3.915639e-18, 3.915295e-18, 3.914387e-18, 3.913868e-18, 3.913368e-18, 
    3.91227e-18, 3.91106e-18, 3.909345e-18, 3.9081e-18, 3.90727e-18, 
    3.907773e-18, 3.90733e-18, 3.907829e-18, 3.908058e-18, 3.905491e-18, 
    3.906939e-18, 3.90475e-18, 3.904868e-18, 3.905865e-18, 3.904855e-18, 
    3.914657e-18, 3.914935e-18, 3.915933e-18, 3.915152e-18, 3.916562e-18, 
    3.915784e-18, 3.915343e-18, 3.913595e-18, 3.913189e-18, 3.912842e-18, 
    3.912135e-18, 3.911239e-18, 3.909676e-18, 3.908303e-18, 3.907039e-18, 
    3.90713e-18, 3.907098e-18, 3.906826e-18, 3.907514e-18, 3.906712e-18, 
    3.906586e-18, 3.906929e-18, 3.904884e-18, 3.905467e-18, 3.904871e-18, 
    3.905247e-18, 3.914842e-18, 3.914369e-18, 3.914626e-18, 3.914148e-18, 
    3.914492e-18, 3.91299e-18, 3.91254e-18, 3.910412e-18, 3.911262e-18, 
    3.909885e-18, 3.911115e-18, 3.910902e-18, 3.909878e-18, 3.911042e-18, 
    3.908397e-18, 3.910224e-18, 3.906815e-18, 3.908673e-18, 3.906701e-18, 
    3.907045e-18, 3.906466e-18, 3.905959e-18, 3.905304e-18, 3.904124e-18, 
    3.904393e-18, 3.903393e-18, 3.913656e-18, 3.913052e-18, 3.913088e-18, 
    3.912444e-18, 3.911972e-18, 3.910929e-18, 3.909277e-18, 3.909892e-18, 
    3.908744e-18, 3.90852e-18, 3.910254e-18, 3.909205e-18, 3.912635e-18, 
    3.912098e-18, 3.912405e-18, 3.913619e-18, 3.909774e-18, 3.911755e-18, 
    3.908083e-18, 3.90915e-18, 3.906034e-18, 3.9076e-18, 3.904546e-18, 
    3.903288e-18, 3.902026e-18, 3.900645e-18, 3.912704e-18, 3.913116e-18, 
    3.912363e-18, 3.911354e-18, 3.910369e-18, 3.909088e-18, 3.908948e-18, 
    3.908714e-18, 3.908085e-18, 3.907565e-18, 3.908656e-18, 3.907433e-18, 
    3.912008e-18, 3.909594e-18, 3.913288e-18, 3.912197e-18, 3.911405e-18, 
    3.911735e-18, 3.909958e-18, 3.909546e-18, 3.907878e-18, 3.90873e-18, 
    3.903613e-18, 3.905876e-18, 3.89954e-18, 3.901317e-18, 3.913264e-18, 
    3.912697e-18, 3.910751e-18, 3.911674e-18, 3.908994e-18, 3.908343e-18, 
    3.907799e-18, 3.907133e-18, 3.907048e-18, 3.906651e-18, 3.907303e-18, 
    3.90667e-18, 3.909086e-18, 3.908003e-18, 3.910953e-18, 3.910244e-18, 
    3.910564e-18, 3.910928e-18, 3.909807e-18, 3.908643e-18, 3.908591e-18, 
    3.908222e-18, 3.907234e-18, 3.908982e-18, 3.903372e-18, 3.90688e-18, 
    3.912081e-18, 3.911029e-18, 3.910844e-18, 3.911258e-18, 3.908409e-18, 
    3.909444e-18, 3.906657e-18, 3.907403e-18, 3.906173e-18, 3.906786e-18, 
    3.906878e-18, 3.90766e-18, 3.908155e-18, 3.909402e-18, 3.910409e-18, 
    3.911194e-18, 3.91101e-18, 3.910146e-18, 3.908565e-18, 3.907053e-18, 
    3.907387e-18, 3.906267e-18, 3.909189e-18, 3.907976e-18, 3.908454e-18, 
    3.907205e-18, 3.909914e-18, 3.90769e-18, 3.910493e-18, 3.910242e-18, 
    3.909464e-18, 3.907913e-18, 3.907529e-18, 3.907169e-18, 3.907385e-18, 
    3.90852e-18, 3.908694e-18, 3.909476e-18, 3.909706e-18, 3.910295e-18, 
    3.910795e-18, 3.910345e-18, 3.909878e-18, 3.908509e-18, 3.907291e-18, 
    3.905956e-18, 3.905619e-18, 3.904131e-18, 3.90538e-18, 3.903358e-18, 
    3.905133e-18, 3.902033e-18, 3.90752e-18, 3.905131e-18, 3.909419e-18, 
    3.90895e-18, 3.90813e-18, 3.906195e-18, 3.90721e-18, 3.906009e-18, 
    3.908698e-18, 3.91013e-18, 3.910467e-18, 3.911151e-18, 3.910451e-18, 
    3.910507e-18, 3.909839e-18, 3.910052e-18, 3.908463e-18, 3.909315e-18, 
    3.906888e-18, 3.906012e-18, 3.903507e-18, 3.901993e-18, 3.900409e-18, 
    3.899725e-18, 3.899515e-18, 3.899428e-18 ;

 MEG_formaldehyde =
  7.832722e-19, 7.829854e-19, 7.830398e-19, 7.828118e-19, 7.829362e-19, 
    7.827885e-19, 7.832116e-19, 7.829762e-19, 7.831251e-19, 7.832431e-19, 
    7.823769e-19, 7.828009e-19, 7.819148e-19, 7.821881e-19, 7.814952e-19, 
    7.819604e-19, 7.814005e-19, 7.815031e-19, 7.811813e-19, 7.812731e-19, 
    7.808734e-19, 7.811388e-19, 7.806579e-19, 7.809338e-19, 7.808927e-19, 
    7.811485e-19, 7.827103e-19, 7.824314e-19, 7.827281e-19, 7.82688e-19, 
    7.827048e-19, 7.829355e-19, 7.830555e-19, 7.832904e-19, 7.832467e-19, 
    7.830722e-19, 7.826698e-19, 7.828027e-19, 7.824574e-19, 7.824651e-19, 
    7.820851e-19, 7.822564e-19, 7.816149e-19, 7.817958e-19, 7.812691e-19, 
    7.814022e-19, 7.812763e-19, 7.813138e-19, 7.812759e-19, 7.814707e-19, 
    7.813875e-19, 7.815574e-19, 7.822254e-19, 7.820306e-19, 7.826152e-19, 
    7.829758e-19, 7.832023e-19, 7.833672e-19, 7.83344e-19, 7.833006e-19, 
    7.830713e-19, 7.828513e-19, 7.826854e-19, 7.825754e-19, 7.824662e-19, 
    7.821506e-19, 7.819717e-19, 7.81581e-19, 7.816469e-19, 7.815317e-19, 
    7.814152e-19, 7.812261e-19, 7.812565e-19, 7.811744e-19, 7.815314e-19, 
    7.812957e-19, 7.816855e-19, 7.815794e-19, 7.824551e-19, 7.82766e-19, 
    7.829142e-19, 7.830301e-19, 7.833263e-19, 7.831228e-19, 7.832034e-19, 
    7.830076e-19, 7.828859e-19, 7.829453e-19, 7.825724e-19, 7.827179e-19, 
    7.819612e-19, 7.822866e-19, 7.814288e-19, 7.816329e-19, 7.813793e-19, 
    7.815077e-19, 7.812891e-19, 7.814858e-19, 7.811423e-19, 7.810696e-19, 
    7.811197e-19, 7.809215e-19, 7.814972e-19, 7.812781e-19, 7.829479e-19, 
    7.829383e-19, 7.828916e-19, 7.830975e-19, 7.831092e-19, 7.832925e-19, 
    7.831277e-19, 7.83059e-19, 7.828774e-19, 7.827736e-19, 7.826737e-19, 
    7.82454e-19, 7.822121e-19, 7.81869e-19, 7.816199e-19, 7.814541e-19, 
    7.815545e-19, 7.81466e-19, 7.815657e-19, 7.816116e-19, 7.810981e-19, 
    7.813878e-19, 7.8095e-19, 7.809735e-19, 7.811731e-19, 7.809709e-19, 
    7.829313e-19, 7.829869e-19, 7.831864e-19, 7.830303e-19, 7.833123e-19, 
    7.831568e-19, 7.830686e-19, 7.82719e-19, 7.826378e-19, 7.825683e-19, 
    7.824269e-19, 7.822478e-19, 7.819351e-19, 7.816607e-19, 7.814077e-19, 
    7.814259e-19, 7.814196e-19, 7.813651e-19, 7.815028e-19, 7.813423e-19, 
    7.813172e-19, 7.813857e-19, 7.809768e-19, 7.810933e-19, 7.809741e-19, 
    7.810494e-19, 7.829684e-19, 7.828738e-19, 7.829252e-19, 7.828296e-19, 
    7.828984e-19, 7.82598e-19, 7.825079e-19, 7.820824e-19, 7.822523e-19, 
    7.819769e-19, 7.822229e-19, 7.821803e-19, 7.819757e-19, 7.822084e-19, 
    7.816794e-19, 7.820447e-19, 7.81363e-19, 7.817346e-19, 7.813401e-19, 
    7.814088e-19, 7.812932e-19, 7.811918e-19, 7.810608e-19, 7.808248e-19, 
    7.808786e-19, 7.806785e-19, 7.827312e-19, 7.826104e-19, 7.826177e-19, 
    7.824888e-19, 7.823944e-19, 7.821857e-19, 7.818554e-19, 7.819783e-19, 
    7.817488e-19, 7.817039e-19, 7.820507e-19, 7.81841e-19, 7.82527e-19, 
    7.824196e-19, 7.82481e-19, 7.827236e-19, 7.819548e-19, 7.82351e-19, 
    7.816165e-19, 7.8183e-19, 7.812067e-19, 7.815199e-19, 7.809091e-19, 
    7.806575e-19, 7.804052e-19, 7.801291e-19, 7.825408e-19, 7.826232e-19, 
    7.824725e-19, 7.822707e-19, 7.820737e-19, 7.818177e-19, 7.817895e-19, 
    7.817427e-19, 7.816169e-19, 7.81513e-19, 7.817312e-19, 7.814866e-19, 
    7.824016e-19, 7.819188e-19, 7.826575e-19, 7.824395e-19, 7.82281e-19, 
    7.82347e-19, 7.819915e-19, 7.819091e-19, 7.815756e-19, 7.81746e-19, 
    7.807226e-19, 7.811752e-19, 7.799079e-19, 7.802634e-19, 7.826528e-19, 
    7.825394e-19, 7.821502e-19, 7.823347e-19, 7.817987e-19, 7.816686e-19, 
    7.815597e-19, 7.814265e-19, 7.814095e-19, 7.813301e-19, 7.814606e-19, 
    7.81334e-19, 7.818171e-19, 7.816005e-19, 7.821905e-19, 7.820488e-19, 
    7.821128e-19, 7.821856e-19, 7.819614e-19, 7.817286e-19, 7.817181e-19, 
    7.816444e-19, 7.814468e-19, 7.817964e-19, 7.806745e-19, 7.813761e-19, 
    7.824161e-19, 7.822057e-19, 7.821689e-19, 7.822515e-19, 7.816819e-19, 
    7.818888e-19, 7.813313e-19, 7.814806e-19, 7.812347e-19, 7.813573e-19, 
    7.813756e-19, 7.81532e-19, 7.81631e-19, 7.818803e-19, 7.820818e-19, 
    7.822388e-19, 7.822018e-19, 7.820293e-19, 7.817131e-19, 7.814105e-19, 
    7.814774e-19, 7.812533e-19, 7.818377e-19, 7.815953e-19, 7.816907e-19, 
    7.814409e-19, 7.819828e-19, 7.81538e-19, 7.820987e-19, 7.820483e-19, 
    7.818928e-19, 7.815826e-19, 7.815057e-19, 7.814338e-19, 7.814771e-19, 
    7.81704e-19, 7.817388e-19, 7.818952e-19, 7.819412e-19, 7.820588e-19, 
    7.821589e-19, 7.820689e-19, 7.819755e-19, 7.817017e-19, 7.814582e-19, 
    7.811912e-19, 7.811237e-19, 7.808262e-19, 7.810759e-19, 7.806716e-19, 
    7.810266e-19, 7.804067e-19, 7.81504e-19, 7.810262e-19, 7.818838e-19, 
    7.817899e-19, 7.81626e-19, 7.812389e-19, 7.81442e-19, 7.812018e-19, 
    7.817397e-19, 7.820261e-19, 7.820933e-19, 7.822303e-19, 7.820902e-19, 
    7.821013e-19, 7.819677e-19, 7.820103e-19, 7.816925e-19, 7.818629e-19, 
    7.813776e-19, 7.812023e-19, 7.807014e-19, 7.803984e-19, 7.800818e-19, 
    7.79945e-19, 7.799029e-19, 7.798856e-19 ;

 MEG_isoprene =
  6.252748e-19, 6.250058e-19, 6.250568e-19, 6.248429e-19, 6.249596e-19, 
    6.24821e-19, 6.25218e-19, 6.249971e-19, 6.251368e-19, 6.252475e-19, 
    6.244349e-19, 6.248327e-19, 6.240013e-19, 6.242577e-19, 6.236076e-19, 
    6.240441e-19, 6.235188e-19, 6.23615e-19, 6.23313e-19, 6.233991e-19, 
    6.230241e-19, 6.232731e-19, 6.228218e-19, 6.230808e-19, 6.230422e-19, 
    6.232822e-19, 6.247476e-19, 6.24486e-19, 6.247644e-19, 6.247268e-19, 
    6.247425e-19, 6.24959e-19, 6.250716e-19, 6.252919e-19, 6.252509e-19, 
    6.250872e-19, 6.247097e-19, 6.248344e-19, 6.245105e-19, 6.245176e-19, 
    6.241611e-19, 6.243219e-19, 6.237199e-19, 6.238897e-19, 6.233955e-19, 
    6.235204e-19, 6.234022e-19, 6.234373e-19, 6.234017e-19, 6.235846e-19, 
    6.235066e-19, 6.23666e-19, 6.242928e-19, 6.2411e-19, 6.246585e-19, 
    6.249967e-19, 6.252092e-19, 6.25364e-19, 6.253421e-19, 6.253014e-19, 
    6.250863e-19, 6.248799e-19, 6.247243e-19, 6.246211e-19, 6.245187e-19, 
    6.242225e-19, 6.240547e-19, 6.236881e-19, 6.237499e-19, 6.236419e-19, 
    6.235326e-19, 6.233551e-19, 6.233836e-19, 6.233065e-19, 6.236416e-19, 
    6.234204e-19, 6.237862e-19, 6.236866e-19, 6.245082e-19, 6.247999e-19, 
    6.24939e-19, 6.250477e-19, 6.253256e-19, 6.251346e-19, 6.252103e-19, 
    6.250266e-19, 6.249125e-19, 6.249681e-19, 6.246182e-19, 6.247548e-19, 
    6.240449e-19, 6.243501e-19, 6.235453e-19, 6.237368e-19, 6.234989e-19, 
    6.236194e-19, 6.234142e-19, 6.235988e-19, 6.232764e-19, 6.232083e-19, 
    6.232552e-19, 6.230692e-19, 6.236095e-19, 6.234038e-19, 6.249705e-19, 
    6.249616e-19, 6.249177e-19, 6.25111e-19, 6.251218e-19, 6.252939e-19, 
    6.251392e-19, 6.250748e-19, 6.249045e-19, 6.24807e-19, 6.247133e-19, 
    6.245072e-19, 6.242802e-19, 6.239584e-19, 6.237246e-19, 6.23569e-19, 
    6.236633e-19, 6.235802e-19, 6.236737e-19, 6.237168e-19, 6.232349e-19, 
    6.235068e-19, 6.230959e-19, 6.231181e-19, 6.233053e-19, 6.231155e-19, 
    6.24955e-19, 6.250072e-19, 6.251944e-19, 6.250479e-19, 6.253124e-19, 
    6.251665e-19, 6.250838e-19, 6.247558e-19, 6.246796e-19, 6.246145e-19, 
    6.244818e-19, 6.243137e-19, 6.240204e-19, 6.237628e-19, 6.235255e-19, 
    6.235426e-19, 6.235367e-19, 6.234855e-19, 6.236147e-19, 6.234642e-19, 
    6.234405e-19, 6.235049e-19, 6.231211e-19, 6.232304e-19, 6.231185e-19, 
    6.231892e-19, 6.249898e-19, 6.249011e-19, 6.249493e-19, 6.248596e-19, 
    6.249241e-19, 6.246423e-19, 6.245578e-19, 6.241586e-19, 6.24318e-19, 
    6.240596e-19, 6.242904e-19, 6.242505e-19, 6.240584e-19, 6.242767e-19, 
    6.237804e-19, 6.241232e-19, 6.234836e-19, 6.238323e-19, 6.234621e-19, 
    6.235266e-19, 6.234181e-19, 6.233229e-19, 6.231999e-19, 6.229784e-19, 
    6.23029e-19, 6.22841e-19, 6.247673e-19, 6.24654e-19, 6.246607e-19, 
    6.245399e-19, 6.244513e-19, 6.242554e-19, 6.239455e-19, 6.240609e-19, 
    6.238455e-19, 6.238034e-19, 6.241288e-19, 6.23932e-19, 6.245756e-19, 
    6.244749e-19, 6.245325e-19, 6.247602e-19, 6.240388e-19, 6.244106e-19, 
    6.237214e-19, 6.239218e-19, 6.233369e-19, 6.236308e-19, 6.230576e-19, 
    6.228214e-19, 6.225845e-19, 6.223254e-19, 6.245886e-19, 6.246659e-19, 
    6.245246e-19, 6.243352e-19, 6.241504e-19, 6.239102e-19, 6.238838e-19, 
    6.238398e-19, 6.237218e-19, 6.236243e-19, 6.23829e-19, 6.235995e-19, 
    6.24458e-19, 6.240051e-19, 6.246982e-19, 6.244936e-19, 6.243449e-19, 
    6.244068e-19, 6.240733e-19, 6.239959e-19, 6.23683e-19, 6.238429e-19, 
    6.228825e-19, 6.233073e-19, 6.221176e-19, 6.224514e-19, 6.246937e-19, 
    6.245873e-19, 6.242222e-19, 6.243953e-19, 6.238924e-19, 6.237703e-19, 
    6.236682e-19, 6.235431e-19, 6.235272e-19, 6.234527e-19, 6.235752e-19, 
    6.234563e-19, 6.239097e-19, 6.237064e-19, 6.2426e-19, 6.241271e-19, 
    6.241871e-19, 6.242554e-19, 6.240451e-19, 6.238266e-19, 6.238167e-19, 
    6.237476e-19, 6.235622e-19, 6.238902e-19, 6.228373e-19, 6.234958e-19, 
    6.244717e-19, 6.242742e-19, 6.242397e-19, 6.243172e-19, 6.237827e-19, 
    6.239769e-19, 6.234538e-19, 6.235939e-19, 6.233631e-19, 6.234782e-19, 
    6.234954e-19, 6.236421e-19, 6.23735e-19, 6.239689e-19, 6.24158e-19, 
    6.243053e-19, 6.242706e-19, 6.241087e-19, 6.23812e-19, 6.235281e-19, 
    6.235909e-19, 6.233805e-19, 6.239289e-19, 6.237015e-19, 6.237911e-19, 
    6.235566e-19, 6.240651e-19, 6.236478e-19, 6.241738e-19, 6.241265e-19, 
    6.239806e-19, 6.236896e-19, 6.236175e-19, 6.2355e-19, 6.235906e-19, 
    6.238035e-19, 6.238361e-19, 6.239829e-19, 6.240261e-19, 6.241365e-19, 
    6.242303e-19, 6.241459e-19, 6.240582e-19, 6.238014e-19, 6.235728e-19, 
    6.233223e-19, 6.23259e-19, 6.229798e-19, 6.232141e-19, 6.228346e-19, 
    6.231679e-19, 6.225859e-19, 6.236159e-19, 6.231674e-19, 6.239723e-19, 
    6.238841e-19, 6.237303e-19, 6.233671e-19, 6.235576e-19, 6.233323e-19, 
    6.23837e-19, 6.241057e-19, 6.241688e-19, 6.242973e-19, 6.241659e-19, 
    6.241763e-19, 6.24051e-19, 6.240909e-19, 6.237927e-19, 6.239526e-19, 
    6.234972e-19, 6.233327e-19, 6.228626e-19, 6.225782e-19, 6.222809e-19, 
    6.221525e-19, 6.22113e-19, 6.220968e-19 ;

 MEG_methanol =
  8.573294e-17, 8.571822e-17, 8.572101e-17, 8.570931e-17, 8.571569e-17, 
    8.570811e-17, 8.572983e-17, 8.571775e-17, 8.572539e-17, 8.573145e-17, 
    8.568699e-17, 8.570875e-17, 8.566329e-17, 8.567731e-17, 8.564175e-17, 
    8.566562e-17, 8.56369e-17, 8.564216e-17, 8.562567e-17, 8.563037e-17, 
    8.56099e-17, 8.56235e-17, 8.559887e-17, 8.561299e-17, 8.561089e-17, 
    8.562399e-17, 8.57041e-17, 8.568978e-17, 8.570502e-17, 8.570295e-17, 
    8.570382e-17, 8.571566e-17, 8.572182e-17, 8.573388e-17, 8.573163e-17, 
    8.572267e-17, 8.570203e-17, 8.570884e-17, 8.569113e-17, 8.569152e-17, 
    8.567203e-17, 8.568082e-17, 8.56479e-17, 8.565719e-17, 8.563017e-17, 
    8.5637e-17, 8.563054e-17, 8.563246e-17, 8.563052e-17, 8.56405e-17, 
    8.563624e-17, 8.564495e-17, 8.567923e-17, 8.566923e-17, 8.569922e-17, 
    8.571772e-17, 8.572936e-17, 8.573782e-17, 8.573663e-17, 8.57344e-17, 
    8.572263e-17, 8.571134e-17, 8.570283e-17, 8.569718e-17, 8.569158e-17, 
    8.567538e-17, 8.566621e-17, 8.564615e-17, 8.564954e-17, 8.564363e-17, 
    8.563766e-17, 8.562797e-17, 8.562953e-17, 8.562532e-17, 8.564361e-17, 
    8.563153e-17, 8.565153e-17, 8.564608e-17, 8.5691e-17, 8.570696e-17, 
    8.571457e-17, 8.572051e-17, 8.573572e-17, 8.572527e-17, 8.572941e-17, 
    8.571936e-17, 8.571312e-17, 8.571616e-17, 8.569702e-17, 8.570449e-17, 
    8.566567e-17, 8.568237e-17, 8.563836e-17, 8.564882e-17, 8.563582e-17, 
    8.56424e-17, 8.56312e-17, 8.564128e-17, 8.562368e-17, 8.561995e-17, 
    8.562252e-17, 8.561237e-17, 8.564186e-17, 8.563063e-17, 8.571629e-17, 
    8.57158e-17, 8.571341e-17, 8.572398e-17, 8.572457e-17, 8.573399e-17, 
    8.572552e-17, 8.5722e-17, 8.571268e-17, 8.570735e-17, 8.570222e-17, 
    8.569095e-17, 8.567854e-17, 8.566094e-17, 8.564815e-17, 8.563965e-17, 
    8.56448e-17, 8.564026e-17, 8.564537e-17, 8.564773e-17, 8.562141e-17, 
    8.563626e-17, 8.561383e-17, 8.561503e-17, 8.562525e-17, 8.561489e-17, 
    8.571544e-17, 8.57183e-17, 8.572854e-17, 8.572052e-17, 8.5735e-17, 
    8.572701e-17, 8.572249e-17, 8.570455e-17, 8.570038e-17, 8.569682e-17, 
    8.568957e-17, 8.568038e-17, 8.566433e-17, 8.565024e-17, 8.563727e-17, 
    8.563821e-17, 8.563789e-17, 8.563509e-17, 8.564214e-17, 8.563393e-17, 
    8.563264e-17, 8.563615e-17, 8.56152e-17, 8.562117e-17, 8.561506e-17, 
    8.561892e-17, 8.571735e-17, 8.571249e-17, 8.571513e-17, 8.571022e-17, 
    8.571375e-17, 8.569833e-17, 8.569371e-17, 8.567189e-17, 8.568061e-17, 
    8.566647e-17, 8.56791e-17, 8.567691e-17, 8.56664e-17, 8.567836e-17, 
    8.565121e-17, 8.566995e-17, 8.563498e-17, 8.565404e-17, 8.563381e-17, 
    8.563733e-17, 8.563141e-17, 8.562621e-17, 8.56195e-17, 8.560742e-17, 
    8.561017e-17, 8.559993e-17, 8.570518e-17, 8.569898e-17, 8.569935e-17, 
    8.569274e-17, 8.56879e-17, 8.567719e-17, 8.566024e-17, 8.566655e-17, 
    8.565477e-17, 8.565247e-17, 8.567026e-17, 8.56595e-17, 8.569469e-17, 
    8.568919e-17, 8.569234e-17, 8.570479e-17, 8.566534e-17, 8.568567e-17, 
    8.564797e-17, 8.565894e-17, 8.562698e-17, 8.564302e-17, 8.561173e-17, 
    8.559885e-17, 8.558594e-17, 8.557182e-17, 8.56954e-17, 8.569963e-17, 
    8.56919e-17, 8.568155e-17, 8.567144e-17, 8.56583e-17, 8.565686e-17, 
    8.565446e-17, 8.5648e-17, 8.564267e-17, 8.565386e-17, 8.564132e-17, 
    8.568826e-17, 8.566349e-17, 8.570139e-17, 8.569021e-17, 8.568208e-17, 
    8.568546e-17, 8.566722e-17, 8.5663e-17, 8.564588e-17, 8.565463e-17, 
    8.560218e-17, 8.562536e-17, 8.556052e-17, 8.557869e-17, 8.570115e-17, 
    8.569534e-17, 8.567537e-17, 8.568483e-17, 8.565734e-17, 8.565066e-17, 
    8.564507e-17, 8.563823e-17, 8.563737e-17, 8.56333e-17, 8.563999e-17, 
    8.56335e-17, 8.565828e-17, 8.564716e-17, 8.567744e-17, 8.567016e-17, 
    8.567345e-17, 8.567718e-17, 8.566568e-17, 8.565374e-17, 8.56532e-17, 
    8.56494e-17, 8.563927e-17, 8.565721e-17, 8.559971e-17, 8.563564e-17, 
    8.568901e-17, 8.567821e-17, 8.567632e-17, 8.568057e-17, 8.565134e-17, 
    8.566195e-17, 8.563336e-17, 8.564101e-17, 8.562841e-17, 8.563469e-17, 
    8.563563e-17, 8.564365e-17, 8.564872e-17, 8.566152e-17, 8.567186e-17, 
    8.567992e-17, 8.567802e-17, 8.566916e-17, 8.565294e-17, 8.563742e-17, 
    8.564085e-17, 8.562936e-17, 8.565933e-17, 8.564689e-17, 8.565179e-17, 
    8.563897e-17, 8.566677e-17, 8.564394e-17, 8.567272e-17, 8.567014e-17, 
    8.566216e-17, 8.564623e-17, 8.56423e-17, 8.563861e-17, 8.564083e-17, 
    8.565247e-17, 8.565426e-17, 8.566229e-17, 8.566464e-17, 8.567068e-17, 
    8.567581e-17, 8.56712e-17, 8.56664e-17, 8.565236e-17, 8.563986e-17, 
    8.562618e-17, 8.562272e-17, 8.560748e-17, 8.562027e-17, 8.559956e-17, 
    8.561774e-17, 8.558601e-17, 8.56422e-17, 8.561772e-17, 8.56617e-17, 
    8.565688e-17, 8.564846e-17, 8.562863e-17, 8.563903e-17, 8.562672e-17, 
    8.565431e-17, 8.566899e-17, 8.567245e-17, 8.567948e-17, 8.567229e-17, 
    8.567286e-17, 8.566601e-17, 8.566819e-17, 8.565189e-17, 8.566063e-17, 
    8.563573e-17, 8.562675e-17, 8.56011e-17, 8.55856e-17, 8.556941e-17, 
    8.556242e-17, 8.556027e-17, 8.555939e-17 ;

 MEG_pinene_a =
  7.460949e-17, 7.459335e-17, 7.45964e-17, 7.458357e-17, 7.459057e-17, 
    7.458225e-17, 7.460608e-17, 7.459282e-17, 7.460121e-17, 7.460785e-17, 
    7.455909e-17, 7.458295e-17, 7.453308e-17, 7.454846e-17, 7.450946e-17, 
    7.453564e-17, 7.450414e-17, 7.450991e-17, 7.449182e-17, 7.449698e-17, 
    7.447451e-17, 7.448943e-17, 7.44624e-17, 7.447791e-17, 7.44756e-17, 
    7.448998e-17, 7.457786e-17, 7.456215e-17, 7.457886e-17, 7.45766e-17, 
    7.457755e-17, 7.459054e-17, 7.459729e-17, 7.461052e-17, 7.460806e-17, 
    7.459823e-17, 7.457557e-17, 7.458306e-17, 7.456362e-17, 7.456405e-17, 
    7.454267e-17, 7.455231e-17, 7.45162e-17, 7.452639e-17, 7.449676e-17, 
    7.450424e-17, 7.449716e-17, 7.449927e-17, 7.449714e-17, 7.45081e-17, 
    7.450342e-17, 7.451297e-17, 7.455057e-17, 7.45396e-17, 7.45725e-17, 
    7.45928e-17, 7.460556e-17, 7.461485e-17, 7.461354e-17, 7.461109e-17, 
    7.459818e-17, 7.458579e-17, 7.457645e-17, 7.457027e-17, 7.456412e-17, 
    7.454635e-17, 7.453629e-17, 7.45143e-17, 7.4518e-17, 7.451152e-17, 
    7.450497e-17, 7.449434e-17, 7.449605e-17, 7.449143e-17, 7.45115e-17, 
    7.449825e-17, 7.452019e-17, 7.45142e-17, 7.456348e-17, 7.458099e-17, 
    7.458933e-17, 7.459586e-17, 7.461254e-17, 7.460108e-17, 7.460562e-17, 
    7.45946e-17, 7.458774e-17, 7.459108e-17, 7.457009e-17, 7.457829e-17, 
    7.45357e-17, 7.455401e-17, 7.450574e-17, 7.451721e-17, 7.450295e-17, 
    7.451017e-17, 7.449788e-17, 7.450894e-17, 7.448963e-17, 7.448554e-17, 
    7.448836e-17, 7.447722e-17, 7.450958e-17, 7.449726e-17, 7.459123e-17, 
    7.459069e-17, 7.458806e-17, 7.459965e-17, 7.460031e-17, 7.461064e-17, 
    7.460135e-17, 7.459748e-17, 7.458727e-17, 7.458142e-17, 7.457579e-17, 
    7.456343e-17, 7.454981e-17, 7.453051e-17, 7.451649e-17, 7.450716e-17, 
    7.451281e-17, 7.450782e-17, 7.451344e-17, 7.451602e-17, 7.448714e-17, 
    7.450343e-17, 7.447882e-17, 7.448014e-17, 7.449135e-17, 7.447999e-17, 
    7.45903e-17, 7.459343e-17, 7.460466e-17, 7.459587e-17, 7.461175e-17, 
    7.460299e-17, 7.459803e-17, 7.457835e-17, 7.457377e-17, 7.456986e-17, 
    7.45619e-17, 7.455183e-17, 7.453423e-17, 7.451878e-17, 7.450455e-17, 
    7.450557e-17, 7.450522e-17, 7.450215e-17, 7.45099e-17, 7.450088e-17, 
    7.449946e-17, 7.450331e-17, 7.448033e-17, 7.448687e-17, 7.448017e-17, 
    7.44844e-17, 7.459238e-17, 7.458706e-17, 7.458995e-17, 7.458457e-17, 
    7.458844e-17, 7.457153e-17, 7.456646e-17, 7.454251e-17, 7.455208e-17, 
    7.453658e-17, 7.455043e-17, 7.454803e-17, 7.45365e-17, 7.454961e-17, 
    7.451983e-17, 7.454039e-17, 7.450203e-17, 7.452294e-17, 7.450075e-17, 
    7.450461e-17, 7.449812e-17, 7.449241e-17, 7.448505e-17, 7.447178e-17, 
    7.447481e-17, 7.446356e-17, 7.457903e-17, 7.457223e-17, 7.457264e-17, 
    7.456539e-17, 7.456008e-17, 7.454833e-17, 7.452973e-17, 7.453666e-17, 
    7.452374e-17, 7.452122e-17, 7.454073e-17, 7.452893e-17, 7.456753e-17, 
    7.456149e-17, 7.456495e-17, 7.45786e-17, 7.453533e-17, 7.455763e-17, 
    7.451629e-17, 7.452831e-17, 7.449325e-17, 7.451085e-17, 7.447652e-17, 
    7.446238e-17, 7.444821e-17, 7.443271e-17, 7.456831e-17, 7.457295e-17, 
    7.456447e-17, 7.455311e-17, 7.454202e-17, 7.452762e-17, 7.452604e-17, 
    7.45234e-17, 7.451631e-17, 7.451047e-17, 7.452275e-17, 7.450899e-17, 
    7.456047e-17, 7.453331e-17, 7.457489e-17, 7.456261e-17, 7.45537e-17, 
    7.455741e-17, 7.45374e-17, 7.453276e-17, 7.451398e-17, 7.452358e-17, 
    7.446603e-17, 7.449147e-17, 7.44203e-17, 7.444025e-17, 7.457462e-17, 
    7.456823e-17, 7.454633e-17, 7.455672e-17, 7.452655e-17, 7.451923e-17, 
    7.45131e-17, 7.45056e-17, 7.450465e-17, 7.450019e-17, 7.450753e-17, 
    7.450041e-17, 7.452758e-17, 7.451539e-17, 7.454861e-17, 7.454063e-17, 
    7.454423e-17, 7.454832e-17, 7.453571e-17, 7.452261e-17, 7.452202e-17, 
    7.451786e-17, 7.450674e-17, 7.452642e-17, 7.446333e-17, 7.450276e-17, 
    7.45613e-17, 7.454945e-17, 7.454738e-17, 7.455203e-17, 7.451997e-17, 
    7.453161e-17, 7.450025e-17, 7.450865e-17, 7.449482e-17, 7.450172e-17, 
    7.450275e-17, 7.451154e-17, 7.451711e-17, 7.453114e-17, 7.454248e-17, 
    7.455132e-17, 7.454924e-17, 7.453952e-17, 7.452173e-17, 7.450471e-17, 
    7.450847e-17, 7.449587e-17, 7.452875e-17, 7.45151e-17, 7.452048e-17, 
    7.450641e-17, 7.453691e-17, 7.451187e-17, 7.454343e-17, 7.45406e-17, 
    7.453185e-17, 7.451438e-17, 7.451006e-17, 7.450602e-17, 7.450845e-17, 
    7.452122e-17, 7.452318e-17, 7.453198e-17, 7.453457e-17, 7.454119e-17, 
    7.454683e-17, 7.454176e-17, 7.45365e-17, 7.452109e-17, 7.450738e-17, 
    7.449238e-17, 7.448858e-17, 7.447186e-17, 7.448589e-17, 7.446317e-17, 
    7.448311e-17, 7.444829e-17, 7.450996e-17, 7.448309e-17, 7.453134e-17, 
    7.452605e-17, 7.451682e-17, 7.449506e-17, 7.450647e-17, 7.449297e-17, 
    7.452323e-17, 7.453934e-17, 7.454313e-17, 7.455084e-17, 7.454296e-17, 
    7.454358e-17, 7.453606e-17, 7.453846e-17, 7.452058e-17, 7.453016e-17, 
    7.450285e-17, 7.449299e-17, 7.446485e-17, 7.444783e-17, 7.443006e-17, 
    7.442239e-17, 7.442002e-17, 7.441905e-17 ;

 MEG_thujene_a =
  1.79764e-18, 1.79728e-18, 1.797348e-18, 1.797063e-18, 1.797219e-18, 
    1.797034e-18, 1.797564e-18, 1.797269e-18, 1.797455e-18, 1.797603e-18, 
    1.796518e-18, 1.797049e-18, 1.79594e-18, 1.796282e-18, 1.795415e-18, 
    1.795997e-18, 1.795297e-18, 1.795425e-18, 1.795023e-18, 1.795137e-18, 
    1.794638e-18, 1.79497e-18, 1.794369e-18, 1.794713e-18, 1.794662e-18, 
    1.794982e-18, 1.796936e-18, 1.796587e-18, 1.796958e-18, 1.796908e-18, 
    1.796929e-18, 1.797218e-18, 1.797368e-18, 1.797662e-18, 1.797608e-18, 
    1.797389e-18, 1.796885e-18, 1.797052e-18, 1.79662e-18, 1.796629e-18, 
    1.796153e-18, 1.796368e-18, 1.795565e-18, 1.795791e-18, 1.795132e-18, 
    1.795299e-18, 1.795141e-18, 1.795188e-18, 1.795141e-18, 1.795384e-18, 
    1.79528e-18, 1.795493e-18, 1.796329e-18, 1.796085e-18, 1.796817e-18, 
    1.797268e-18, 1.797552e-18, 1.797759e-18, 1.79773e-18, 1.797675e-18, 
    1.797388e-18, 1.797113e-18, 1.796905e-18, 1.796767e-18, 1.796631e-18, 
    1.796235e-18, 1.796011e-18, 1.795522e-18, 1.795605e-18, 1.795461e-18, 
    1.795315e-18, 1.795079e-18, 1.795117e-18, 1.795014e-18, 1.79546e-18, 
    1.795166e-18, 1.795653e-18, 1.79552e-18, 1.796616e-18, 1.797006e-18, 
    1.797191e-18, 1.797336e-18, 1.797707e-18, 1.797452e-18, 1.797553e-18, 
    1.797308e-18, 1.797156e-18, 1.79723e-18, 1.796763e-18, 1.796945e-18, 
    1.795998e-18, 1.796406e-18, 1.795332e-18, 1.795587e-18, 1.79527e-18, 
    1.795431e-18, 1.795157e-18, 1.795403e-18, 1.794974e-18, 1.794883e-18, 
    1.794946e-18, 1.794698e-18, 1.795418e-18, 1.795144e-18, 1.797233e-18, 
    1.797221e-18, 1.797163e-18, 1.797421e-18, 1.797435e-18, 1.797665e-18, 
    1.797459e-18, 1.797372e-18, 1.797145e-18, 1.797015e-18, 1.79689e-18, 
    1.796615e-18, 1.796312e-18, 1.795883e-18, 1.795571e-18, 1.795364e-18, 
    1.795489e-18, 1.795379e-18, 1.795503e-18, 1.795561e-18, 1.794919e-18, 
    1.795281e-18, 1.794734e-18, 1.794763e-18, 1.795012e-18, 1.79476e-18, 
    1.797213e-18, 1.797282e-18, 1.797532e-18, 1.797337e-18, 1.79769e-18, 
    1.797495e-18, 1.797385e-18, 1.796947e-18, 1.796845e-18, 1.796758e-18, 
    1.796581e-18, 1.796357e-18, 1.795966e-18, 1.795622e-18, 1.795306e-18, 
    1.795329e-18, 1.795321e-18, 1.795252e-18, 1.795424e-18, 1.795224e-18, 
    1.795192e-18, 1.795278e-18, 1.794767e-18, 1.794913e-18, 1.794764e-18, 
    1.794858e-18, 1.797259e-18, 1.797141e-18, 1.797205e-18, 1.797085e-18, 
    1.797171e-18, 1.796795e-18, 1.796683e-18, 1.79615e-18, 1.796363e-18, 
    1.796018e-18, 1.796326e-18, 1.796273e-18, 1.796016e-18, 1.796308e-18, 
    1.795646e-18, 1.796103e-18, 1.79525e-18, 1.795715e-18, 1.795221e-18, 
    1.795307e-18, 1.795162e-18, 1.795036e-18, 1.794872e-18, 1.794577e-18, 
    1.794644e-18, 1.794394e-18, 1.796962e-18, 1.796811e-18, 1.79682e-18, 
    1.796659e-18, 1.796541e-18, 1.796279e-18, 1.795866e-18, 1.79602e-18, 
    1.795732e-18, 1.795676e-18, 1.79611e-18, 1.795848e-18, 1.796706e-18, 
    1.796572e-18, 1.796649e-18, 1.796953e-18, 1.79599e-18, 1.796486e-18, 
    1.795567e-18, 1.795834e-18, 1.795054e-18, 1.795446e-18, 1.794682e-18, 
    1.794368e-18, 1.794053e-18, 1.793708e-18, 1.796724e-18, 1.796827e-18, 
    1.796638e-18, 1.796386e-18, 1.796139e-18, 1.795819e-18, 1.795783e-18, 
    1.795725e-18, 1.795567e-18, 1.795437e-18, 1.79571e-18, 1.795404e-18, 
    1.796549e-18, 1.795945e-18, 1.79687e-18, 1.796597e-18, 1.796399e-18, 
    1.796481e-18, 1.796036e-18, 1.795933e-18, 1.795515e-18, 1.795729e-18, 
    1.794449e-18, 1.795015e-18, 1.793433e-18, 1.793876e-18, 1.796864e-18, 
    1.796722e-18, 1.796235e-18, 1.796466e-18, 1.795795e-18, 1.795632e-18, 
    1.795496e-18, 1.795329e-18, 1.795308e-18, 1.795209e-18, 1.795372e-18, 
    1.795214e-18, 1.795818e-18, 1.795547e-18, 1.796285e-18, 1.796108e-18, 
    1.796188e-18, 1.796279e-18, 1.795999e-18, 1.795707e-18, 1.795694e-18, 
    1.795602e-18, 1.795354e-18, 1.795792e-18, 1.794389e-18, 1.795266e-18, 
    1.796568e-18, 1.796304e-18, 1.796258e-18, 1.796362e-18, 1.795649e-18, 
    1.795908e-18, 1.79521e-18, 1.795397e-18, 1.795089e-18, 1.795243e-18, 
    1.795265e-18, 1.795461e-18, 1.795585e-18, 1.795897e-18, 1.796149e-18, 
    1.796346e-18, 1.7963e-18, 1.796084e-18, 1.795688e-18, 1.795309e-18, 
    1.795393e-18, 1.795113e-18, 1.795844e-18, 1.79554e-18, 1.79566e-18, 
    1.795347e-18, 1.796025e-18, 1.795469e-18, 1.79617e-18, 1.796107e-18, 
    1.795913e-18, 1.795524e-18, 1.795428e-18, 1.795338e-18, 1.795392e-18, 
    1.795676e-18, 1.79572e-18, 1.795916e-18, 1.795973e-18, 1.796121e-18, 
    1.796246e-18, 1.796133e-18, 1.796016e-18, 1.795674e-18, 1.795369e-18, 
    1.795035e-18, 1.794951e-18, 1.794579e-18, 1.794891e-18, 1.794386e-18, 
    1.794829e-18, 1.794055e-18, 1.795426e-18, 1.794828e-18, 1.795902e-18, 
    1.795784e-18, 1.795579e-18, 1.795095e-18, 1.795348e-18, 1.795048e-18, 
    1.795721e-18, 1.796079e-18, 1.796164e-18, 1.796335e-18, 1.79616e-18, 
    1.796174e-18, 1.796006e-18, 1.79606e-18, 1.795662e-18, 1.795875e-18, 
    1.795268e-18, 1.795049e-18, 1.794423e-18, 1.794045e-18, 1.79365e-18, 
    1.793479e-18, 1.793427e-18, 1.793405e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  9.889298e-26, -1.455922e-25, 1.593275e-25, -3.43378e-25, 1.373521e-26, 
    8.515785e-26, 2.060269e-25, -3.488721e-25, -1.098809e-25, -9.889281e-26, 
    -2.36244e-25, -1.400982e-25, -6.098394e-25, -2.746942e-27, -2.747024e-25, 
    -4.395239e-25, -4.285358e-25, -1.016398e-25, -2.664613e-25, 
    -1.071339e-25, -1.840506e-25, -4.944636e-26, -2.3075e-25, -3.983185e-25, 
    3.433782e-25, -4.395231e-26, 1.758097e-25, -3.928245e-25, -3.790893e-25, 
    1.400983e-25, 3.351371e-25, 3.57114e-26, 4.532592e-25, -4.724882e-25, 
    -5.493967e-27, 2.719555e-25, 3.351371e-25, 2.747107e-27, -1.318571e-25, 
    4.120538e-25, 4.010657e-25, -3.571124e-26, -5.301757e-25, -3.186548e-25, 
    -1.126279e-25, 2.582204e-25, -4.944636e-26, -2.746942e-27, -1.895446e-25, 
    -4.120536e-25, -9.614578e-26, -7.691661e-26, -3.571131e-25, 
    -9.614578e-26, -1.098802e-26, 2.197628e-26, 1.758097e-25, 2.197621e-25, 
    -1.263631e-25, -1.813036e-25, -4.175477e-25, -1.346041e-25, 
    -1.318571e-25, -3.571124e-26, -3.598602e-25, 4.202949e-25, -1.758095e-25, 
    -1.483393e-25, -3.845826e-26, 2.280031e-25, 1.455924e-25, -1.346041e-25, 
    -4.230417e-25, 2.08774e-25, 4.807294e-25, 3.681014e-25, -2.060268e-25, 
    1.263632e-25, 2.747033e-26, 3.296438e-26, 3.296438e-26, -3.37884e-25, 
    3.131609e-25, 3.708484e-25, -9.339876e-26, 2.747026e-25, 1.291103e-25, 
    1.04387e-25, -7.966364e-26, 1.098811e-25, 1.428454e-25, 1.428454e-25, 
    5.76876e-26, -1.593274e-25, 4.120545e-26, 2.774496e-25, 1.126281e-25, 
    -7.691661e-26, -9.065174e-26, 3.818365e-25, -2.856905e-25, -1.098802e-26, 
    1.263632e-25, -1.126279e-25, -1.400982e-25, 4.395248e-26, -2.719554e-25, 
    -2.472314e-26, -2.746942e-27, 1.977859e-25, -1.785565e-25, -2.746942e-27, 
    1.400983e-25, 2.856907e-25, -7.142256e-26, -2.472321e-25, 1.730626e-25, 
    -1.922916e-25, 3.57114e-26, -3.845826e-26, 4.669943e-25, 3.57114e-26, 
    -2.554732e-25, 1.703156e-25, 2.252561e-25, 1.922926e-26, -2.197612e-26, 
    -3.021727e-25, 3.845843e-26, 8.241157e-27, 2.472331e-26, -3.571131e-25, 
    8.515785e-26, -4.395231e-26, 2.307502e-25, -4.065596e-25, 1.428454e-25, 
    -5.686341e-25, 1.813037e-25, 2.692085e-25, 1.0164e-25, -4.202947e-25, 
    1.593275e-25, -3.516191e-25, -8.790471e-26, -3.543661e-25, 1.373521e-26, 
    -3.186548e-25, -2.444851e-25, 9.614595e-26, -1.758095e-25, 1.181221e-25, 
    2.856907e-25, -3.37884e-25, -3.983185e-25, -5.768744e-26, -2.554732e-25, 
    -7.691661e-26, -4.50512e-25, 2.417383e-25, -4.724882e-25, -1.977857e-25, 
    -4.395231e-26, -2.747016e-26, -1.263631e-25, -5.439108e-25, -1.20869e-25, 
    3.57114e-26, -4.285358e-25, -2.472321e-25, 2.472331e-26, -6.318148e-26, 
    2.747107e-27, -1.291101e-25, -6.867554e-26, -3.571124e-26, -2.746942e-27, 
    -2.36244e-25, -6.867554e-26, 4.66995e-26, 1.648223e-26, -6.043446e-26, 
    1.867978e-25, -2.856905e-25, 6.070926e-25, -4.834763e-25, 4.175478e-25, 
    2.994258e-25, 1.098818e-26, -2.444851e-25, -1.895446e-25, -1.813036e-25, 
    -1.675684e-25, -5.301757e-25, -1.20869e-25, -3.021719e-26, -2.472321e-25, 
    5.494058e-26, 5.46658e-25, -1.428452e-25, -4.175477e-25, -1.703155e-25, 
    -1.043869e-25, 2.334972e-25, 2.856907e-25, 4.175478e-25, 3.18655e-25, 
    -4.202947e-25, -1.373504e-26, 1.153751e-25, 2.444853e-25, -1.098809e-25, 
    -2.554732e-25, 5.494132e-27, 4.917175e-25, 3.681014e-25, 2.14268e-25, 
    2.719555e-25, -1.813036e-25, 4.3403e-25, 2.609674e-25, 4.560062e-25, 
    -8.515768e-26, 2.801966e-25, -1.648207e-26, 3.845843e-26, -3.186548e-25, 
    3.076668e-25, -5.494041e-26, 1.620745e-25, -3.241488e-25, -5.219346e-25, 
    -6.867561e-25, -2.170149e-25, -7.142256e-26, -5.164406e-25, 
    -7.691661e-26, -9.065174e-26, 5.76876e-26, -9.614578e-26, -1.785565e-25, 
    -3.955715e-25, 3.57114e-26, -2.747016e-26, -6.592851e-26, -9.339876e-26, 
    -4.038125e-25, -4.093066e-25, 6.318165e-26, -8.790471e-26, -1.373504e-26, 
    1.510864e-25, 3.928246e-25, 1.648216e-25, -1.895446e-25, -4.450179e-25, 
    -1.071339e-25, 3.159079e-25, 3.296438e-26, 2.554734e-25, -2.225089e-25, 
    6.318165e-26, -3.268959e-25, -3.46125e-25, 2.994258e-25, 7.96638e-26, 
    6.86757e-26, -2.527262e-25, -5.493967e-27, -7.938901e-25, -2.170149e-25, 
    4.175478e-25, -4.312828e-25, 1.758097e-25, -1.15375e-25, -3.900774e-25, 
    -1.126279e-25, 1.867978e-25, -2.36244e-25, 2.747026e-25, 1.620745e-25, 
    1.455924e-25, 2.994258e-25, 2.197628e-26, -2.087738e-25, 5.384169e-25, 
    2.939317e-25, 1.648223e-26, 7.142273e-26, -1.648214e-25, 5.76876e-26, 
    -1.23616e-25, -1.483393e-25, 2.527264e-25, 4.944653e-26, -2.582203e-25, 
    -5.219339e-26, 3.57114e-26, -1.895446e-25, -5.493967e-27, -1.346041e-25, 
    -4.669934e-26, 8.790487e-26, -2.005327e-25, -3.351369e-25, -3.241488e-25, 
    8.241157e-27, -4.395231e-26, -5.219339e-26, 1.840507e-25, 1.483394e-25, 
    -1.263631e-25, -3.323899e-25, 5.76876e-26, 1.236162e-25, -2.966786e-25, 
    -2.527262e-25, 3.131609e-25, 1.208692e-25, 5.494058e-26, 3.681014e-25, 
    -2.142679e-25, 7.142273e-26, -3.653542e-25, 2.11521e-25, 2.005329e-25, 
    1.977859e-25, 1.181221e-25, 6.318165e-26, -2.747016e-26, -1.648207e-26, 
    -2.582203e-25, -1.15375e-25, -5.768744e-26, -6.318148e-26, -1.071339e-25, 
    3.433782e-25, 3.406311e-25 ;

 M_LITR2C_TO_LEACHING =
  -2.087738e-25, -1.098809e-25, -2.334971e-25, -2.362441e-25, 8.515782e-26, 
    -1.373507e-26, -1.703155e-25, -3.021722e-26, -9.339879e-26, 2.280031e-25, 
    -7.142259e-26, -2.692084e-25, -1.593274e-25, -2.527262e-25, 
    -2.005328e-25, 4.94465e-26, -9.614581e-26, -1.20869e-25, 7.691675e-26, 
    5.494103e-27, 2.005329e-25, -1.867976e-25, 2.14268e-25, 6.592865e-26, 
    -1.318571e-25, -3.104137e-25, -1.538333e-25, 1.373518e-26, 3.790895e-25, 
    1.318572e-25, -3.790894e-25, 3.790895e-25, -2.197614e-26, -2.472317e-26, 
    -7.966367e-26, -1.867976e-25, 4.395245e-26, 1.922923e-26, 2.417382e-25, 
    -1.373512e-25, -1.18122e-25, 1.208691e-25, 1.730626e-25, -2.609673e-25, 
    -1.977857e-25, -2.3075e-25, 2.197625e-26, -2.746971e-27, -3.076667e-25, 
    -7.416961e-26, -1.922912e-26, 2.087739e-25, 1.318572e-25, -2.719554e-25, 
    -7.966367e-26, -4.285358e-25, -1.291101e-25, -1.098809e-25, 7.966377e-26, 
    -2.115208e-25, 1.0164e-25, -6.592854e-26, -6.592854e-26, -4.724882e-25, 
    -2.527262e-25, -5.494044e-26, -1.373512e-25, -1.15375e-25, -4.010656e-25, 
    3.571138e-26, 2.747078e-27, 1.07134e-25, 1.64822e-26, -5.493996e-27, 
    1.236162e-25, 3.84584e-26, -4.257888e-25, -1.263631e-25, 3.296435e-26, 
    3.021733e-26, 1.593275e-25, 2.747025e-25, -5.493996e-27, 2.252561e-25, 
    -2.472322e-25, 5.494055e-26, -1.373512e-25, -2.334971e-25, -4.944639e-26, 
    -1.455923e-25, -1.895447e-25, -4.669937e-26, -6.867557e-26, 3.29643e-25, 
    -2.746971e-27, -3.40631e-25, -6.867557e-26, -9.339879e-26, 1.09881e-25, 
    2.472328e-26, -3.845829e-26, 6.04346e-26, -1.428452e-25, -1.098805e-26, 
    1.620745e-25, -2.3075e-25, -2.142679e-25, 4.395245e-26, 8.24108e-26, 
    -9.339879e-26, 9.339889e-26, -6.043449e-26, -1.867976e-25, 1.208691e-25, 
    6.592865e-26, 1.758096e-25, -4.395234e-26, -2.884375e-25, -9.889284e-26, 
    -3.845829e-26, -1.538333e-25, -7.142259e-26, 6.04346e-26, -2.197614e-26, 
    -3.021727e-25, 2.252561e-25, -1.346042e-25, 3.296435e-26, -1.098805e-26, 
    -3.845829e-26, -1.373512e-25, -5.494044e-26, -1.428452e-25, 
    -2.005328e-25, -1.098805e-26, 8.24108e-26, -4.010656e-25, -4.944639e-26, 
    -3.626072e-25, -2.746971e-27, 6.592865e-26, -2.499792e-25, -3.241489e-25, 
    -1.263631e-25, 2.719555e-25, -2.362441e-25, 1.153751e-25, -2.746971e-27, 
    -9.339879e-26, 6.592865e-26, -1.922917e-25, 7.14227e-26, 2.637144e-25, 
    1.318572e-25, -1.922912e-26, 1.181221e-25, -3.241489e-25, 2.280031e-25, 
    1.922918e-25, 2.966787e-25, -1.510863e-25, 1.208691e-25, -2.582203e-25, 
    -1.071339e-25, -1.840506e-25, -1.703155e-25, 5.219352e-26, -2.115208e-25, 
    9.889295e-26, 2.692085e-25, -1.098809e-25, -1.098809e-25, 5.494055e-26, 
    -1.263631e-25, -2.774495e-25, 7.14227e-26, -5.494044e-26, 3.021728e-25, 
    -2.637143e-25, -2.032798e-25, 4.175478e-25, 1.373518e-26, -2.197619e-25, 
    3.104139e-25, 1.648215e-25, 1.648215e-25, 1.373513e-25, -2.637143e-25, 
    1.346043e-25, -2.472317e-26, 1.510864e-25, 1.785567e-25, -1.373507e-26, 
    -1.703155e-25, 1.758096e-25, 3.29643e-25, -1.867976e-25, 6.04346e-26, 
    2.472328e-26, -1.922912e-26, 1.455924e-25, 2.472328e-26, -3.35137e-25, 
    7.691675e-26, -9.339879e-26, 2.74703e-26, 1.648215e-25, -2.664613e-25, 
    8.515782e-26, -1.18122e-25, -1.483393e-25, -9.065177e-26, -2.362441e-25, 
    2.801966e-25, -4.395234e-26, -1.703155e-25, 9.889295e-26, 8.790485e-26, 
    -2.74702e-26, -1.538333e-25, -1.428452e-25, 1.703156e-25, -3.076667e-25, 
    -1.428452e-25, 5.494103e-27, 5.494055e-26, -1.346042e-25, 4.669947e-26, 
    -8.790474e-26, -4.148007e-25, 1.950388e-25, -2.197619e-25, -3.296424e-26, 
    1.538334e-25, -2.939316e-25, 7.14227e-26, -7.691664e-26, -5.219342e-26, 
    1.64822e-26, -1.510863e-25, -1.538333e-25, -4.669937e-26, 1.867977e-25, 
    -4.944639e-26, 8.241128e-27, 9.614592e-26, 1.675686e-25, 2.307501e-25, 
    -2.637143e-25, 1.09881e-25, 2.252561e-25, 1.648215e-25, 6.592865e-26, 
    -6.867557e-26, 8.241128e-27, 6.318163e-26, -9.339879e-26, -5.493996e-27, 
    -2.856905e-25, -7.416961e-26, 9.614592e-26, -1.20869e-25, 2.801966e-25, 
    -4.120532e-26, -2.829435e-25, -7.691664e-26, -2.994256e-25, 2.527263e-25, 
    8.24108e-26, 1.373518e-26, -2.692084e-25, -5.493996e-27, -5.493996e-27, 
    -1.428452e-25, -2.74702e-26, -2.115208e-25, -1.510863e-25, -1.758095e-25, 
    -1.977857e-25, 1.09881e-25, -2.087738e-25, -4.120532e-26, -1.400982e-25, 
    -1.840506e-25, 1.64822e-26, -2.087738e-25, -2.25256e-25, -2.74702e-26, 
    -2.417381e-25, 3.571138e-26, 3.681014e-25, 1.648215e-25, 5.494103e-27, 
    8.515782e-26, 1.64822e-26, 4.669947e-26, -5.219342e-26, -1.098805e-26, 
    -3.35137e-25, -9.339879e-26, -2.74702e-26, -2.527262e-25, 7.14227e-26, 
    8.790485e-26, -2.582203e-25, 2.911847e-25, -1.593274e-25, -8.241069e-26, 
    -1.840506e-25, -2.197619e-25, -1.346042e-25, 1.208691e-25, 8.790485e-26, 
    2.966787e-25, -4.944639e-26, -9.065177e-26, -2.362441e-25, 1.922923e-26, 
    -7.691664e-26, -5.768747e-26, 2.801966e-25, -2.087738e-25, 6.867567e-26, 
    1.510864e-25, -3.268959e-25, 2.252561e-25, 2.74703e-26, 3.653543e-25, 
    -2.856905e-25, -1.455923e-25, -3.571132e-25, -1.098805e-26, 
    -1.483393e-25, 6.04346e-26, 8.515782e-26, -9.889284e-26, -3.845829e-26, 
    -1.346042e-25 ;

 M_LITR3C_TO_LEACHING =
  -3.57113e-26, 4.395242e-26, -7.279613e-26, -6.592857e-26, 3.159081e-26, 
    9.75194e-26, -1.373512e-25, -8.241071e-26, -6.318154e-26, 1.373513e-25, 
    -6.867559e-26, 1.92292e-26, 3.571135e-26, -1.15375e-25, -1.016399e-25, 
    -1.455923e-25, 2.22509e-25, -3.57113e-26, -2.884373e-26, -9.065179e-26, 
    6.180808e-26, -1.030134e-25, -3.57113e-26, -2.747022e-26, -2.609671e-26, 
    -3.57113e-26, 7.966375e-26, -3.845832e-26, 6.867589e-27, -6.867535e-27, 
    -2.47232e-26, -2.884373e-26, -6.867535e-27, -3.159076e-26, -2.156414e-25, 
    2.197622e-26, -1.648212e-26, 3.296432e-26, 4.12054e-26, -7.966369e-26, 
    -3.021725e-26, -7.966369e-26, -1.002664e-25, -4.532588e-26, 
    -1.758096e-25, -1.208691e-25, -1.785563e-26, 5.081998e-26, -8.241047e-27, 
    -1.140015e-25, -7.691667e-26, -2.609671e-26, 8.653131e-26, -4.807291e-26, 
    1.92292e-26, 5.631404e-26, 3.845837e-26, -7.691667e-26, 1.09881e-25, 
    -1.194956e-25, -4.944642e-26, -7.691667e-26, -1.455923e-25, 
    -2.609671e-26, -7.142262e-26, -5.631398e-26, 4.944647e-26, 1.648217e-26, 
    2.747052e-27, -2.747022e-26, -7.416964e-26, -1.414718e-25, -2.747022e-26, 
    1.09881e-25, 6.043457e-26, 1.277367e-25, -1.648212e-26, -1.414718e-25, 
    6.867565e-26, -6.318154e-26, 9.614614e-27, 1.565804e-25, -6.592857e-26, 
    -1.043869e-25, 9.614614e-27, 1.92292e-26, 1.098813e-26, 1.497129e-25, 
    -1.318572e-25, 7.966375e-26, -5.494023e-27, -1.18122e-25, -6.867559e-26, 
    -3.845832e-26, 1.483394e-25, 8.241101e-27, 2.609676e-26, 3.708486e-26, 
    -2.884373e-26, 1.236164e-26, -5.081993e-26, 2.675708e-32, -2.609671e-26, 
    -8.241071e-26, -1.510863e-25, -5.494047e-26, 1.373515e-26, -3.845832e-26, 
    -8.515774e-26, -1.346042e-25, 8.241101e-27, -1.373486e-27, 3.571135e-26, 
    -4.532588e-26, 1.66195e-25, -7.416964e-26, 7.966375e-26, -1.497128e-25, 
    -8.653126e-26, 2.675714e-32, 2.472325e-26, -9.20253e-26, 5.494076e-27, 
    1.098813e-26, 3.159081e-26, -2.746998e-27, -2.197617e-26, -3.296427e-26, 
    -3.433778e-26, -6.043452e-26, 4.395242e-26, -1.071339e-25, -1.15375e-25, 
    -2.609671e-26, -1.387247e-25, 3.02173e-26, -7.966369e-26, -1.057604e-25, 
    6.180808e-26, -1.922915e-26, 5.494076e-27, -1.428453e-25, -6.592857e-26, 
    -5.494047e-26, -2.417381e-25, -7.966369e-26, -8.378423e-26, 
    -4.669939e-26, 4.257891e-26, -1.359777e-25, 3.159081e-26, 7.416969e-26, 
    -1.455923e-25, 2.472325e-26, 4.944647e-26, -3.433778e-26, -1.510861e-26, 
    -3.845832e-26, 4.395242e-26, -5.494047e-26, 9.614589e-26, 8.515779e-26, 
    -6.867559e-26, -3.021725e-26, 1.593275e-25, 2.675718e-32, 2.197622e-26, 
    -1.208691e-25, -1.400982e-25, 6.31816e-26, -6.867559e-26, -1.675685e-25, 
    1.112545e-25, -1.922915e-26, 1.09881e-25, 2.197622e-26, -7.142262e-26, 
    4.395242e-26, -8.10372e-26, -1.318572e-25, -9.61456e-27, -8.653126e-26, 
    4.12054e-26, -8.378423e-26, 1.04387e-25, -5.631398e-26, -9.614584e-26, 
    -4.257886e-26, 8.241077e-26, -9.339881e-26, 1.112545e-25, -1.400982e-25, 
    1.318572e-25, -3.021725e-26, -5.494047e-26, -3.57113e-26, -5.219344e-26, 
    -1.373486e-27, -1.387247e-25, -1.043869e-25, -1.112545e-25, 
    -6.455506e-26, -5.768749e-26, -1.098807e-26, -6.592857e-26, 
    -1.318572e-25, 6.455511e-26, 1.60701e-25, -1.510861e-26, 4.669945e-26, 
    2.472325e-26, -7.691667e-26, -4.120535e-26, 6.31816e-26, 5.356701e-26, 
    3.845837e-26, -6.318154e-26, -1.236158e-26, 1.785569e-26, 2.197622e-26, 
    -7.279613e-26, -2.747022e-26, 3.983189e-26, 6.31816e-26, -1.648212e-26, 
    -4.944642e-26, 2.747052e-27, -3.021725e-26, 2.472325e-26, 2.197622e-26, 
    2.197622e-26, 1.497129e-25, 1.648217e-26, -2.609671e-26, -8.241047e-27, 
    1.373515e-26, 8.378428e-26, 8.241101e-27, 1.194956e-25, 6.043457e-26, 
    1.565804e-25, -9.889287e-26, -2.060266e-26, 2.675713e-32, 3.571135e-26, 
    -9.339881e-26, 3.296432e-26, -6.318154e-26, -4.120535e-26, 6.592862e-26, 
    5.768755e-26, -6.867535e-27, -2.747022e-26, 4.669945e-26, 7.004916e-26, 
    -1.043869e-25, 7.004916e-26, 1.112545e-25, 1.181221e-25, 2.747028e-26, 
    -1.236161e-25, -1.12628e-25, -1.510861e-26, 6.867589e-27, 6.31816e-26, 
    -1.249896e-25, -3.021725e-26, -1.565804e-25, -3.159076e-26, 8.241101e-27, 
    -5.494023e-27, -3.708481e-26, -4.807291e-26, 1.098813e-26, -2.334968e-26, 
    9.614614e-27, -9.61456e-27, 5.21935e-26, 1.510866e-26, 4.120564e-27, 
    -3.708481e-26, 1.510866e-26, 1.373515e-26, -1.291101e-25, 1.12628e-25, 
    -5.494047e-26, -2.211355e-25, 2.197622e-26, 7.416969e-26, 1.648215e-25, 
    -3.021725e-26, 9.614614e-27, -1.648212e-26, 1.648217e-26, -1.620744e-25, 
    1.236164e-26, -1.37351e-26, -4.257886e-26, 1.016399e-25, -1.098807e-26, 
    4.532594e-26, 5.906106e-26, 5.21935e-26, -2.334968e-26, 2.060271e-26, 
    2.884379e-26, 3.159081e-26, 2.197622e-26, -1.208691e-25, 4.12054e-26, 
    2.197622e-26, -9.889287e-26, -9.614584e-26, -1.675685e-25, -2.746998e-27, 
    3.433784e-26, -1.12628e-25, -9.61456e-27, -2.197617e-26, 2.197622e-26, 
    -2.747022e-26, 8.241101e-27, 3.571135e-26, -2.197617e-26, -7.416964e-26, 
    -3.57113e-26, -1.730625e-25, 2.884379e-26, -4.120535e-26, 1.030135e-25, 
    -6.592857e-26, 9.614589e-26, 1.648217e-26, 1.181221e-25, -2.25256e-25, 
    -2.747022e-26, 4.669945e-26, 9.339887e-26 ;

 M_SOIL1C_TO_LEACHING =
  -4.222318e-21, 2.792506e-20, 3.748973e-22, 1.70597e-20, 2.676189e-20, 
    2.347145e-20, 4.484401e-21, 2.559853e-21, -1.325642e-20, -1.650951e-20, 
    1.428694e-20, -7.925507e-21, -1.737863e-20, 1.155549e-20, -8.323295e-21, 
    -3.944632e-20, 2.821571e-20, 1.765059e-20, 3.659554e-20, 8.786148e-21, 
    -5.881915e-21, -1.124873e-20, 9.405606e-21, -5.841781e-21, 2.091217e-20, 
    -4.586748e-21, -2.403777e-20, -2.680856e-21, 1.416086e-20, 4.608775e-23, 
    2.424756e-20, -3.831849e-20, -2.281977e-20, -2.899291e-20, 1.662061e-20, 
    1.85986e-20, -2.037917e-21, -1.386624e-20, -2.25769e-20, -7.273807e-21, 
    1.072426e-20, -1.940154e-20, 3.257993e-20, 3.26472e-20, 1.288404e-20, 
    5.510147e-21, -8.908964e-22, -4.002363e-20, -1.191088e-20, 1.329344e-20, 
    7.831087e-21, -1.253205e-20, -1.482132e-20, -8.569018e-21, 2.114149e-20, 
    -2.642798e-20, -9.438686e-21, 8.255172e-21, -2.451615e-20, 4.883892e-20, 
    -3.546583e-21, -7.275513e-21, 1.631441e-20, -2.207553e-21, 4.697204e-20, 
    1.608683e-20, 3.946639e-20, -2.429619e-20, 3.306169e-20, 2.790919e-20, 
    4.831304e-20, 4.219248e-20, 1.749453e-20, 7.305903e-20, -3.622043e-21, 
    -2.134931e-20, -3.20659e-20, 8.267608e-21, 8.739488e-21, -4.817462e-21, 
    -1.285208e-20, -1.348512e-20, 2.897396e-20, 2.248021e-20, 1.471911e-21, 
    -6.825097e-21, -4.653578e-20, 1.393493e-20, 5.11599e-21, -2.847106e-21, 
    -1.702625e-21, -3.494837e-21, -3.977259e-20, -2.415312e-20, 1.094308e-20, 
    -1.526294e-20, -3.212244e-20, -4.313849e-20, 2.560131e-21, 1.086787e-20, 
    -2.009933e-20, -1.134203e-20, -3.200145e-20, -2.583595e-20, -4.92633e-20, 
    1.604611e-20, -2.893155e-20, 1.980357e-20, 4.456102e-21, -1.732745e-20, 
    -2.195404e-20, 7.156469e-21, -1.775262e-21, -1.187157e-20, 8.040289e-21, 
    -9.844689e-21, 1.154504e-20, -5.204907e-22, 2.792983e-20, 1.812529e-20, 
    9.481378e-21, 2.606241e-20, 1.916944e-20, 3.034836e-21, 1.119163e-20, 
    -3.518784e-20, 6.474824e-21, 2.801721e-20, -2.875597e-20, -1.159678e-20, 
    1.332087e-20, 3.291554e-21, -4.354343e-21, -3.423644e-20, 2.192011e-20, 
    -3.910365e-20, -6.450772e-21, -2.739781e-22, -4.788324e-21, 2.418773e-21, 
    -7.320173e-21, 7.470608e-21, -2.793265e-20, 6.060338e-21, -3.561643e-20, 
    6.792651e-24, -2.540331e-21, -2.823605e-20, -2.726599e-20, 8.227249e-22, 
    -2.099332e-20, 2.187234e-20, 9.132484e-21, 1.334538e-22, -2.002297e-21, 
    -4.411148e-21, -2.952726e-20, -4.055546e-20, 8.451956e-21, -1.441531e-20, 
    4.875135e-21, 2.573869e-20, 6.9775e-21, 2.800985e-20, -3.392515e-20, 
    7.095417e-21, 2.212356e-21, 1.269091e-20, 8.423407e-21, -7.807606e-21, 
    1.318742e-20, 1.1886e-20, 5.266703e-21, -1.181531e-20, -4.565257e-21, 
    1.481085e-20, -4.503323e-21, 2.405755e-20, 1.237483e-20, 1.676622e-20, 
    3.76683e-21, 2.880942e-20, 1.228692e-20, -1.48643e-20, -2.014119e-20, 
    -2.024694e-20, -1.9088e-20, -1.709956e-20, -1.166151e-20, 2.279671e-21, 
    -1.82135e-21, 1.829861e-20, 1.163152e-20, -5.667989e-20, -3.350105e-20, 
    -8.693972e-21, 3.667442e-20, 1.81957e-20, 1.681087e-20, -4.191757e-21, 
    1.848181e-20, -8.890201e-21, -1.082856e-21, 2.795075e-20, -2.432502e-20, 
    3.732606e-21, -3.064235e-21, -4.084329e-20, 1.053681e-20, 3.524407e-20, 
    1.778235e-20, 1.737184e-20, 1.72689e-20, -4.452722e-21, -3.044983e-20, 
    4.308537e-20, 1.862037e-20, -5.980598e-21, 7.495494e-21, 2.387888e-20, 
    1.123261e-20, -7.753893e-21, -9.464968e-21, -5.211855e-21, 1.993194e-20, 
    4.566402e-21, 3.266926e-20, -1.093434e-20, 4.975775e-21, -8.583618e-22, 
    -2.750235e-20, -4.369858e-20, 1.892617e-21, 4.343614e-21, -2.855294e-21, 
    -7.621583e-21, -2.473554e-20, -2.357132e-21, -3.0563e-22, -5.500471e-20, 
    2.411214e-20, 1.339606e-20, -1.740066e-20, -9.765806e-21, 3.521151e-21, 
    -1.455753e-20, 6.114052e-21, 1.260119e-21, -2.181043e-20, 7.387552e-22, 
    1.060213e-20, -2.900167e-20, 1.992392e-21, 1.677271e-20, 4.344752e-20, 
    -2.235524e-20, 1.682276e-20, 1.231293e-20, -8.966806e-21, -3.79983e-22, 
    -3.384513e-20, -2.771618e-21, 8.865576e-21, -4.083499e-21, -2.716365e-20, 
    -4.758869e-20, -2.087401e-21, 1.109237e-20, -1.039434e-20, -2.410846e-21, 
    2.465666e-20, -2.594904e-20, 2.204055e-20, 1.30401e-20, 1.697523e-21, 
    -1.569156e-20, 4.769375e-21, 4.365078e-21, 1.771732e-20, -2.447457e-20, 
    3.548979e-20, -1.877077e-20, 6.269541e-21, 1.997379e-20, 2.351275e-20, 
    1.84626e-20, -3.149309e-20, -7.343637e-21, 7.656059e-21, 2.822362e-20, 
    3.709173e-20, -7.373909e-21, 3.145943e-21, 3.297202e-21, 1.242543e-20, 
    -2.319667e-20, -4.902608e-20, -2.63802e-20, 3.33956e-20, -3.572298e-21, 
    -1.84134e-20, -7.589904e-21, -3.493441e-21, -3.654776e-20, -2.411157e-20, 
    9.620767e-21, 2.180333e-20, -3.356664e-20, -8.467769e-22, 1.879563e-20, 
    1.125747e-20, 1.638059e-20, -3.233817e-20, 2.503288e-21, 3.801342e-20, 
    -4.111193e-21, 2.54582e-20, 1.087637e-20, 1.80405e-20, -7.746555e-21, 
    -3.265005e-20, -1.408169e-20, -1.350293e-20, 1.306952e-20, 1.568563e-20, 
    -9.336911e-21, -5.848573e-21, -4.842322e-21, 1.049977e-20, 3.400064e-20, 
    -6.536996e-22, 5.834709e-21, 9.168409e-21, -1.332113e-20, 2.968785e-20, 
    -4.459514e-21, -2.467109e-20, 6.009426e-21 ;

 M_SOIL2C_TO_LEACHING =
  3.710925e-20, -1.018198e-20, -1.205396e-20, 4.096007e-20, 3.385729e-20, 
    2.868616e-20, -1.995458e-20, -9.666456e-22, 1.988956e-20, 6.2853e-22, 
    -5.238714e-21, -3.627324e-20, -1.232817e-20, -7.409246e-21, 
    -3.541399e-20, 1.774334e-20, -3.824555e-20, 2.986343e-20, 2.937234e-20, 
    -3.816469e-20, 4.033802e-20, 1.958984e-20, 1.100755e-20, 3.064744e-20, 
    -9.411827e-21, 1.907755e-20, -4.278284e-21, -1.226881e-20, -2.711756e-20, 
    1.737464e-20, -4.435706e-20, 6.882518e-21, 2.827584e-21, 1.625051e-20, 
    7.33602e-21, 2.660694e-20, 7.056695e-21, 2.211293e-20, -1.75344e-20, 
    3.127766e-20, 7.814971e-21, 5.55679e-21, -1.616117e-20, 9.893039e-21, 
    2.324556e-20, 1.646002e-20, -2.904468e-21, 2.580341e-20, 3.436367e-20, 
    -4.282298e-20, 6.924637e-21, 6.896381e-21, 2.668921e-20, 1.041158e-20, 
    8.105848e-22, -7.704409e-21, -1.711681e-20, -2.096845e-20, 1.501074e-20, 
    -6.331492e-21, 2.5042e-20, -5.586905e-22, -9.326722e-21, 2.007981e-20, 
    -1.517841e-20, -2.930051e-20, -3.003729e-21, 1.096317e-20, 8.768316e-21, 
    -6.78808e-21, 1.795282e-20, 2.886256e-20, -3.663055e-21, 2.432813e-20, 
    -2.820324e-20, 2.245081e-20, 2.378981e-20, -1.564266e-20, -6.989967e-21, 
    1.135334e-20, -1.716316e-20, -3.660599e-20, 1.206244e-20, 4.57091e-20, 
    4.663022e-20, 2.541466e-21, -2.094328e-20, 1.505815e-21, 7.650721e-21, 
    6.977705e-22, 2.390432e-20, 1.033111e-21, 2.699059e-20, 8.563343e-21, 
    2.567027e-20, 4.940748e-20, -2.689786e-20, 2.527077e-20, 9.630957e-21, 
    1.259849e-20, -2.37375e-20, 1.24571e-21, -1.792627e-20, 1.883919e-20, 
    -4.72019e-20, 3.031184e-20, -1.812897e-20, -1.974421e-20, 1.213567e-20, 
    -1.18945e-21, 1.078223e-20, -8.494364e-21, -2.279546e-20, -2.645219e-21, 
    2.807377e-20, 1.614394e-20, -2.918857e-20, 2.117796e-20, 6.740286e-22, 
    6.252046e-21, 1.472745e-20, -3.516594e-21, 1.80207e-20, -4.071664e-20, 
    -8.982359e-21, 1.027436e-21, 2.018923e-20, -5.522303e-21, -1.028597e-21, 
    2.633693e-20, -3.536992e-20, 6.203697e-21, 1.770404e-20, 3.132318e-20, 
    -8.61112e-21, 1.80419e-20, -5.642466e-21, 2.618396e-20, 3.409676e-20, 
    -1.715043e-20, 1.534669e-21, 3.705611e-20, 4.604536e-21, 1.764522e-20, 
    2.991971e-20, 1.289592e-20, -1.82558e-21, -1.05682e-20, 2.069758e-20, 
    -4.081221e-21, -8.893008e-21, 3.676068e-21, 1.853612e-20, -1.384842e-20, 
    1.251168e-20, -3.032911e-20, -3.714519e-20, 2.220454e-20, 3.161497e-21, 
    1.50468e-21, -7.764343e-21, 2.296878e-20, 3.238426e-20, 6.248078e-21, 
    2.313163e-20, -2.417639e-21, -2.640563e-20, -1.005135e-20, -1.245138e-21, 
    -2.083189e-20, -1.516286e-20, 3.901134e-21, -1.801476e-20, 3.860957e-21, 
    1.7354e-20, 3.495682e-20, -3.105545e-20, 2.306151e-20, 9.468937e-21, 
    -1.012684e-20, 1.926237e-21, 2.145842e-20, -9.252924e-21, -5.041569e-20, 
    -3.305293e-20, -9.439536e-21, 4.42898e-21, -4.162645e-21, 1.158942e-20, 
    2.316525e-20, 3.286468e-21, 2.362046e-20, 2.437111e-20, 2.006286e-20, 
    8.023912e-21, -9.491241e-22, 3.02214e-20, -1.229116e-20, -1.31071e-20, 
    -2.503723e-20, -1.732178e-20, 3.036613e-20, 1.310428e-20, -1.815131e-20, 
    -9.168676e-21, -1.152979e-21, -7.886507e-21, 8.838749e-21, 5.689099e-21, 
    1.941791e-21, 1.925481e-20, -4.038668e-20, 3.874684e-20, 5.790329e-21, 
    1.720728e-20, -3.400572e-20, -5.645314e-20, 1.695545e-21, 1.120433e-20, 
    6.849721e-21, 1.608709e-20, 2.038972e-20, -5.580531e-21, -9.423983e-21, 
    -6.656388e-20, 3.468271e-21, -2.441324e-20, 4.81858e-21, 3.548011e-21, 
    -2.873126e-21, 1.097305e-20, 1.996474e-20, 1.90931e-20, -5.537578e-21, 
    -2.59168e-20, -5.47904e-21, -1.095555e-20, 2.10182e-20, 3.069579e-20, 
    1.064398e-20, 3.522547e-21, -2.117457e-20, 1.121328e-21, 3.521158e-20, 
    -6.547461e-21, -1.431805e-20, -1.368361e-20, 5.568374e-21, 3.319711e-20, 
    -1.812135e-20, 7.982355e-21, 1.221227e-20, 1.428046e-20, 1.259396e-20, 
    -1.066998e-20, 3.052475e-20, 2.275134e-20, 1.351677e-20, 2.97068e-20, 
    3.483923e-20, 3.10492e-20, -4.781815e-21, -3.633826e-20, -2.136313e-21, 
    3.166528e-22, -3.25347e-20, 1.703681e-20, 2.254636e-20, 2.434226e-20, 
    -3.916089e-21, -4.224028e-20, 1.177179e-20, -5.094526e-21, -1.470622e-20, 
    8.051596e-21, 1.667544e-20, 4.052655e-21, -5.222037e-20, -1.644586e-20, 
    3.01196e-20, 2.184463e-20, -1.225893e-20, -1.453915e-20, -1.415464e-20, 
    -4.256512e-20, -1.987427e-20, 2.151582e-20, -3.591358e-20, 2.414548e-20, 
    -3.291639e-20, -4.572901e-21, -2.575903e-20, -9.899832e-21, 3.880255e-20, 
    4.148227e-20, -1.99441e-20, 5.519764e-21, -3.32266e-21, 4.59115e-20, 
    -9.466112e-21, 2.881298e-21, 1.977675e-20, 1.480038e-20, 2.150789e-20, 
    -1.650723e-20, 2.173069e-20, -1.204489e-20, -8.133875e-21, -6.167226e-21, 
    -6.891823e-21, 3.246315e-20, 6.544947e-21, -2.43222e-20, 1.625844e-20, 
    -1.531215e-20, 2.424121e-21, -9.16044e-22, -1.399687e-20, -2.097947e-20, 
    4.086478e-20, -2.074621e-20, 1.431465e-20, 2.424953e-20, 4.508933e-20, 
    -4.976347e-21, -7.545524e-21, -4.49553e-20, -1.560816e-20, 2.189637e-20, 
    3.726674e-20, 1.040421e-20, 1.725197e-20, 2.344433e-20, -6.114052e-21, 
    4.070701e-20, 3.464527e-20, -8.433858e-21, -1.94179e-21 ;

 M_SOIL3C_TO_LEACHING =
  8.839893e-21, 9.766379e-21, 2.357777e-20, 7.557365e-22, 4.385269e-20, 
    2.37966e-20, -8.846759e-22, -2.683653e-20, 6.525998e-21, -5.498747e-20, 
    -3.910704e-20, -5.818008e-20, 2.674066e-20, 2.518453e-20, 1.165332e-20, 
    -5.764586e-21, -4.552844e-20, -3.782089e-21, -4.497396e-21, 5.023195e-20, 
    3.286887e-20, 5.117371e-23, -1.480859e-20, 2.913797e-20, -5.516141e-22, 
    1.451315e-20, 9.465563e-21, 4.637938e-21, 2.84823e-20, 1.81564e-20, 
    7.871509e-21, 3.918562e-20, -2.405162e-20, -1.185263e-20, -4.252541e-21, 
    -7.651528e-21, 2.408272e-20, -1.051712e-22, -3.163079e-20, 2.745372e-20, 
    -1.990651e-20, -2.537931e-20, -8.051334e-21, 6.042533e-21, 7.10644e-21, 
    2.720445e-21, 7.629493e-21, -1.877315e-21, 1.97216e-20, 2.061051e-20, 
    6.106563e-20, 1.614099e-21, -3.717935e-21, -8.231709e-21, 1.260894e-20, 
    1.310034e-20, 1.165614e-20, 1.276785e-20, -1.446957e-20, 3.722858e-20, 
    -1.549817e-20, -6.973825e-21, -6.513841e-21, -4.564546e-20, 1.857965e-20, 
    -2.819448e-20, -3.932214e-21, -1.862234e-20, -7.321601e-21, 2.739915e-20, 
    -3.098166e-21, 2.820124e-20, -2.429846e-20, -1.542551e-20, 4.143279e-20, 
    -8.985445e-21, 6.9795e-21, -1.674605e-21, 1.213486e-21, -2.070298e-20, 
    -3.014672e-20, 1.608683e-20, 3.139217e-20, -1.259567e-20, -5.575167e-21, 
    2.074398e-20, -2.305868e-20, -1.603452e-20, -1.534437e-20, -2.213188e-20, 
    2.994967e-20, -2.715149e-20, -8.281193e-21, -4.376812e-20, -1.413203e-20, 
    -4.162927e-20, 2.149601e-20, 2.009648e-20, -2.356758e-20, -1.396406e-21, 
    1.500167e-21, -1.008897e-20, 3.301191e-20, 3.146515e-21, -1.286397e-20, 
    6.216399e-21, 1.630224e-21, 3.511432e-20, -1.716544e-20, -3.526237e-21, 
    -1.226926e-22, 1.492196e-20, -2.331596e-20, -1.111684e-21, 3.894531e-20, 
    -1.753243e-20, 4.163763e-21, 5.21694e-21, 1.553096e-20, -2.787535e-22, 
    -3.432548e-20, 1.902692e-20, 2.777434e-20, 1.231553e-21, 6.021877e-21, 
    -1.907866e-20, -2.123619e-20, -4.323604e-20, -8.823736e-21, 2.793654e-21, 
    -2.038828e-20, -7.178541e-22, -7.938798e-21, -1.286172e-20, 2.208919e-20, 
    -1.569918e-20, -3.831011e-21, -8.903476e-21, 2.190796e-20, -1.051985e-20, 
    4.036322e-20, -1.245372e-20, 4.124484e-21, -2.110247e-20, 1.630225e-20, 
    -1.237654e-20, -5.341929e-21, -1.159818e-20, -2.358344e-20, 
    -6.880828e-21, 3.132884e-20, 3.362292e-20, -1.34235e-20, -1.167737e-20, 
    5.903143e-21, -2.788205e-20, 2.219409e-20, 2.163624e-20, -1.420355e-20, 
    2.930673e-20, 1.45547e-20, 1.60543e-20, -1.665172e-20, 7.025016e-21, 
    1.067872e-20, 1.23262e-20, 1.467203e-20, -1.846966e-20, -9.90802e-21, 
    -1.16343e-21, -3.560994e-20, -1.764411e-20, -2.754052e-20, 8.4217e-21, 
    1.607495e-20, -1.262053e-20, 7.289377e-21, -9.119471e-21, 7.025588e-21, 
    -1.236325e-20, 9.866752e-21, 5.876871e-20, -2.970001e-20, -6.602881e-21, 
    -2.778422e-20, -2.903617e-20, -4.017566e-22, -1.221227e-20, 5.304602e-21, 
    1.237766e-20, 9.288251e-21, 9.404755e-21, -2.152515e-20, 1.317835e-20, 
    -1.703056e-20, -4.222007e-21, 5.570937e-21, -2.262128e-20, 1.473707e-20, 
    4.900487e-20, 1.538593e-20, -1.28829e-20, -1.327252e-20, -2.271456e-21, 
    -3.545642e-20, -3.563877e-20, -2.547657e-20, -5.267924e-20, 1.008303e-20, 
    -3.385786e-20, -1.049722e-20, 1.25705e-20, -3.460334e-21, -5.15446e-21, 
    -1.26505e-20, -2.144287e-20, -5.085193e-21, 3.660996e-20, -2.864033e-20, 
    3.525993e-20, 7.792053e-21, 4.826638e-20, 1.219221e-20, 9.855953e-22, 
    3.751669e-20, -1.652109e-20, 5.749605e-21, 1.559233e-20, 1.555308e-21, 
    4.797376e-20, -3.481688e-20, 1.124111e-20, -4.08823e-20, 2.338438e-20, 
    -2.114685e-20, -1.111867e-20, 2.703162e-20, -2.751026e-20, -1.154164e-20, 
    -9.719718e-21, 1.288689e-20, -1.759405e-20, -2.037191e-20, 3.348126e-20, 
    -3.508607e-20, -1.234997e-20, -5.952888e-21, -7.360879e-21, 1.800571e-20, 
    7.809034e-21, -9.535974e-21, 3.232741e-20, -2.413417e-20, -1.404612e-21, 
    1.370425e-20, -5.675252e-21, -5.59072e-21, -2.773846e-20, -1.436414e-20, 
    -8.213894e-21, -1.678178e-20, -5.573477e-21, 1.416256e-20, -3.155333e-20, 
    2.828721e-20, -4.877982e-20, 3.809521e-21, -4.173951e-21, -1.014919e-20, 
    -2.055722e-21, -1.849737e-20, -1.073924e-20, 3.273542e-20, 4.608775e-23, 
    -1.102282e-20, -9.391733e-21, -2.44307e-21, -2.558656e-20, 5.145389e-21, 
    5.49968e-21, -1.855761e-20, 1.180064e-20, -1.10231e-20, 1.649874e-20, 
    -1.30093e-20, 7.580288e-21, 1.91406e-20, -9.85595e-22, 2.039281e-20, 
    8.848344e-21, 3.065353e-21, -4.617827e-21, 1.98845e-21, -1.011696e-20, 
    2.128397e-20, 1.896049e-20, -2.768501e-20, 2.305275e-20, 5.043917e-20, 
    -3.068648e-20, -2.687751e-20, -2.968163e-20, -4.687405e-21, 7.113232e-21, 
    -3.874091e-20, -2.189834e-20, -1.200164e-20, 3.449427e-20, -1.985166e-20, 
    3.803803e-20, 9.254631e-21, 1.753072e-20, -1.109519e-20, 1.190438e-20, 
    6.928605e-21, -2.540731e-20, -1.815837e-20, -1.85951e-21, 5.373591e-21, 
    9.063866e-20, -5.063825e-22, -1.763986e-20, 8.008359e-21, -2.263261e-20, 
    -5.963649e-21, -1.543062e-20, -1.207234e-20, 3.919411e-20, -8.852302e-21, 
    1.282325e-20, 2.37769e-22, -1.881855e-20, -1.382922e-20, -5.034276e-20, 
    -2.236146e-20, 1.895768e-20, 1.130922e-20, -2.108464e-20 ;

 NBP =
  -6.35703e-08, -6.384985e-08, -6.379551e-08, -6.402099e-08, -6.389591e-08, 
    -6.404356e-08, -6.362697e-08, -6.386096e-08, -6.371158e-08, 
    -6.359546e-08, -6.445858e-08, -6.403105e-08, -6.490264e-08, 
    -6.462999e-08, -6.531489e-08, -6.486022e-08, -6.540657e-08, 
    -6.530176e-08, -6.561717e-08, -6.552681e-08, -6.593026e-08, 
    -6.565888e-08, -6.613939e-08, -6.586544e-08, -6.59083e-08, -6.564993e-08, 
    -6.411708e-08, -6.440536e-08, -6.410001e-08, -6.414111e-08, 
    -6.412267e-08, -6.38985e-08, -6.378554e-08, -6.354892e-08, -6.359188e-08, 
    -6.376565e-08, -6.41596e-08, -6.402587e-08, -6.436288e-08, -6.435527e-08, 
    -6.473046e-08, -6.45613e-08, -6.519191e-08, -6.501268e-08, -6.553059e-08, 
    -6.540034e-08, -6.552447e-08, -6.548683e-08, -6.552496e-08, 
    -6.533394e-08, -6.541578e-08, -6.524769e-08, -6.459298e-08, -6.47854e-08, 
    -6.421152e-08, -6.386645e-08, -6.363724e-08, -6.347459e-08, 
    -6.349758e-08, -6.354141e-08, -6.376668e-08, -6.397845e-08, 
    -6.413985e-08, -6.424781e-08, -6.435418e-08, -6.467617e-08, 
    -6.484658e-08, -6.522815e-08, -6.515928e-08, -6.527594e-08, 
    -6.538738e-08, -6.557449e-08, -6.554369e-08, -6.562612e-08, 
    -6.527286e-08, -6.550764e-08, -6.512006e-08, -6.522607e-08, 
    -6.438312e-08, -6.406194e-08, -6.392545e-08, -6.380596e-08, 
    -6.351526e-08, -6.371601e-08, -6.363688e-08, -6.382514e-08, 
    -6.394477e-08, -6.38856e-08, -6.425076e-08, -6.41088e-08, -6.485669e-08, 
    -6.453455e-08, -6.537438e-08, -6.517342e-08, -6.542255e-08, 
    -6.529542e-08, -6.551326e-08, -6.531721e-08, -6.565681e-08, 
    -6.573075e-08, -6.568022e-08, -6.587433e-08, -6.530634e-08, 
    -6.552447e-08, -6.388395e-08, -6.389359e-08, -6.393855e-08, 
    -6.374094e-08, -6.372885e-08, -6.354775e-08, -6.370889e-08, 
    -6.377751e-08, -6.39517e-08, -6.405474e-08, -6.415268e-08, -6.436803e-08, 
    -6.460854e-08, -6.494484e-08, -6.518644e-08, -6.53484e-08, -6.524908e-08, 
    -6.533676e-08, -6.523875e-08, -6.519281e-08, -6.570305e-08, 
    -6.541654e-08, -6.584641e-08, -6.582263e-08, -6.562809e-08, -6.58253e-08, 
    -6.390037e-08, -6.384484e-08, -6.365205e-08, -6.380292e-08, 
    -6.352803e-08, -6.36819e-08, -6.377039e-08, -6.411177e-08, -6.418676e-08, 
    -6.425632e-08, -6.439367e-08, -6.456996e-08, -6.48792e-08, -6.514825e-08, 
    -6.539386e-08, -6.537586e-08, -6.53822e-08, -6.543707e-08, -6.530116e-08, 
    -6.545939e-08, -6.548594e-08, -6.541651e-08, -6.581944e-08, 
    -6.570433e-08, -6.582212e-08, -6.574717e-08, -6.386289e-08, 
    -6.395633e-08, -6.390584e-08, -6.400078e-08, -6.39339e-08, -6.423132e-08, 
    -6.432049e-08, -6.473773e-08, -6.456649e-08, -6.483902e-08, 
    -6.459417e-08, -6.463756e-08, -6.484792e-08, -6.46074e-08, -6.513343e-08, 
    -6.477681e-08, -6.543921e-08, -6.508311e-08, -6.546152e-08, -6.53928e-08, 
    -6.550658e-08, -6.560848e-08, -6.573668e-08, -6.597322e-08, 
    -6.591844e-08, -6.611626e-08, -6.409562e-08, -6.421681e-08, 
    -6.420614e-08, -6.433297e-08, -6.442676e-08, -6.463005e-08, -6.49561e-08, 
    -6.483349e-08, -6.505858e-08, -6.510377e-08, -6.47618e-08, -6.497177e-08, 
    -6.429792e-08, -6.44068e-08, -6.434197e-08, -6.410518e-08, -6.486175e-08, 
    -6.447348e-08, -6.519043e-08, -6.498011e-08, -6.559395e-08, 
    -6.528868e-08, -6.588829e-08, -6.614464e-08, -6.638587e-08, -6.66678e-08, 
    -6.428295e-08, -6.42006e-08, -6.434804e-08, -6.455205e-08, -6.474131e-08, 
    -6.499293e-08, -6.501867e-08, -6.506582e-08, -6.518791e-08, 
    -6.529058e-08, -6.508073e-08, -6.531631e-08, -6.443206e-08, 
    -6.489545e-08, -6.416948e-08, -6.438809e-08, -6.454002e-08, 
    -6.447337e-08, -6.481947e-08, -6.490105e-08, -6.523254e-08, 
    -6.506118e-08, -6.608137e-08, -6.563001e-08, -6.688245e-08, 
    -6.653246e-08, -6.417183e-08, -6.428267e-08, -6.466841e-08, 
    -6.448487e-08, -6.500973e-08, -6.513893e-08, -6.524394e-08, -6.53782e-08, 
    -6.539269e-08, -6.547224e-08, -6.534189e-08, -6.546708e-08, 
    -6.499347e-08, -6.520511e-08, -6.462431e-08, -6.476568e-08, 
    -6.470064e-08, -6.46293e-08, -6.484947e-08, -6.508403e-08, -6.508903e-08, 
    -6.516425e-08, -6.537621e-08, -6.501185e-08, -6.613964e-08, 
    -6.544317e-08, -6.440352e-08, -6.461701e-08, -6.464749e-08, 
    -6.456479e-08, -6.512597e-08, -6.492264e-08, -6.54703e-08, -6.532228e-08, 
    -6.55648e-08, -6.544429e-08, -6.542655e-08, -6.527178e-08, -6.517542e-08, 
    -6.493197e-08, -6.473388e-08, -6.457679e-08, -6.461332e-08, 
    -6.478587e-08, -6.509838e-08, -6.5394e-08, -6.532925e-08, -6.554637e-08, 
    -6.497167e-08, -6.521266e-08, -6.511952e-08, -6.536237e-08, 
    -6.483023e-08, -6.528341e-08, -6.471441e-08, -6.476429e-08, -6.49186e-08, 
    -6.522901e-08, -6.529767e-08, -6.5371e-08, -6.532575e-08, -6.510631e-08, 
    -6.507035e-08, -6.491485e-08, -6.487192e-08, -6.475343e-08, 
    -6.465533e-08, -6.474496e-08, -6.483909e-08, -6.51064e-08, -6.534729e-08, 
    -6.560993e-08, -6.56742e-08, -6.598109e-08, -6.573129e-08, -6.614352e-08, 
    -6.579306e-08, -6.639972e-08, -6.530966e-08, -6.578274e-08, 
    -6.492562e-08, -6.501796e-08, -6.518498e-08, -6.556804e-08, 
    -6.536123e-08, -6.560308e-08, -6.506895e-08, -6.479183e-08, 
    -6.472012e-08, -6.458635e-08, -6.472317e-08, -6.471205e-08, 
    -6.484298e-08, -6.480091e-08, -6.511527e-08, -6.494641e-08, 
    -6.542611e-08, -6.560117e-08, -6.609553e-08, -6.639859e-08, 
    -6.670707e-08, -6.684326e-08, -6.688472e-08, -6.690204e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.35703e-08, 6.384985e-08, 6.379551e-08, 6.402099e-08, 6.389591e-08, 
    6.404356e-08, 6.362697e-08, 6.386096e-08, 6.371158e-08, 6.359546e-08, 
    6.445858e-08, 6.403105e-08, 6.490264e-08, 6.462999e-08, 6.531489e-08, 
    6.486022e-08, 6.540657e-08, 6.530176e-08, 6.561717e-08, 6.552681e-08, 
    6.593026e-08, 6.565888e-08, 6.613939e-08, 6.586544e-08, 6.59083e-08, 
    6.564993e-08, 6.411708e-08, 6.440536e-08, 6.410001e-08, 6.414111e-08, 
    6.412267e-08, 6.38985e-08, 6.378554e-08, 6.354892e-08, 6.359188e-08, 
    6.376565e-08, 6.41596e-08, 6.402587e-08, 6.436288e-08, 6.435527e-08, 
    6.473046e-08, 6.45613e-08, 6.519191e-08, 6.501268e-08, 6.553059e-08, 
    6.540034e-08, 6.552447e-08, 6.548683e-08, 6.552496e-08, 6.533394e-08, 
    6.541578e-08, 6.524769e-08, 6.459298e-08, 6.47854e-08, 6.421152e-08, 
    6.386645e-08, 6.363724e-08, 6.347459e-08, 6.349758e-08, 6.354141e-08, 
    6.376668e-08, 6.397845e-08, 6.413985e-08, 6.424781e-08, 6.435418e-08, 
    6.467617e-08, 6.484658e-08, 6.522815e-08, 6.515928e-08, 6.527594e-08, 
    6.538738e-08, 6.557449e-08, 6.554369e-08, 6.562612e-08, 6.527286e-08, 
    6.550764e-08, 6.512006e-08, 6.522607e-08, 6.438312e-08, 6.406194e-08, 
    6.392545e-08, 6.380596e-08, 6.351526e-08, 6.371601e-08, 6.363688e-08, 
    6.382514e-08, 6.394477e-08, 6.38856e-08, 6.425076e-08, 6.41088e-08, 
    6.485669e-08, 6.453455e-08, 6.537438e-08, 6.517342e-08, 6.542255e-08, 
    6.529542e-08, 6.551326e-08, 6.531721e-08, 6.565681e-08, 6.573075e-08, 
    6.568022e-08, 6.587433e-08, 6.530634e-08, 6.552447e-08, 6.388395e-08, 
    6.389359e-08, 6.393855e-08, 6.374094e-08, 6.372885e-08, 6.354775e-08, 
    6.370889e-08, 6.377751e-08, 6.39517e-08, 6.405474e-08, 6.415268e-08, 
    6.436803e-08, 6.460854e-08, 6.494484e-08, 6.518644e-08, 6.53484e-08, 
    6.524908e-08, 6.533676e-08, 6.523875e-08, 6.519281e-08, 6.570305e-08, 
    6.541654e-08, 6.584641e-08, 6.582263e-08, 6.562809e-08, 6.58253e-08, 
    6.390037e-08, 6.384484e-08, 6.365205e-08, 6.380292e-08, 6.352803e-08, 
    6.36819e-08, 6.377039e-08, 6.411177e-08, 6.418676e-08, 6.425632e-08, 
    6.439367e-08, 6.456996e-08, 6.48792e-08, 6.514825e-08, 6.539386e-08, 
    6.537586e-08, 6.53822e-08, 6.543707e-08, 6.530116e-08, 6.545939e-08, 
    6.548594e-08, 6.541651e-08, 6.581944e-08, 6.570433e-08, 6.582212e-08, 
    6.574717e-08, 6.386289e-08, 6.395633e-08, 6.390584e-08, 6.400078e-08, 
    6.39339e-08, 6.423132e-08, 6.432049e-08, 6.473773e-08, 6.456649e-08, 
    6.483902e-08, 6.459417e-08, 6.463756e-08, 6.484792e-08, 6.46074e-08, 
    6.513343e-08, 6.477681e-08, 6.543921e-08, 6.508311e-08, 6.546152e-08, 
    6.53928e-08, 6.550658e-08, 6.560848e-08, 6.573668e-08, 6.597322e-08, 
    6.591844e-08, 6.611626e-08, 6.409562e-08, 6.421681e-08, 6.420614e-08, 
    6.433297e-08, 6.442676e-08, 6.463005e-08, 6.49561e-08, 6.483349e-08, 
    6.505858e-08, 6.510377e-08, 6.47618e-08, 6.497177e-08, 6.429792e-08, 
    6.44068e-08, 6.434197e-08, 6.410518e-08, 6.486175e-08, 6.447348e-08, 
    6.519043e-08, 6.498011e-08, 6.559395e-08, 6.528868e-08, 6.588829e-08, 
    6.614464e-08, 6.638587e-08, 6.66678e-08, 6.428295e-08, 6.42006e-08, 
    6.434804e-08, 6.455205e-08, 6.474131e-08, 6.499293e-08, 6.501867e-08, 
    6.506582e-08, 6.518791e-08, 6.529058e-08, 6.508073e-08, 6.531631e-08, 
    6.443206e-08, 6.489545e-08, 6.416948e-08, 6.438809e-08, 6.454002e-08, 
    6.447337e-08, 6.481947e-08, 6.490105e-08, 6.523254e-08, 6.506118e-08, 
    6.608137e-08, 6.563001e-08, 6.688245e-08, 6.653246e-08, 6.417183e-08, 
    6.428267e-08, 6.466841e-08, 6.448487e-08, 6.500973e-08, 6.513893e-08, 
    6.524394e-08, 6.53782e-08, 6.539269e-08, 6.547224e-08, 6.534189e-08, 
    6.546708e-08, 6.499347e-08, 6.520511e-08, 6.462431e-08, 6.476568e-08, 
    6.470064e-08, 6.46293e-08, 6.484947e-08, 6.508403e-08, 6.508903e-08, 
    6.516425e-08, 6.537621e-08, 6.501185e-08, 6.613964e-08, 6.544317e-08, 
    6.440352e-08, 6.461701e-08, 6.464749e-08, 6.456479e-08, 6.512597e-08, 
    6.492264e-08, 6.54703e-08, 6.532228e-08, 6.55648e-08, 6.544429e-08, 
    6.542655e-08, 6.527178e-08, 6.517542e-08, 6.493197e-08, 6.473388e-08, 
    6.457679e-08, 6.461332e-08, 6.478587e-08, 6.509838e-08, 6.5394e-08, 
    6.532925e-08, 6.554637e-08, 6.497167e-08, 6.521266e-08, 6.511952e-08, 
    6.536237e-08, 6.483023e-08, 6.528341e-08, 6.471441e-08, 6.476429e-08, 
    6.49186e-08, 6.522901e-08, 6.529767e-08, 6.5371e-08, 6.532575e-08, 
    6.510631e-08, 6.507035e-08, 6.491485e-08, 6.487192e-08, 6.475343e-08, 
    6.465533e-08, 6.474496e-08, 6.483909e-08, 6.51064e-08, 6.534729e-08, 
    6.560993e-08, 6.56742e-08, 6.598109e-08, 6.573129e-08, 6.614352e-08, 
    6.579306e-08, 6.639972e-08, 6.530966e-08, 6.578274e-08, 6.492562e-08, 
    6.501796e-08, 6.518498e-08, 6.556804e-08, 6.536123e-08, 6.560308e-08, 
    6.506895e-08, 6.479183e-08, 6.472012e-08, 6.458635e-08, 6.472317e-08, 
    6.471205e-08, 6.484298e-08, 6.480091e-08, 6.511527e-08, 6.494641e-08, 
    6.542611e-08, 6.560117e-08, 6.609553e-08, 6.639859e-08, 6.670707e-08, 
    6.684326e-08, 6.688472e-08, 6.690204e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.35703e-08, -6.384985e-08, -6.379551e-08, -6.402099e-08, -6.389591e-08, 
    -6.404356e-08, -6.362697e-08, -6.386096e-08, -6.371158e-08, 
    -6.359546e-08, -6.445858e-08, -6.403105e-08, -6.490264e-08, 
    -6.462999e-08, -6.531489e-08, -6.486022e-08, -6.540657e-08, 
    -6.530176e-08, -6.561717e-08, -6.552681e-08, -6.593026e-08, 
    -6.565888e-08, -6.613939e-08, -6.586544e-08, -6.59083e-08, -6.564993e-08, 
    -6.411708e-08, -6.440536e-08, -6.410001e-08, -6.414111e-08, 
    -6.412267e-08, -6.38985e-08, -6.378554e-08, -6.354892e-08, -6.359188e-08, 
    -6.376565e-08, -6.41596e-08, -6.402587e-08, -6.436288e-08, -6.435527e-08, 
    -6.473046e-08, -6.45613e-08, -6.519191e-08, -6.501268e-08, -6.553059e-08, 
    -6.540034e-08, -6.552447e-08, -6.548683e-08, -6.552496e-08, 
    -6.533394e-08, -6.541578e-08, -6.524769e-08, -6.459298e-08, -6.47854e-08, 
    -6.421152e-08, -6.386645e-08, -6.363724e-08, -6.347459e-08, 
    -6.349758e-08, -6.354141e-08, -6.376668e-08, -6.397845e-08, 
    -6.413985e-08, -6.424781e-08, -6.435418e-08, -6.467617e-08, 
    -6.484658e-08, -6.522815e-08, -6.515928e-08, -6.527594e-08, 
    -6.538738e-08, -6.557449e-08, -6.554369e-08, -6.562612e-08, 
    -6.527286e-08, -6.550764e-08, -6.512006e-08, -6.522607e-08, 
    -6.438312e-08, -6.406194e-08, -6.392545e-08, -6.380596e-08, 
    -6.351526e-08, -6.371601e-08, -6.363688e-08, -6.382514e-08, 
    -6.394477e-08, -6.38856e-08, -6.425076e-08, -6.41088e-08, -6.485669e-08, 
    -6.453455e-08, -6.537438e-08, -6.517342e-08, -6.542255e-08, 
    -6.529542e-08, -6.551326e-08, -6.531721e-08, -6.565681e-08, 
    -6.573075e-08, -6.568022e-08, -6.587433e-08, -6.530634e-08, 
    -6.552447e-08, -6.388395e-08, -6.389359e-08, -6.393855e-08, 
    -6.374094e-08, -6.372885e-08, -6.354775e-08, -6.370889e-08, 
    -6.377751e-08, -6.39517e-08, -6.405474e-08, -6.415268e-08, -6.436803e-08, 
    -6.460854e-08, -6.494484e-08, -6.518644e-08, -6.53484e-08, -6.524908e-08, 
    -6.533676e-08, -6.523875e-08, -6.519281e-08, -6.570305e-08, 
    -6.541654e-08, -6.584641e-08, -6.582263e-08, -6.562809e-08, -6.58253e-08, 
    -6.390037e-08, -6.384484e-08, -6.365205e-08, -6.380292e-08, 
    -6.352803e-08, -6.36819e-08, -6.377039e-08, -6.411177e-08, -6.418676e-08, 
    -6.425632e-08, -6.439367e-08, -6.456996e-08, -6.48792e-08, -6.514825e-08, 
    -6.539386e-08, -6.537586e-08, -6.53822e-08, -6.543707e-08, -6.530116e-08, 
    -6.545939e-08, -6.548594e-08, -6.541651e-08, -6.581944e-08, 
    -6.570433e-08, -6.582212e-08, -6.574717e-08, -6.386289e-08, 
    -6.395633e-08, -6.390584e-08, -6.400078e-08, -6.39339e-08, -6.423132e-08, 
    -6.432049e-08, -6.473773e-08, -6.456649e-08, -6.483902e-08, 
    -6.459417e-08, -6.463756e-08, -6.484792e-08, -6.46074e-08, -6.513343e-08, 
    -6.477681e-08, -6.543921e-08, -6.508311e-08, -6.546152e-08, -6.53928e-08, 
    -6.550658e-08, -6.560848e-08, -6.573668e-08, -6.597322e-08, 
    -6.591844e-08, -6.611626e-08, -6.409562e-08, -6.421681e-08, 
    -6.420614e-08, -6.433297e-08, -6.442676e-08, -6.463005e-08, -6.49561e-08, 
    -6.483349e-08, -6.505858e-08, -6.510377e-08, -6.47618e-08, -6.497177e-08, 
    -6.429792e-08, -6.44068e-08, -6.434197e-08, -6.410518e-08, -6.486175e-08, 
    -6.447348e-08, -6.519043e-08, -6.498011e-08, -6.559395e-08, 
    -6.528868e-08, -6.588829e-08, -6.614464e-08, -6.638587e-08, -6.66678e-08, 
    -6.428295e-08, -6.42006e-08, -6.434804e-08, -6.455205e-08, -6.474131e-08, 
    -6.499293e-08, -6.501867e-08, -6.506582e-08, -6.518791e-08, 
    -6.529058e-08, -6.508073e-08, -6.531631e-08, -6.443206e-08, 
    -6.489545e-08, -6.416948e-08, -6.438809e-08, -6.454002e-08, 
    -6.447337e-08, -6.481947e-08, -6.490105e-08, -6.523254e-08, 
    -6.506118e-08, -6.608137e-08, -6.563001e-08, -6.688245e-08, 
    -6.653246e-08, -6.417183e-08, -6.428267e-08, -6.466841e-08, 
    -6.448487e-08, -6.500973e-08, -6.513893e-08, -6.524394e-08, -6.53782e-08, 
    -6.539269e-08, -6.547224e-08, -6.534189e-08, -6.546708e-08, 
    -6.499347e-08, -6.520511e-08, -6.462431e-08, -6.476568e-08, 
    -6.470064e-08, -6.46293e-08, -6.484947e-08, -6.508403e-08, -6.508903e-08, 
    -6.516425e-08, -6.537621e-08, -6.501185e-08, -6.613964e-08, 
    -6.544317e-08, -6.440352e-08, -6.461701e-08, -6.464749e-08, 
    -6.456479e-08, -6.512597e-08, -6.492264e-08, -6.54703e-08, -6.532228e-08, 
    -6.55648e-08, -6.544429e-08, -6.542655e-08, -6.527178e-08, -6.517542e-08, 
    -6.493197e-08, -6.473388e-08, -6.457679e-08, -6.461332e-08, 
    -6.478587e-08, -6.509838e-08, -6.5394e-08, -6.532925e-08, -6.554637e-08, 
    -6.497167e-08, -6.521266e-08, -6.511952e-08, -6.536237e-08, 
    -6.483023e-08, -6.528341e-08, -6.471441e-08, -6.476429e-08, -6.49186e-08, 
    -6.522901e-08, -6.529767e-08, -6.5371e-08, -6.532575e-08, -6.510631e-08, 
    -6.507035e-08, -6.491485e-08, -6.487192e-08, -6.475343e-08, 
    -6.465533e-08, -6.474496e-08, -6.483909e-08, -6.51064e-08, -6.534729e-08, 
    -6.560993e-08, -6.56742e-08, -6.598109e-08, -6.573129e-08, -6.614352e-08, 
    -6.579306e-08, -6.639972e-08, -6.530966e-08, -6.578274e-08, 
    -6.492562e-08, -6.501796e-08, -6.518498e-08, -6.556804e-08, 
    -6.536123e-08, -6.560308e-08, -6.506895e-08, -6.479183e-08, 
    -6.472012e-08, -6.458635e-08, -6.472317e-08, -6.471205e-08, 
    -6.484298e-08, -6.480091e-08, -6.511527e-08, -6.494641e-08, 
    -6.542611e-08, -6.560117e-08, -6.609553e-08, -6.639859e-08, 
    -6.670707e-08, -6.684326e-08, -6.688472e-08, -6.690204e-08 ;

 NET_NMIN =
  8.955642e-09, 8.995023e-09, 8.987367e-09, 9.019131e-09, 9.001511e-09, 
    9.02231e-09, 8.963626e-09, 8.996587e-09, 8.975546e-09, 8.959187e-09, 
    9.080773e-09, 9.020548e-09, 9.143326e-09, 9.104919e-09, 9.201399e-09, 
    9.13735e-09, 9.214313e-09, 9.19955e-09, 9.243981e-09, 9.231252e-09, 
    9.288083e-09, 9.249855e-09, 9.317541e-09, 9.278954e-09, 9.284991e-09, 
    9.248595e-09, 9.032667e-09, 9.073275e-09, 9.030261e-09, 9.036052e-09, 
    9.033453e-09, 9.001875e-09, 8.985962e-09, 8.952632e-09, 8.958683e-09, 
    8.983163e-09, 9.038656e-09, 9.019818e-09, 9.067292e-09, 9.06622e-09, 
    9.119073e-09, 9.095243e-09, 9.184074e-09, 9.158827e-09, 9.231783e-09, 
    9.213435e-09, 9.230922e-09, 9.225619e-09, 9.230991e-09, 9.204082e-09, 
    9.215611e-09, 9.191933e-09, 9.099706e-09, 9.126811e-09, 9.04597e-09, 
    8.997361e-09, 8.965072e-09, 8.94216e-09, 8.945399e-09, 8.951574e-09, 
    8.983306e-09, 9.013139e-09, 9.035873e-09, 9.051082e-09, 9.066066e-09, 
    9.111425e-09, 9.135429e-09, 9.18918e-09, 9.179479e-09, 9.195912e-09, 
    9.21161e-09, 9.237968e-09, 9.233629e-09, 9.245241e-09, 9.195478e-09, 
    9.228551e-09, 9.173953e-09, 9.188886e-09, 9.070144e-09, 9.0249e-09, 
    9.005673e-09, 8.988839e-09, 8.94789e-09, 8.976169e-09, 8.965021e-09, 
    8.991542e-09, 9.008393e-09, 9.000058e-09, 9.051497e-09, 9.0315e-09, 
    9.136852e-09, 9.091474e-09, 9.20978e-09, 9.18147e-09, 9.216564e-09, 
    9.198656e-09, 9.229342e-09, 9.201725e-09, 9.249563e-09, 9.25998e-09, 
    9.252862e-09, 9.280205e-09, 9.200194e-09, 9.230922e-09, 8.999825e-09, 
    9.001185e-09, 9.007517e-09, 8.97968e-09, 8.977977e-09, 8.952466e-09, 
    8.975165e-09, 8.984832e-09, 9.00937e-09, 9.023885e-09, 9.037682e-09, 
    9.068017e-09, 9.101898e-09, 9.149272e-09, 9.183305e-09, 9.206119e-09, 
    9.192129e-09, 9.20448e-09, 9.190673e-09, 9.184202e-09, 9.256077e-09, 
    9.215719e-09, 9.276272e-09, 9.272921e-09, 9.245518e-09, 9.273299e-09, 
    9.002139e-09, 8.994316e-09, 8.967159e-09, 8.988412e-09, 8.949688e-09, 
    8.971364e-09, 8.983829e-09, 9.031918e-09, 9.042483e-09, 9.052281e-09, 
    9.071631e-09, 9.096462e-09, 9.140024e-09, 9.177925e-09, 9.212523e-09, 
    9.209988e-09, 9.210881e-09, 9.218611e-09, 9.199464e-09, 9.221753e-09, 
    9.225495e-09, 9.215714e-09, 9.272473e-09, 9.256257e-09, 9.27285e-09, 
    9.262292e-09, 8.996859e-09, 9.010021e-09, 9.00291e-09, 9.016284e-09, 
    9.006862e-09, 9.048759e-09, 9.061321e-09, 9.120097e-09, 9.095974e-09, 
    9.134364e-09, 9.099874e-09, 9.105985e-09, 9.135618e-09, 9.101737e-09, 
    9.175836e-09, 9.125601e-09, 9.218911e-09, 9.168748e-09, 9.222054e-09, 
    9.212374e-09, 9.228401e-09, 9.242756e-09, 9.260814e-09, 9.294135e-09, 
    9.28642e-09, 9.314284e-09, 9.029644e-09, 9.046715e-09, 9.045212e-09, 
    9.063077e-09, 9.076291e-09, 9.104927e-09, 9.150858e-09, 9.133585e-09, 
    9.165293e-09, 9.171659e-09, 9.123487e-09, 9.153064e-09, 9.058141e-09, 
    9.073478e-09, 9.064346e-09, 9.03099e-09, 9.137567e-09, 9.082872e-09, 
    9.183867e-09, 9.154238e-09, 9.24071e-09, 9.197707e-09, 9.282171e-09, 
    9.318281e-09, 9.352263e-09, 9.391978e-09, 9.056032e-09, 9.044432e-09, 
    9.065202e-09, 9.093939e-09, 9.1206e-09, 9.156046e-09, 9.159672e-09, 
    9.166313e-09, 9.183513e-09, 9.197974e-09, 9.168413e-09, 9.201599e-09, 
    9.077037e-09, 9.142314e-09, 9.040047e-09, 9.070844e-09, 9.092245e-09, 
    9.082856e-09, 9.131611e-09, 9.143103e-09, 9.189798e-09, 9.165659e-09, 
    9.30937e-09, 9.245789e-09, 9.422214e-09, 9.372912e-09, 9.040379e-09, 
    9.055992e-09, 9.11033e-09, 9.084476e-09, 9.158412e-09, 9.176611e-09, 
    9.191405e-09, 9.210317e-09, 9.212358e-09, 9.223563e-09, 9.205202e-09, 
    9.222838e-09, 9.156121e-09, 9.185936e-09, 9.104118e-09, 9.124033e-09, 
    9.114872e-09, 9.104823e-09, 9.135836e-09, 9.168879e-09, 9.169583e-09, 
    9.180178e-09, 9.210037e-09, 9.158711e-09, 9.317579e-09, 9.219469e-09, 
    9.073017e-09, 9.103091e-09, 9.107385e-09, 9.095736e-09, 9.174786e-09, 
    9.146143e-09, 9.223291e-09, 9.20244e-09, 9.236603e-09, 9.219627e-09, 
    9.217129e-09, 9.195325e-09, 9.181751e-09, 9.147457e-09, 9.119553e-09, 
    9.097425e-09, 9.10257e-09, 9.126877e-09, 9.1709e-09, 9.212544e-09, 
    9.203421e-09, 9.234006e-09, 9.153051e-09, 9.186998e-09, 9.173878e-09, 
    9.208088e-09, 9.133127e-09, 9.196964e-09, 9.11681e-09, 9.123838e-09, 
    9.145575e-09, 9.189301e-09, 9.198973e-09, 9.209303e-09, 9.202928e-09, 
    9.172017e-09, 9.166952e-09, 9.145046e-09, 9.138999e-09, 9.122307e-09, 
    9.108489e-09, 9.121115e-09, 9.134374e-09, 9.172029e-09, 9.205963e-09, 
    9.24296e-09, 9.252014e-09, 9.295244e-09, 9.260054e-09, 9.318125e-09, 
    9.268756e-09, 9.354214e-09, 9.200661e-09, 9.267302e-09, 9.146564e-09, 
    9.159571e-09, 9.183099e-09, 9.237058e-09, 9.207926e-09, 9.241996e-09, 
    9.166754e-09, 9.127716e-09, 9.117615e-09, 9.098771e-09, 9.118046e-09, 
    9.116478e-09, 9.134922e-09, 9.128995e-09, 9.17328e-09, 9.149492e-09, 
    9.217066e-09, 9.241726e-09, 9.311365e-09, 9.354055e-09, 9.397509e-09, 
    9.416694e-09, 9.422533e-09, 9.424974e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.485607e-14, 4.497747e-14, 4.495389e-14, 4.505172e-14, 4.499748e-14, 
    4.506151e-14, 4.488071e-14, 4.498227e-14, 4.491746e-14, 4.486703e-14, 
    4.524128e-14, 4.505608e-14, 4.54335e-14, 4.53156e-14, 4.561158e-14, 
    4.541514e-14, 4.565116e-14, 4.560596e-14, 4.574206e-14, 4.570309e-14, 
    4.58769e-14, 4.576004e-14, 4.596696e-14, 4.584903e-14, 4.586747e-14, 
    4.575618e-14, 4.509342e-14, 4.521822e-14, 4.508601e-14, 4.510382e-14, 
    4.509583e-14, 4.499858e-14, 4.494952e-14, 4.484682e-14, 4.486548e-14, 
    4.494092e-14, 4.511182e-14, 4.505386e-14, 4.519997e-14, 4.519667e-14, 
    4.535908e-14, 4.528588e-14, 4.555852e-14, 4.548112e-14, 4.570472e-14, 
    4.564851e-14, 4.570207e-14, 4.568584e-14, 4.570228e-14, 4.561985e-14, 
    4.565517e-14, 4.558262e-14, 4.529958e-14, 4.538283e-14, 4.513434e-14, 
    4.498462e-14, 4.488516e-14, 4.481451e-14, 4.48245e-14, 4.484354e-14, 
    4.494136e-14, 4.50333e-14, 4.51033e-14, 4.51501e-14, 4.519619e-14, 
    4.53355e-14, 4.540926e-14, 4.557415e-14, 4.554444e-14, 4.559479e-14, 
    4.564292e-14, 4.572364e-14, 4.571036e-14, 4.57459e-14, 4.559349e-14, 
    4.569479e-14, 4.552753e-14, 4.557328e-14, 4.520858e-14, 4.506951e-14, 
    4.501023e-14, 4.495842e-14, 4.483218e-14, 4.491936e-14, 4.4885e-14, 
    4.496677e-14, 4.501868e-14, 4.499301e-14, 4.515138e-14, 4.508983e-14, 
    4.541363e-14, 4.527427e-14, 4.563731e-14, 4.555054e-14, 4.56581e-14, 
    4.560324e-14, 4.569722e-14, 4.561264e-14, 4.575914e-14, 4.579099e-14, 
    4.576922e-14, 4.585288e-14, 4.560794e-14, 4.570206e-14, 4.499229e-14, 
    4.499647e-14, 4.501599e-14, 4.493019e-14, 4.492494e-14, 4.48463e-14, 
    4.491629e-14, 4.494607e-14, 4.50217e-14, 4.506638e-14, 4.510885e-14, 
    4.520218e-14, 4.53063e-14, 4.545177e-14, 4.555617e-14, 4.56261e-14, 
    4.558323e-14, 4.562108e-14, 4.557876e-14, 4.555893e-14, 4.577905e-14, 
    4.565549e-14, 4.584085e-14, 4.583061e-14, 4.574674e-14, 4.583176e-14, 
    4.499941e-14, 4.497533e-14, 4.48916e-14, 4.495713e-14, 4.483773e-14, 
    4.490456e-14, 4.494296e-14, 4.509108e-14, 4.512364e-14, 4.515377e-14, 
    4.52133e-14, 4.528963e-14, 4.54234e-14, 4.553966e-14, 4.564573e-14, 
    4.563796e-14, 4.56407e-14, 4.566436e-14, 4.560571e-14, 4.567399e-14, 
    4.568543e-14, 4.565549e-14, 4.582924e-14, 4.577963e-14, 4.583039e-14, 
    4.57981e-14, 4.498316e-14, 4.50237e-14, 4.500179e-14, 4.504297e-14, 
    4.501395e-14, 4.51429e-14, 4.518154e-14, 4.536219e-14, 4.528812e-14, 
    4.540601e-14, 4.530011e-14, 4.531887e-14, 4.54098e-14, 4.530584e-14, 
    4.553325e-14, 4.537907e-14, 4.566528e-14, 4.551147e-14, 4.567491e-14, 
    4.564527e-14, 4.569436e-14, 4.57383e-14, 4.579357e-14, 4.589544e-14, 
    4.587187e-14, 4.595703e-14, 4.508411e-14, 4.513663e-14, 4.513204e-14, 
    4.5187e-14, 4.522762e-14, 4.531564e-14, 4.545666e-14, 4.540366e-14, 
    4.550097e-14, 4.552048e-14, 4.537265e-14, 4.546342e-14, 4.517179e-14, 
    4.521893e-14, 4.519088e-14, 4.508824e-14, 4.541584e-14, 4.524782e-14, 
    4.555789e-14, 4.546704e-14, 4.573203e-14, 4.560028e-14, 4.585888e-14, 
    4.596918e-14, 4.607301e-14, 4.619408e-14, 4.516532e-14, 4.512964e-14, 
    4.519354e-14, 4.528184e-14, 4.536377e-14, 4.547258e-14, 4.548372e-14, 
    4.550408e-14, 4.555682e-14, 4.560114e-14, 4.551049e-14, 4.561226e-14, 
    4.52298e-14, 4.543042e-14, 4.511612e-14, 4.521082e-14, 4.527664e-14, 
    4.52478e-14, 4.53976e-14, 4.543288e-14, 4.557605e-14, 4.550209e-14, 
    4.594194e-14, 4.574753e-14, 4.628626e-14, 4.613596e-14, 4.511717e-14, 
    4.516521e-14, 4.533221e-14, 4.525279e-14, 4.547985e-14, 4.553566e-14, 
    4.558101e-14, 4.563894e-14, 4.564522e-14, 4.567953e-14, 4.56233e-14, 
    4.567732e-14, 4.547281e-14, 4.556424e-14, 4.531317e-14, 4.537431e-14, 
    4.53462e-14, 4.531533e-14, 4.541057e-14, 4.551191e-14, 4.551412e-14, 
    4.554656e-14, 4.563793e-14, 4.548077e-14, 4.596693e-14, 4.566685e-14, 
    4.521757e-14, 4.530994e-14, 4.532318e-14, 4.528741e-14, 4.553007e-14, 
    4.54422e-14, 4.56787e-14, 4.561483e-14, 4.571947e-14, 4.566748e-14, 
    4.565983e-14, 4.559303e-14, 4.555141e-14, 4.544622e-14, 4.536055e-14, 
    4.52926e-14, 4.530841e-14, 4.538304e-14, 4.551812e-14, 4.564577e-14, 
    4.56178e-14, 4.571152e-14, 4.54634e-14, 4.556747e-14, 4.552726e-14, 
    4.563213e-14, 4.540224e-14, 4.55979e-14, 4.535215e-14, 4.537373e-14, 
    4.544045e-14, 4.55745e-14, 4.56042e-14, 4.563583e-14, 4.561633e-14, 
    4.552156e-14, 4.550604e-14, 4.543884e-14, 4.542026e-14, 4.536904e-14, 
    4.532659e-14, 4.536536e-14, 4.540605e-14, 4.552161e-14, 4.56256e-14, 
    4.573892e-14, 4.576664e-14, 4.589875e-14, 4.579116e-14, 4.596859e-14, 
    4.581767e-14, 4.607883e-14, 4.560929e-14, 4.581332e-14, 4.54435e-14, 
    4.548341e-14, 4.55555e-14, 4.57208e-14, 4.563163e-14, 4.573593e-14, 
    4.550543e-14, 4.538559e-14, 4.535462e-14, 4.529672e-14, 4.535594e-14, 
    4.535113e-14, 4.540777e-14, 4.538958e-14, 4.552545e-14, 4.545249e-14, 
    4.565962e-14, 4.573512e-14, 4.59481e-14, 4.607843e-14, 4.621101e-14, 
    4.626946e-14, 4.628725e-14, 4.629468e-14 ;

 POT_F_DENIT =
  1.021875e-12, 1.024719e-12, 1.024165e-12, 1.026459e-12, 1.025186e-12, 
    1.026687e-12, 1.022448e-12, 1.024829e-12, 1.023308e-12, 1.022126e-12, 
    1.030908e-12, 1.026558e-12, 1.035418e-12, 1.032645e-12, 1.039603e-12, 
    1.034986e-12, 1.040533e-12, 1.039467e-12, 1.042669e-12, 1.041751e-12, 
    1.045846e-12, 1.04309e-12, 1.047964e-12, 1.045186e-12, 1.045621e-12, 
    1.042997e-12, 1.027436e-12, 1.03037e-12, 1.027261e-12, 1.027679e-12, 
    1.027491e-12, 1.02521e-12, 1.024062e-12, 1.021652e-12, 1.022088e-12, 
    1.023857e-12, 1.027864e-12, 1.026502e-12, 1.029929e-12, 1.029851e-12, 
    1.033664e-12, 1.031945e-12, 1.038351e-12, 1.03653e-12, 1.041788e-12, 
    1.040466e-12, 1.041726e-12, 1.041342e-12, 1.041729e-12, 1.03979e-12, 
    1.04062e-12, 1.038913e-12, 1.032273e-12, 1.034228e-12, 1.028394e-12, 
    1.024885e-12, 1.022551e-12, 1.020895e-12, 1.021128e-12, 1.021575e-12, 
    1.023867e-12, 1.02602e-12, 1.027661e-12, 1.028758e-12, 1.029839e-12, 
    1.033115e-12, 1.034844e-12, 1.038719e-12, 1.038018e-12, 1.039203e-12, 
    1.040334e-12, 1.042232e-12, 1.041919e-12, 1.042755e-12, 1.039168e-12, 
    1.041552e-12, 1.037615e-12, 1.038692e-12, 1.030142e-12, 1.026872e-12, 
    1.025485e-12, 1.024267e-12, 1.021308e-12, 1.023351e-12, 1.022545e-12, 
    1.024459e-12, 1.025676e-12, 1.025073e-12, 1.028787e-12, 1.027343e-12, 
    1.034946e-12, 1.031672e-12, 1.040202e-12, 1.038161e-12, 1.04069e-12, 
    1.039399e-12, 1.04161e-12, 1.039619e-12, 1.043065e-12, 1.043816e-12, 
    1.043302e-12, 1.045271e-12, 1.039506e-12, 1.041721e-12, 1.02506e-12, 
    1.025158e-12, 1.025615e-12, 1.023604e-12, 1.023481e-12, 1.021637e-12, 
    1.023276e-12, 1.023975e-12, 1.025745e-12, 1.026793e-12, 1.027788e-12, 
    1.029978e-12, 1.032423e-12, 1.03584e-12, 1.038293e-12, 1.039936e-12, 
    1.038927e-12, 1.039817e-12, 1.038822e-12, 1.038354e-12, 1.043534e-12, 
    1.040626e-12, 1.044987e-12, 1.044745e-12, 1.042771e-12, 1.044771e-12, 
    1.025226e-12, 1.02466e-12, 1.022699e-12, 1.024233e-12, 1.021435e-12, 
    1.023001e-12, 1.023901e-12, 1.027373e-12, 1.028134e-12, 1.028842e-12, 
    1.030238e-12, 1.032029e-12, 1.035172e-12, 1.037904e-12, 1.040397e-12, 
    1.040213e-12, 1.040278e-12, 1.040834e-12, 1.039454e-12, 1.04106e-12, 
    1.041329e-12, 1.040624e-12, 1.044712e-12, 1.043544e-12, 1.044738e-12, 
    1.043977e-12, 1.024843e-12, 1.025793e-12, 1.025279e-12, 1.026245e-12, 
    1.025564e-12, 1.028589e-12, 1.029496e-12, 1.033736e-12, 1.031994e-12, 
    1.034764e-12, 1.032274e-12, 1.032716e-12, 1.034855e-12, 1.032407e-12, 
    1.037753e-12, 1.03413e-12, 1.040855e-12, 1.037241e-12, 1.041081e-12, 
    1.040382e-12, 1.041536e-12, 1.042571e-12, 1.043871e-12, 1.046271e-12, 
    1.045714e-12, 1.04772e-12, 1.027209e-12, 1.028442e-12, 1.028332e-12, 
    1.029621e-12, 1.030574e-12, 1.03264e-12, 1.035953e-12, 1.034706e-12, 
    1.036992e-12, 1.037452e-12, 1.033976e-12, 1.03611e-12, 1.029261e-12, 
    1.030368e-12, 1.029708e-12, 1.027299e-12, 1.03499e-12, 1.031044e-12, 
    1.038327e-12, 1.03619e-12, 1.042422e-12, 1.039324e-12, 1.045408e-12, 
    1.048009e-12, 1.050452e-12, 1.05331e-12, 1.029113e-12, 1.028275e-12, 
    1.029773e-12, 1.031848e-12, 1.03377e-12, 1.036327e-12, 1.036587e-12, 
    1.037065e-12, 1.038304e-12, 1.039347e-12, 1.037216e-12, 1.039607e-12, 
    1.030626e-12, 1.035332e-12, 1.027952e-12, 1.030176e-12, 1.031719e-12, 
    1.031041e-12, 1.034557e-12, 1.035385e-12, 1.038752e-12, 1.037011e-12, 
    1.047367e-12, 1.042787e-12, 1.055482e-12, 1.051937e-12, 1.027982e-12, 
    1.029108e-12, 1.033029e-12, 1.031163e-12, 1.036495e-12, 1.037808e-12, 
    1.038873e-12, 1.040237e-12, 1.040382e-12, 1.04119e-12, 1.039865e-12, 
    1.041137e-12, 1.036327e-12, 1.038476e-12, 1.032574e-12, 1.034011e-12, 
    1.033349e-12, 1.032623e-12, 1.03486e-12, 1.037244e-12, 1.037293e-12, 
    1.038057e-12, 1.040213e-12, 1.036507e-12, 1.047958e-12, 1.04089e-12, 
    1.030336e-12, 1.032507e-12, 1.032815e-12, 1.031974e-12, 1.037675e-12, 
    1.03561e-12, 1.04117e-12, 1.039667e-12, 1.042128e-12, 1.040905e-12, 
    1.040724e-12, 1.039152e-12, 1.038173e-12, 1.035701e-12, 1.033687e-12, 
    1.03209e-12, 1.03246e-12, 1.034214e-12, 1.037388e-12, 1.04039e-12, 
    1.039732e-12, 1.041934e-12, 1.036098e-12, 1.038547e-12, 1.0376e-12, 
    1.040065e-12, 1.034671e-12, 1.039278e-12, 1.033493e-12, 1.034e-12, 
    1.035567e-12, 1.038721e-12, 1.039416e-12, 1.040161e-12, 1.0397e-12, 
    1.037473e-12, 1.037106e-12, 1.035525e-12, 1.035089e-12, 1.033885e-12, 
    1.032887e-12, 1.033798e-12, 1.034754e-12, 1.037469e-12, 1.039915e-12, 
    1.04258e-12, 1.043231e-12, 1.046347e-12, 1.043812e-12, 1.047995e-12, 
    1.04444e-12, 1.05059e-12, 1.039541e-12, 1.044344e-12, 1.035638e-12, 
    1.036575e-12, 1.038273e-12, 1.042161e-12, 1.04006e-12, 1.042516e-12, 
    1.037091e-12, 1.034276e-12, 1.033546e-12, 1.032186e-12, 1.033576e-12, 
    1.033463e-12, 1.034792e-12, 1.034364e-12, 1.037557e-12, 1.035842e-12, 
    1.040713e-12, 1.04249e-12, 1.047505e-12, 1.050577e-12, 1.053701e-12, 
    1.05508e-12, 1.055499e-12, 1.055674e-12 ;

 POT_F_NIT =
  4.01379e-11, 4.04843e-11, 4.041683e-11, 4.069712e-11, 4.05415e-11, 
    4.072521e-11, 4.020798e-11, 4.049806e-11, 4.031275e-11, 4.016898e-11, 
    4.124388e-11, 4.070961e-11, 4.180262e-11, 4.145908e-11, 4.232481e-11, 
    4.174906e-11, 4.244139e-11, 4.230813e-11, 4.270985e-11, 4.259455e-11, 
    4.311054e-11, 4.27631e-11, 4.337926e-11, 4.302742e-11, 4.308236e-11, 
    4.275164e-11, 4.081686e-11, 4.11772e-11, 4.079555e-11, 4.084683e-11, 
    4.082381e-11, 4.05447e-11, 4.040443e-11, 4.011144e-11, 4.016454e-11, 
    4.037977e-11, 4.086986e-11, 4.070314e-11, 4.112395e-11, 4.111443e-11, 
    4.158549e-11, 4.137275e-11, 4.216865e-11, 4.194164e-11, 4.259935e-11, 
    4.243344e-11, 4.259155e-11, 4.254357e-11, 4.259216e-11, 4.234898e-11, 
    4.245307e-11, 4.223941e-11, 4.141261e-11, 4.165474e-11, 4.093471e-11, 
    4.050488e-11, 4.022066e-11, 4.001962e-11, 4.0048e-11, 4.010215e-11, 
    4.038102e-11, 4.064411e-11, 4.084521e-11, 4.098e-11, 4.111304e-11, 
    4.151715e-11, 4.173184e-11, 4.221463e-11, 4.212728e-11, 4.22753e-11, 
    4.241695e-11, 4.265533e-11, 4.261604e-11, 4.272124e-11, 4.227136e-11, 
    4.257008e-11, 4.207753e-11, 4.221195e-11, 4.114933e-11, 4.07481e-11, 
    4.05782e-11, 4.042976e-11, 4.006983e-11, 4.031821e-11, 4.02202e-11, 
    4.045355e-11, 4.06022e-11, 4.052864e-11, 4.098369e-11, 4.080646e-11, 
    4.174457e-11, 4.133914e-11, 4.240042e-11, 4.214519e-11, 4.24617e-11, 
    4.230004e-11, 4.257723e-11, 4.232771e-11, 4.276041e-11, 4.285494e-11, 
    4.279032e-11, 4.303877e-11, 4.231387e-11, 4.259151e-11, 4.05266e-11, 
    4.05386e-11, 4.059448e-11, 4.03491e-11, 4.033411e-11, 4.010996e-11, 
    4.030937e-11, 4.039444e-11, 4.061081e-11, 4.073908e-11, 4.08612e-11, 
    4.113038e-11, 4.143208e-11, 4.185587e-11, 4.21617e-11, 4.236735e-11, 
    4.224118e-11, 4.235256e-11, 4.222805e-11, 4.216976e-11, 4.28195e-11, 
    4.245403e-11, 4.300298e-11, 4.297251e-11, 4.272371e-11, 4.297593e-11, 
    4.054701e-11, 4.047801e-11, 4.023897e-11, 4.042598e-11, 4.008558e-11, 
    4.027594e-11, 4.038559e-11, 4.081016e-11, 4.090374e-11, 4.099062e-11, 
    4.116248e-11, 4.138359e-11, 4.177297e-11, 4.211327e-11, 4.242518e-11, 
    4.240228e-11, 4.241034e-11, 4.248016e-11, 4.23073e-11, 4.250857e-11, 
    4.25424e-11, 4.245397e-11, 4.296841e-11, 4.282111e-11, 4.297184e-11, 
    4.287589e-11, 4.050043e-11, 4.061657e-11, 4.055378e-11, 4.067188e-11, 
    4.058865e-11, 4.095938e-11, 4.107087e-11, 4.159462e-11, 4.137924e-11, 
    4.172227e-11, 4.141401e-11, 4.146854e-11, 4.173349e-11, 4.143062e-11, 
    4.209447e-11, 4.164381e-11, 4.248287e-11, 4.203071e-11, 4.251128e-11, 
    4.242379e-11, 4.256868e-11, 4.269867e-11, 4.286247e-11, 4.31656e-11, 
    4.309529e-11, 4.334942e-11, 4.079003e-11, 4.094126e-11, 4.092793e-11, 
    4.108647e-11, 4.120394e-11, 4.145912e-11, 4.18701e-11, 4.171529e-11, 
    4.199969e-11, 4.205691e-11, 4.162491e-11, 4.188988e-11, 4.10426e-11, 
    4.117888e-11, 4.10977e-11, 4.080189e-11, 4.175092e-11, 4.126246e-11, 
    4.216672e-11, 4.190038e-11, 4.268011e-11, 4.229141e-11, 4.305662e-11, 
    4.338594e-11, 4.369702e-11, 4.406205e-11, 4.102392e-11, 4.092101e-11, 
    4.110534e-11, 4.13611e-11, 4.159911e-11, 4.191665e-11, 4.19492e-11, 
    4.200885e-11, 4.216355e-11, 4.229386e-11, 4.202771e-11, 4.232655e-11, 
    4.121053e-11, 4.179345e-11, 4.088209e-11, 4.115544e-11, 4.134594e-11, 
    4.126231e-11, 4.169757e-11, 4.180049e-11, 4.222012e-11, 4.200292e-11, 
    4.330453e-11, 4.272613e-11, 4.434102e-11, 4.388661e-11, 4.088508e-11, 
    4.102354e-11, 4.150734e-11, 4.127678e-11, 4.193788e-11, 4.210144e-11, 
    4.223463e-11, 4.240524e-11, 4.242366e-11, 4.252493e-11, 4.235904e-11, 
    4.251836e-11, 4.191728e-11, 4.218534e-11, 4.145184e-11, 4.162975e-11, 
    4.154785e-11, 4.14581e-11, 4.173538e-11, 4.203185e-11, 4.203818e-11, 
    4.213347e-11, 4.240265e-11, 4.194049e-11, 4.337948e-11, 4.248784e-11, 
    4.11748e-11, 4.144271e-11, 4.148103e-11, 4.137709e-11, 4.208502e-11, 
    4.182779e-11, 4.252246e-11, 4.233413e-11, 4.264292e-11, 4.248933e-11, 
    4.246675e-11, 4.226995e-11, 4.214766e-11, 4.183954e-11, 4.158968e-11, 
    4.139211e-11, 4.1438e-11, 4.165518e-11, 4.205001e-11, 4.242529e-11, 
    4.234293e-11, 4.261936e-11, 4.188967e-11, 4.219486e-11, 4.207676e-11, 
    4.238502e-11, 4.171117e-11, 4.228475e-11, 4.156521e-11, 4.162803e-11, 
    4.182268e-11, 4.221566e-11, 4.230284e-11, 4.239606e-11, 4.233851e-11, 
    4.206008e-11, 4.201455e-11, 4.181792e-11, 4.176371e-11, 4.161431e-11, 
    4.149082e-11, 4.160363e-11, 4.172227e-11, 4.206016e-11, 4.236586e-11, 
    4.270047e-11, 4.278256e-11, 4.317565e-11, 4.285552e-11, 4.338446e-11, 
    4.293457e-11, 4.371487e-11, 4.231808e-11, 4.292144e-11, 4.183155e-11, 
    4.194826e-11, 4.21598e-11, 4.264705e-11, 4.238362e-11, 4.269177e-11, 
    4.201276e-11, 4.16627e-11, 4.157235e-11, 4.14041e-11, 4.15762e-11, 
    4.156218e-11, 4.172718e-11, 4.167412e-11, 4.207139e-11, 4.185775e-11, 
    4.246613e-11, 4.268928e-11, 4.332271e-11, 4.371341e-11, 4.411298e-11, 
    4.428997e-11, 4.434392e-11, 4.436648e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001208392, 0.00120832, 0.001208334, 0.001208277, 0.001208308, 
    0.001208271, 0.001208376, 0.001208318, 0.001208355, 0.001208384, 
    0.001208168, 0.001208274, 0.001208053, 0.001208121, 0.001207947, 
    0.001208064, 0.001207923, 0.001207949, 0.001207868, 0.001207891, 
    0.001207791, 0.001207858, 0.001207737, 0.001207806, 0.001207796, 
    0.00120786, 0.001208251, 0.001208182, 0.001208256, 0.001208246, 
    0.00120825, 0.001208308, 0.001208337, 0.001208396, 0.001208385, 
    0.001208342, 0.001208241, 0.001208275, 0.001208188, 0.00120819, 
    0.001208096, 0.001208138, 0.001207977, 0.001208023, 0.00120789, 
    0.001207924, 0.001207892, 0.001207901, 0.001207892, 0.001207941, 
    0.00120792, 0.001207962, 0.001208131, 0.001208082, 0.001208228, 
    0.001208318, 0.001208374, 0.001208415, 0.001208409, 0.001208398, 
    0.001208341, 0.001208287, 0.001208245, 0.001208218, 0.001208191, 
    0.001208112, 0.001208067, 0.001207968, 0.001207985, 0.001207956, 
    0.001207927, 0.00120788, 0.001207887, 0.001207867, 0.001207956, 
    0.001207897, 0.001207996, 0.001207968, 0.001208188, 0.001208265, 
    0.001208302, 0.001208331, 0.001208405, 0.001208354, 0.001208374, 
    0.001208325, 0.001208295, 0.00120831, 0.001208217, 0.001208253, 
    0.001208065, 0.001208146, 0.00120793, 0.001207981, 0.001207918, 
    0.00120795, 0.001207895, 0.001207944, 0.001207859, 0.00120784, 
    0.001207853, 0.001207803, 0.001207947, 0.001207892, 0.001208311, 
    0.001208308, 0.001208297, 0.001208348, 0.001208351, 0.001208397, 
    0.001208355, 0.001208338, 0.001208293, 0.001208267, 0.001208242, 
    0.001208188, 0.001208127, 0.001208042, 0.001207978, 0.001207936, 
    0.001207961, 0.001207939, 0.001207964, 0.001207976, 0.001207847, 
    0.00120792, 0.00120781, 0.001207816, 0.001207866, 0.001207816, 
    0.001208307, 0.00120832, 0.00120837, 0.001208331, 0.001208401, 
    0.001208363, 0.001208341, 0.001208254, 0.001208233, 0.001208216, 
    0.001208181, 0.001208136, 0.001208058, 0.001207988, 0.001207925, 
    0.001207929, 0.001207928, 0.001207914, 0.001207949, 0.001207908, 
    0.001207902, 0.001207919, 0.001207817, 0.001207846, 0.001207817, 
    0.001207835, 0.001208316, 0.001208292, 0.001208305, 0.001208281, 
    0.001208298, 0.001208223, 0.001208201, 0.001208095, 0.001208137, 
    0.001208069, 0.00120813, 0.001208119, 0.001208068, 0.001208126, 
    0.001207994, 0.001208085, 0.001207914, 0.001208008, 0.001207908, 
    0.001207925, 0.001207896, 0.001207871, 0.001207838, 0.001207779, 
    0.001207793, 0.001207743, 0.001208257, 0.001208227, 0.001208228, 
    0.001208196, 0.001208173, 0.001208121, 0.001208038, 0.001208069, 
    0.001208012, 0.001208, 0.001208087, 0.001208035, 0.001208206, 
    0.001208179, 0.001208194, 0.001208255, 0.001208063, 0.001208162, 
    0.001207977, 0.001208032, 0.001207875, 0.001207953, 0.0012078, 
    0.001207737, 0.001207674, 0.001207605, 0.001208209, 0.00120823, 
    0.001208192, 0.001208142, 0.001208093, 0.001208029, 0.001208022, 
    0.00120801, 0.001207977, 0.001207951, 0.001208007, 0.001207945, 
    0.001208175, 0.001208054, 0.001208238, 0.001208184, 0.001208144, 
    0.001208161, 0.001208072, 0.001208052, 0.001207967, 0.001208011, 
    0.001207754, 0.001207867, 0.00120755, 0.001207639, 0.001208237, 
    0.001208209, 0.001208112, 0.001208158, 0.001208024, 0.001207992, 
    0.001207963, 0.00120793, 0.001207925, 0.001207905, 0.001207938, 
    0.001207906, 0.001208029, 0.001207973, 0.001208122, 0.001208086, 
    0.001208102, 0.001208121, 0.001208065, 0.001208007, 0.001208004, 
    0.001207984, 0.001207935, 0.001208024, 0.001207742, 0.001207917, 
    0.001208178, 0.001208126, 0.001208116, 0.001208137, 0.001207995, 
    0.001208047, 0.001207906, 0.001207943, 0.001207882, 0.001207912, 
    0.001207917, 0.001207956, 0.001207981, 0.001208044, 0.001208095, 
    0.001208134, 0.001208125, 0.001208082, 0.001208003, 0.001207926, 
    0.001207942, 0.001207886, 0.001208034, 0.001207972, 0.001207997, 
    0.001207933, 0.00120807, 0.001207957, 0.001208099, 0.001208086, 
    0.001208048, 0.001207969, 0.001207949, 0.001207931, 0.001207942, 
    0.001208, 0.001208009, 0.001208048, 0.00120806, 0.001208089, 0.001208114, 
    0.001208092, 0.001208068, 0.001208, 0.001207937, 0.001207871, 
    0.001207854, 0.00120778, 0.001207842, 0.001207741, 0.00120783, 
    0.001207675, 0.001207949, 0.00120783, 0.001208045, 0.001208022, 
    0.001207979, 0.001207883, 0.001207933, 0.001207873, 0.001208009, 
    0.001208081, 0.001208098, 0.001208132, 0.001208097, 0.0012081, 
    0.001208066, 0.001208077, 0.001207998, 0.00120804, 0.001207917, 
    0.001207874, 0.001207748, 0.001207673, 0.001207593, 0.001207559, 
    0.001207548, 0.001207544 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  -1.287405e-07, -1.290487e-07, -1.289887e-07, -1.292371e-07, -1.290991e-07, 
    -1.292618e-07, -1.288028e-07, -1.290611e-07, -1.288961e-07, 
    -1.287679e-07, -1.297172e-07, -1.292481e-07, -1.302e-07, -1.299027e-07, 
    -1.306518e-07, -1.301541e-07, -1.307511e-07, -1.306369e-07, 
    -1.309787e-07, -1.308809e-07, -1.313181e-07, -1.310238e-07, 
    -1.315432e-07, -1.312476e-07, -1.312941e-07, -1.310142e-07, 
    -1.293421e-07, -1.296591e-07, -1.293234e-07, -1.293686e-07, 
    -1.293482e-07, -1.291022e-07, -1.289782e-07, -1.287165e-07, -1.28764e-07, 
    -1.28956e-07, -1.293889e-07, -1.29242e-07, -1.296108e-07, -1.296025e-07, 
    -1.300121e-07, -1.298276e-07, -1.305176e-07, -1.303189e-07, 
    -1.308849e-07, -1.307438e-07, -1.308784e-07, -1.308375e-07, 
    -1.308789e-07, -1.306719e-07, -1.307607e-07, -1.305782e-07, 
    -1.298623e-07, -1.300721e-07, -1.294456e-07, -1.290677e-07, 
    -1.288142e-07, -1.286345e-07, -1.286599e-07, -1.287085e-07, 
    -1.289571e-07, -1.291899e-07, -1.293668e-07, -1.29485e-07, -1.296013e-07, 
    -1.29954e-07, -1.30139e-07, -1.305573e-07, -1.30482e-07, -1.306092e-07, 
    -1.307298e-07, -1.309327e-07, -1.308992e-07, -1.309886e-07, 
    -1.306054e-07, -1.308604e-07, -1.304356e-07, -1.305547e-07, 
    -1.296349e-07, -1.292816e-07, -1.291325e-07, -1.290003e-07, 
    -1.286795e-07, -1.289012e-07, -1.288139e-07, -1.290211e-07, 
    -1.291529e-07, -1.290876e-07, -1.294883e-07, -1.293329e-07, -1.3015e-07, 
    -1.297987e-07, -1.307157e-07, -1.304975e-07, -1.307679e-07, 
    -1.306299e-07, -1.308664e-07, -1.306535e-07, -1.310217e-07, -1.31102e-07, 
    -1.310472e-07, -1.312568e-07, -1.306418e-07, -1.308786e-07, 
    -1.290859e-07, -1.290965e-07, -1.291459e-07, -1.289287e-07, 
    -1.289153e-07, -1.287153e-07, -1.288931e-07, -1.289689e-07, 
    -1.291603e-07, -1.292737e-07, -1.29381e-07, -1.296167e-07, -1.298795e-07, 
    -1.302456e-07, -1.305116e-07, -1.306874e-07, -1.305795e-07, 
    -1.306748e-07, -1.305684e-07, -1.305184e-07, -1.31072e-07, -1.307616e-07, 
    -1.312267e-07, -1.312009e-07, -1.309908e-07, -1.312038e-07, -1.29104e-07, 
    -1.290428e-07, -1.288305e-07, -1.289966e-07, -1.286935e-07, 
    -1.288635e-07, -1.289613e-07, -1.293366e-07, -1.294182e-07, 
    -1.294945e-07, -1.296446e-07, -1.298371e-07, -1.301741e-07, 
    -1.304703e-07, -1.307367e-07, -1.307172e-07, -1.307241e-07, 
    -1.307837e-07, -1.306362e-07, -1.308079e-07, -1.308369e-07, 
    -1.307614e-07, -1.311975e-07, -1.310731e-07, -1.312004e-07, 
    -1.311193e-07, -1.290626e-07, -1.291655e-07, -1.2911e-07, -1.292146e-07, 
    -1.29141e-07, -1.294676e-07, -1.295652e-07, -1.300205e-07, -1.298334e-07, 
    -1.301305e-07, -1.298635e-07, -1.299109e-07, -1.30141e-07, -1.298778e-07, 
    -1.304509e-07, -1.300633e-07, -1.30786e-07, -1.303966e-07, -1.308102e-07, 
    -1.307356e-07, -1.308589e-07, -1.309695e-07, -1.311081e-07, 
    -1.313639e-07, -1.313046e-07, -1.31518e-07, -1.293184e-07, -1.294515e-07, 
    -1.294394e-07, -1.295782e-07, -1.296809e-07, -1.299025e-07, 
    -1.302576e-07, -1.301241e-07, -1.303688e-07, -1.304181e-07, -1.30046e-07, 
    -1.302748e-07, -1.295401e-07, -1.296596e-07, -1.295882e-07, 
    -1.293291e-07, -1.301554e-07, -1.297323e-07, -1.30516e-07, -1.302836e-07, 
    -1.309538e-07, -1.306231e-07, -1.312721e-07, -1.315494e-07, -1.31808e-07, 
    -1.321114e-07, -1.295236e-07, -1.294333e-07, -1.295946e-07, -1.29818e-07, 
    -1.300239e-07, -1.302976e-07, -1.303254e-07, -1.303768e-07, 
    -1.305131e-07, -1.306246e-07, -1.303934e-07, -1.306526e-07, 
    -1.296879e-07, -1.301919e-07, -1.293995e-07, -1.296392e-07, 
    -1.298047e-07, -1.297318e-07, -1.301087e-07, -1.301975e-07, -1.30562e-07, 
    -1.303716e-07, -1.314813e-07, -1.309933e-07, -1.323407e-07, 
    -1.319661e-07, -1.294019e-07, -1.295231e-07, -1.299447e-07, 
    -1.297443e-07, -1.303157e-07, -1.304563e-07, -1.305739e-07, -1.3072e-07, 
    -1.307355e-07, -1.308219e-07, -1.306803e-07, -1.308162e-07, 
    -1.302982e-07, -1.305319e-07, -1.298961e-07, -1.300504e-07, 
    -1.299793e-07, -1.299016e-07, -1.301414e-07, -1.303971e-07, -1.30402e-07, 
    -1.304877e-07, -1.307198e-07, -1.303179e-07, -1.315453e-07, 
    -1.307921e-07, -1.296553e-07, -1.29889e-07, -1.299216e-07, -1.298313e-07, 
    -1.304423e-07, -1.302212e-07, -1.308197e-07, -1.30659e-07, -1.30922e-07, 
    -1.307915e-07, -1.307723e-07, -1.306042e-07, -1.304996e-07, 
    -1.302314e-07, -1.300158e-07, -1.298443e-07, -1.298842e-07, 
    -1.300725e-07, -1.304126e-07, -1.307372e-07, -1.30667e-07, -1.309021e-07, 
    -1.302743e-07, -1.305403e-07, -1.304355e-07, -1.307027e-07, 
    -1.301206e-07, -1.306187e-07, -1.299943e-07, -1.300487e-07, 
    -1.302167e-07, -1.305585e-07, -1.306323e-07, -1.307122e-07, 
    -1.306628e-07, -1.304211e-07, -1.303818e-07, -1.302125e-07, 
    -1.301661e-07, -1.300368e-07, -1.2993e-07, -1.300277e-07, -1.301304e-07, 
    -1.30421e-07, -1.306865e-07, -1.309711e-07, -1.310405e-07, -1.313734e-07, 
    -1.311033e-07, -1.315496e-07, -1.311715e-07, -1.318245e-07, 
    -1.306465e-07, -1.311592e-07, -1.302242e-07, -1.303246e-07, 
    -1.305105e-07, -1.309263e-07, -1.307014e-07, -1.309641e-07, 
    -1.303802e-07, -1.300793e-07, -1.300006e-07, -1.298549e-07, 
    -1.300039e-07, -1.299918e-07, -1.301343e-07, -1.300885e-07, 
    -1.304306e-07, -1.302468e-07, -1.30772e-07, -1.309619e-07, -1.314958e-07, 
    -1.318223e-07, -1.321527e-07, -1.322985e-07, -1.323428e-07, -1.323614e-07 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.022795e-06, 3.029914e-06, 3.028535e-06, 3.034268e-06, 3.031096e-06, 
    3.034841e-06, 3.024248e-06, 3.030189e-06, 3.026402e-06, 3.023449e-06, 
    3.045301e-06, 3.034525e-06, 3.056584e-06, 3.049695e-06, 3.067742e-06, 
    3.055499e-06, 3.070077e-06, 3.067429e-06, 3.075451e-06, 3.073154e-06, 
    3.083377e-06, 3.076512e-06, 3.088716e-06, 3.081749e-06, 3.08283e-06, 
    3.076282e-06, 3.036713e-06, 3.043952e-06, 3.03628e-06, 3.037313e-06, 
    3.036854e-06, 3.031153e-06, 3.028259e-06, 3.022266e-06, 3.023358e-06, 
    3.027768e-06, 3.037778e-06, 3.034408e-06, 3.042944e-06, 3.042752e-06, 
    3.052241e-06, 3.047963e-06, 3.064639e-06, 3.059399e-06, 3.07325e-06, 
    3.069937e-06, 3.073091e-06, 3.072137e-06, 3.073103e-06, 3.068245e-06, 
    3.070325e-06, 3.066059e-06, 3.04876e-06, 3.053628e-06, 3.039099e-06, 
    3.030307e-06, 3.024505e-06, 3.020373e-06, 3.020956e-06, 3.022065e-06, 
    3.027793e-06, 3.033201e-06, 3.037296e-06, 3.040028e-06, 3.042724e-06, 
    3.050827e-06, 3.055163e-06, 3.065548e-06, 3.063816e-06, 3.066764e-06, 
    3.069608e-06, 3.07436e-06, 3.07358e-06, 3.07567e-06, 3.066699e-06, 
    3.072654e-06, 3.062126e-06, 3.06551e-06, 3.043385e-06, 3.03532e-06, 
    3.031815e-06, 3.028797e-06, 3.021404e-06, 3.026505e-06, 3.024492e-06, 
    3.029298e-06, 3.032342e-06, 3.030839e-06, 3.040103e-06, 3.036507e-06, 
    3.05542e-06, 3.047274e-06, 3.069276e-06, 3.064173e-06, 3.070503e-06, 
    3.067275e-06, 3.0728e-06, 3.067828e-06, 3.076454e-06, 3.078325e-06, 
    3.077045e-06, 3.081988e-06, 3.06755e-06, 3.073084e-06, 3.030793e-06, 
    3.031038e-06, 3.032186e-06, 3.027138e-06, 3.026834e-06, 3.022232e-06, 
    3.026334e-06, 3.028074e-06, 3.032524e-06, 3.035137e-06, 3.037615e-06, 
    3.043067e-06, 3.049144e-06, 3.057664e-06, 3.064503e-06, 3.068621e-06, 
    3.0661e-06, 3.068325e-06, 3.065835e-06, 3.064672e-06, 3.077619e-06, 
    3.07034e-06, 3.081277e-06, 3.080674e-06, 3.075717e-06, 3.080742e-06, 
    3.031211e-06, 3.029801e-06, 3.024884e-06, 3.028732e-06, 3.021733e-06, 
    3.025641e-06, 3.027883e-06, 3.036566e-06, 3.038482e-06, 3.040237e-06, 
    3.043721e-06, 3.048181e-06, 3.056003e-06, 3.063526e-06, 3.069777e-06, 
    3.06932e-06, 3.06948e-06, 3.070869e-06, 3.067418e-06, 3.071437e-06, 
    3.072105e-06, 3.070348e-06, 3.080593e-06, 3.077666e-06, 3.080661e-06, 
    3.078757e-06, 3.030261e-06, 3.032637e-06, 3.031352e-06, 3.033765e-06, 
    3.032059e-06, 3.039588e-06, 3.041842e-06, 3.052407e-06, 3.04809e-06, 
    3.054982e-06, 3.048795e-06, 3.049887e-06, 3.055177e-06, 3.049134e-06, 
    3.062436e-06, 3.053388e-06, 3.070924e-06, 3.061143e-06, 3.071491e-06, 
    3.069749e-06, 3.072641e-06, 3.075224e-06, 3.078487e-06, 3.084491e-06, 
    3.083103e-06, 3.088139e-06, 3.036174e-06, 3.03923e-06, 3.038974e-06, 
    3.042183e-06, 3.044554e-06, 3.049706e-06, 3.057958e-06, 3.054858e-06, 
    3.060564e-06, 3.061706e-06, 3.053045e-06, 3.058349e-06, 3.041286e-06, 
    3.044029e-06, 3.042406e-06, 3.036407e-06, 3.055554e-06, 3.04572e-06, 
    3.064602e-06, 3.05857e-06, 3.074854e-06, 3.067083e-06, 3.082336e-06, 
    3.08883e-06, 3.095009e-06, 3.102163e-06, 3.040913e-06, 3.038834e-06, 
    3.042569e-06, 3.04771e-06, 3.052518e-06, 3.058892e-06, 3.059552e-06, 
    3.060743e-06, 3.064546e-06, 3.067151e-06, 3.061106e-06, 3.067806e-06, 
    3.044638e-06, 3.056414e-06, 3.038036e-06, 3.043552e-06, 3.047413e-06, 
    3.045734e-06, 3.054507e-06, 3.056572e-06, 3.065663e-06, 3.060631e-06, 
    3.087215e-06, 3.07575e-06, 3.10766e-06, 3.098721e-06, 3.038105e-06, 
    3.040912e-06, 3.050662e-06, 3.046027e-06, 3.059325e-06, 3.062595e-06, 
    3.06597e-06, 3.069367e-06, 3.069744e-06, 3.07176e-06, 3.068455e-06, 
    3.071635e-06, 3.058906e-06, 3.064979e-06, 3.049564e-06, 3.053135e-06, 
    3.051497e-06, 3.04969e-06, 3.055266e-06, 3.061187e-06, 3.061335e-06, 
    3.063932e-06, 3.069243e-06, 3.059379e-06, 3.088655e-06, 3.070955e-06, 
    3.043973e-06, 3.04935e-06, 3.050144e-06, 3.048057e-06, 3.062267e-06, 
    3.057113e-06, 3.071714e-06, 3.067957e-06, 3.074119e-06, 3.071055e-06, 
    3.070603e-06, 3.066674e-06, 3.064224e-06, 3.057345e-06, 3.052327e-06, 
    3.048362e-06, 3.049286e-06, 3.053643e-06, 3.061554e-06, 3.069769e-06, 
    3.068118e-06, 3.073651e-06, 3.058359e-06, 3.065161e-06, 3.062093e-06, 
    3.068972e-06, 3.054771e-06, 3.066899e-06, 3.051846e-06, 3.053107e-06, 
    3.05701e-06, 3.06556e-06, 3.067331e-06, 3.069184e-06, 3.068046e-06, 
    3.061759e-06, 3.060855e-06, 3.056921e-06, 3.055824e-06, 3.052834e-06, 
    3.05035e-06, 3.052614e-06, 3.054989e-06, 3.061771e-06, 3.068581e-06, 
    3.075257e-06, 3.0769e-06, 3.084654e-06, 3.078311e-06, 3.08875e-06, 
    3.079829e-06, 3.0953e-06, 3.067594e-06, 3.079611e-06, 3.057195e-06, 
    3.059535e-06, 3.064447e-06, 3.074171e-06, 3.068943e-06, 3.075068e-06, 
    3.060821e-06, 3.053782e-06, 3.051989e-06, 3.048599e-06, 3.052066e-06, 
    3.051785e-06, 3.055103e-06, 3.054038e-06, 3.061996e-06, 3.057721e-06, 
    3.070586e-06, 3.075025e-06, 3.087603e-06, 3.095309e-06, 3.103196e-06, 
    3.106669e-06, 3.107728e-06, 3.108169e-06 ;

 QVEGE =
  -6.482325e-07, -6.477935e-07, -6.478768e-07, -6.475265e-07, -6.477176e-07, 
    -6.474905e-07, -6.481396e-07, -6.477796e-07, -6.480072e-07, 
    -6.481876e-07, -6.468545e-07, -6.475098e-07, -6.461386e-07, -6.46561e-07, 
    -6.454867e-07, -6.462099e-07, -6.45338e-07, -6.454985e-07, -6.449918e-07, 
    -6.451367e-07, -6.445046e-07, -6.449247e-07, -6.441597e-07, 
    -6.446002e-07, -6.44535e-07, -6.4494e-07, -6.473695e-07, -6.469393e-07, 
    -6.47397e-07, -6.473354e-07, -6.473609e-07, -6.477168e-07, -6.479016e-07, 
    -6.482597e-07, -6.481932e-07, -6.479266e-07, -6.473073e-07, -6.47512e-07, 
    -6.469774e-07, -6.469893e-07, -6.464019e-07, -6.466663e-07, 
    -6.456734e-07, -6.45953e-07, -6.451305e-07, -6.453401e-07, -6.451419e-07, 
    -6.452009e-07, -6.451411e-07, -6.454478e-07, -6.453171e-07, 
    -6.455834e-07, -6.466184e-07, -6.463177e-07, -6.472226e-07, 
    -6.477799e-07, -6.481255e-07, -6.483768e-07, -6.483414e-07, 
    -6.482755e-07, -6.479253e-07, -6.475868e-07, -6.473308e-07, 
    -6.471606e-07, -6.469912e-07, -6.465045e-07, -6.462271e-07, 
    -6.456208e-07, -6.457232e-07, -6.455437e-07, -6.453605e-07, 
    -6.450628e-07, -6.451107e-07, -6.449811e-07, -6.455427e-07, 
    -6.451727e-07, -6.457811e-07, -6.456178e-07, -6.469763e-07, 
    -6.474554e-07, -6.476849e-07, -6.47862e-07, -6.483147e-07, -6.48004e-07, 
    -6.481274e-07, -6.478271e-07, -6.476403e-07, -6.477314e-07, 
    -6.471558e-07, -6.473812e-07, -6.462107e-07, -6.467133e-07, 
    -6.453818e-07, -6.457015e-07, -6.453039e-07, -6.455055e-07, 
    -6.451623e-07, -6.454712e-07, -6.449303e-07, -6.448157e-07, 
    -6.448947e-07, -6.445799e-07, -6.454891e-07, -6.45145e-07, -6.477354e-07, 
    -6.477208e-07, -6.476487e-07, -6.479655e-07, -6.479831e-07, 
    -6.482631e-07, -6.480112e-07, -6.479062e-07, -6.476269e-07, 
    -6.474671e-07, -6.473129e-07, -6.469724e-07, -6.465984e-07, 
    -6.460671e-07, -6.456812e-07, -6.454213e-07, -6.455787e-07, -6.4544e-07, 
    -6.455962e-07, -6.45668e-07, -6.448607e-07, -6.453178e-07, -6.446253e-07, 
    -6.446627e-07, -6.449793e-07, -6.446584e-07, -6.4771e-07, -6.477953e-07, 
    -6.481012e-07, -6.478618e-07, -6.482931e-07, -6.480559e-07, 
    -6.479215e-07, -6.473833e-07, -6.472572e-07, -6.471498e-07, -6.4693e-07, 
    -6.466529e-07, -6.461698e-07, -6.457449e-07, -6.453486e-07, -6.45377e-07, 
    -6.453673e-07, -6.452817e-07, -6.454978e-07, -6.452459e-07, 
    -6.452066e-07, -6.453141e-07, -6.446679e-07, -6.448527e-07, 
    -6.446635e-07, -6.447831e-07, -6.477668e-07, -6.476215e-07, 
    -6.477006e-07, -6.475536e-07, -6.476596e-07, -6.471963e-07, -6.47057e-07, 
    -6.463983e-07, -6.466601e-07, -6.462346e-07, -6.466144e-07, -6.46549e-07, 
    -6.462338e-07, -6.46592e-07, -6.457724e-07, -6.463405e-07, -6.452784e-07, 
    -6.458594e-07, -6.452424e-07, -6.453503e-07, -6.451684e-07, 
    -6.450086e-07, -6.448013e-07, -6.444264e-07, -6.445121e-07, 
    -6.441924e-07, -6.474017e-07, -6.472153e-07, -6.472259e-07, 
    -6.470263e-07, -6.468798e-07, -6.465569e-07, -6.460456e-07, 
    -6.462363e-07, -6.458797e-07, -6.4581e-07, -6.463483e-07, -6.460236e-07, 
    -6.470859e-07, -6.469195e-07, -6.470143e-07, -6.473904e-07, 
    -6.462005e-07, -6.468131e-07, -6.456759e-07, -6.460063e-07, 
    -6.450322e-07, -6.455254e-07, -6.445606e-07, -6.441599e-07, 
    -6.437531e-07, -6.433075e-07, -6.47107e-07, -6.472345e-07, -6.470009e-07, 
    -6.466889e-07, -6.463843e-07, -6.459871e-07, -6.459433e-07, 
    -6.458704e-07, -6.456762e-07, -6.455137e-07, -6.45853e-07, -6.454723e-07, 
    -6.468927e-07, -6.461444e-07, -6.472881e-07, -6.469506e-07, 
    -6.467046e-07, -6.468061e-07, -6.462566e-07, -6.461288e-07, 
    -6.456122e-07, -6.458753e-07, -6.442642e-07, -6.449831e-07, 
    -6.429465e-07, -6.43525e-07, -6.472805e-07, -6.471047e-07, -6.465028e-07, 
    -6.467872e-07, -6.459575e-07, -6.457549e-07, -6.455869e-07, 
    -6.453783e-07, -6.453515e-07, -6.452269e-07, -6.454317e-07, 
    -6.452327e-07, -6.459863e-07, -6.456507e-07, -6.465643e-07, 
    -6.463457e-07, -6.464443e-07, -6.465567e-07, -6.462101e-07, 
    -6.458492e-07, -6.45832e-07, -6.457196e-07, -6.454129e-07, -6.459539e-07, 
    -6.441885e-07, -6.453016e-07, -6.469132e-07, -6.465887e-07, 
    -6.465311e-07, -6.466584e-07, -6.457756e-07, -6.460974e-07, 
    -6.452286e-07, -6.45463e-07, -6.45076e-07, -6.452694e-07, -6.452983e-07, 
    -6.455435e-07, -6.456984e-07, -6.460845e-07, -6.463968e-07, 
    -6.466387e-07, -6.465818e-07, -6.463155e-07, -6.458249e-07, 
    -6.453533e-07, -6.454586e-07, -6.451053e-07, -6.460182e-07, -6.45643e-07, 
    -6.457901e-07, -6.454007e-07, -6.462435e-07, -6.455554e-07, 
    -6.464225e-07, -6.463446e-07, -6.461037e-07, -6.456236e-07, 
    -6.455024e-07, -6.453898e-07, -6.454573e-07, -6.458106e-07, 
    -6.458645e-07, -6.461073e-07, -6.46179e-07, -6.463609e-07, -6.465156e-07, 
    -6.463766e-07, -6.462324e-07, -6.458066e-07, -6.454282e-07, 
    -6.450078e-07, -6.449009e-07, -6.444299e-07, -6.448266e-07, 
    -6.441842e-07, -6.447505e-07, -6.437576e-07, -6.455012e-07, 
    -6.447478e-07, -6.460896e-07, -6.459438e-07, -6.456914e-07, 
    -6.450838e-07, -6.454025e-07, -6.450251e-07, -6.458658e-07, -6.46311e-07, 
    -6.464143e-07, -6.466258e-07, -6.464094e-07, -6.464267e-07, 
    -6.462197e-07, -6.462857e-07, -6.457922e-07, -6.460571e-07, 
    -6.453015e-07, -6.450257e-07, -6.442294e-07, -6.437432e-07, 
    -6.432296e-07, -6.43007e-07, -6.429382e-07, -6.4291e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.7115, 84.71105, 84.71114, 84.71078, 84.71098, 84.71075, 84.71141, 
    84.71104, 84.71127, 84.71146, 84.71015, 84.71077, 84.70958, 84.70992, 
    84.70865, 84.70963, 84.70854, 84.70866, 84.7083, 84.7084, 84.70796, 
    84.70825, 84.70773, 84.70803, 84.70798, 84.70827, 84.71064, 84.71023, 
    84.71066, 84.7106, 84.71063, 84.71098, 84.71116, 84.71153, 84.71146, 
    84.71119, 84.71058, 84.71078, 84.71027, 84.71029, 84.70979, 84.71001, 
    84.70879, 84.70944, 84.7084, 84.70855, 84.7084, 84.70845, 84.7084, 
    84.70863, 84.70853, 84.70872, 84.70996, 84.70972, 84.7105, 84.71104, 
    84.7114, 84.71166, 84.71162, 84.71155, 84.71119, 84.71085, 84.7106, 
    84.71044, 84.71029, 84.70986, 84.70965, 84.70875, 84.70883, 84.70869, 
    84.70856, 84.70835, 84.70838, 84.70829, 84.70869, 84.70843, 84.70931, 
    84.70875, 84.71026, 84.71072, 84.71094, 84.71112, 84.71159, 84.71127, 
    84.7114, 84.71109, 84.7109, 84.71099, 84.71044, 84.71065, 84.70963, 
    84.71004, 84.70858, 84.70881, 84.70852, 84.70867, 84.70842, 84.70864, 
    84.70826, 84.70818, 84.70823, 84.70802, 84.70866, 84.7084, 84.711, 
    84.71098, 84.71091, 84.71123, 84.71124, 84.71154, 84.71127, 84.71117, 
    84.71089, 84.71073, 84.71059, 84.71027, 84.70995, 84.70953, 84.70879, 
    84.70861, 84.70872, 84.70862, 84.70873, 84.70879, 84.70821, 84.70853, 
    84.70805, 84.70808, 84.70829, 84.70807, 84.71097, 84.71106, 84.71137, 
    84.71113, 84.71157, 84.71132, 84.71118, 84.71065, 84.71053, 84.71043, 
    84.71024, 84.70999, 84.70961, 84.70884, 84.70856, 84.70857, 84.70857, 
    84.7085, 84.70866, 84.70848, 84.70845, 84.70853, 84.70808, 84.70821, 
    84.70808, 84.70815, 84.71103, 84.71088, 84.71096, 84.71082, 84.71092, 
    84.71047, 84.71034, 84.70979, 84.71, 84.70966, 84.70996, 84.70991, 
    84.70965, 84.70995, 84.7093, 84.70974, 84.7085, 84.70937, 84.70848, 
    84.70856, 84.70843, 84.70831, 84.70817, 84.70791, 84.70797, 84.70776, 
    84.71067, 84.71049, 84.7105, 84.71032, 84.71019, 84.70992, 84.70951, 
    84.70966, 84.70939, 84.70934, 84.70975, 84.7095, 84.71037, 84.71022, 
    84.71031, 84.71066, 84.70963, 84.71012, 84.70879, 84.70948, 84.70833, 
    84.70868, 84.708, 84.70773, 84.70747, 84.70719, 84.7104, 84.71052, 
    84.7103, 84.71002, 84.70978, 84.70947, 84.70943, 84.70938, 84.70879, 
    84.70867, 84.70937, 84.70865, 84.71019, 84.70959, 84.71056, 84.71024, 
    84.71004, 84.71012, 84.70968, 84.70958, 84.70875, 84.70939, 84.7078, 
    84.70829, 84.70698, 84.70733, 84.71056, 84.7104, 84.70987, 84.71011, 
    84.70945, 84.7093, 84.70873, 84.70857, 84.70856, 84.70847, 84.70862, 
    84.70847, 84.70947, 84.70878, 84.70992, 84.70975, 84.70982, 84.70992, 
    84.70964, 84.70936, 84.70935, 84.70882, 84.70859, 84.70944, 84.70774, 
    84.70851, 84.71022, 84.70994, 84.70989, 84.71, 84.70931, 84.70955, 
    84.70847, 84.70864, 84.70836, 84.7085, 84.70852, 84.70869, 84.70881, 
    84.70954, 84.70979, 84.70998, 84.70994, 84.70972, 84.70934, 84.70856, 
    84.70863, 84.70838, 84.7095, 84.70877, 84.70932, 84.7086, 84.70966, 
    84.70869, 84.70981, 84.70975, 84.70956, 84.70875, 84.70866, 84.70858, 
    84.70863, 84.70934, 84.70937, 84.70956, 84.70962, 84.70976, 84.70988, 
    84.70977, 84.70966, 84.70934, 84.70861, 84.70831, 84.70824, 84.70791, 
    84.70818, 84.70774, 84.70811, 84.70747, 84.70866, 84.70812, 84.70955, 
    84.70943, 84.7088, 84.70836, 84.7086, 84.70832, 84.70938, 84.70972, 
    84.7098, 84.70997, 84.7098, 84.70982, 84.70965, 84.7097, 84.70932, 
    84.70953, 84.70852, 84.70832, 84.70778, 84.70747, 84.70715, 84.70702, 
    84.70698, 84.70696 ;

 RH2M_R =
  84.7115, 84.71105, 84.71114, 84.71078, 84.71098, 84.71075, 84.71141, 
    84.71104, 84.71127, 84.71146, 84.71015, 84.71077, 84.70958, 84.70992, 
    84.70865, 84.70963, 84.70854, 84.70866, 84.7083, 84.7084, 84.70796, 
    84.70825, 84.70773, 84.70803, 84.70798, 84.70827, 84.71064, 84.71023, 
    84.71066, 84.7106, 84.71063, 84.71098, 84.71116, 84.71153, 84.71146, 
    84.71119, 84.71058, 84.71078, 84.71027, 84.71029, 84.70979, 84.71001, 
    84.70879, 84.70944, 84.7084, 84.70855, 84.7084, 84.70845, 84.7084, 
    84.70863, 84.70853, 84.70872, 84.70996, 84.70972, 84.7105, 84.71104, 
    84.7114, 84.71166, 84.71162, 84.71155, 84.71119, 84.71085, 84.7106, 
    84.71044, 84.71029, 84.70986, 84.70965, 84.70875, 84.70883, 84.70869, 
    84.70856, 84.70835, 84.70838, 84.70829, 84.70869, 84.70843, 84.70931, 
    84.70875, 84.71026, 84.71072, 84.71094, 84.71112, 84.71159, 84.71127, 
    84.7114, 84.71109, 84.7109, 84.71099, 84.71044, 84.71065, 84.70963, 
    84.71004, 84.70858, 84.70881, 84.70852, 84.70867, 84.70842, 84.70864, 
    84.70826, 84.70818, 84.70823, 84.70802, 84.70866, 84.7084, 84.711, 
    84.71098, 84.71091, 84.71123, 84.71124, 84.71154, 84.71127, 84.71117, 
    84.71089, 84.71073, 84.71059, 84.71027, 84.70995, 84.70953, 84.70879, 
    84.70861, 84.70872, 84.70862, 84.70873, 84.70879, 84.70821, 84.70853, 
    84.70805, 84.70808, 84.70829, 84.70807, 84.71097, 84.71106, 84.71137, 
    84.71113, 84.71157, 84.71132, 84.71118, 84.71065, 84.71053, 84.71043, 
    84.71024, 84.70999, 84.70961, 84.70884, 84.70856, 84.70857, 84.70857, 
    84.7085, 84.70866, 84.70848, 84.70845, 84.70853, 84.70808, 84.70821, 
    84.70808, 84.70815, 84.71103, 84.71088, 84.71096, 84.71082, 84.71092, 
    84.71047, 84.71034, 84.70979, 84.71, 84.70966, 84.70996, 84.70991, 
    84.70965, 84.70995, 84.7093, 84.70974, 84.7085, 84.70937, 84.70848, 
    84.70856, 84.70843, 84.70831, 84.70817, 84.70791, 84.70797, 84.70776, 
    84.71067, 84.71049, 84.7105, 84.71032, 84.71019, 84.70992, 84.70951, 
    84.70966, 84.70939, 84.70934, 84.70975, 84.7095, 84.71037, 84.71022, 
    84.71031, 84.71066, 84.70963, 84.71012, 84.70879, 84.70948, 84.70833, 
    84.70868, 84.708, 84.70773, 84.70747, 84.70719, 84.7104, 84.71052, 
    84.7103, 84.71002, 84.70978, 84.70947, 84.70943, 84.70938, 84.70879, 
    84.70867, 84.70937, 84.70865, 84.71019, 84.70959, 84.71056, 84.71024, 
    84.71004, 84.71012, 84.70968, 84.70958, 84.70875, 84.70939, 84.7078, 
    84.70829, 84.70698, 84.70733, 84.71056, 84.7104, 84.70987, 84.71011, 
    84.70945, 84.7093, 84.70873, 84.70857, 84.70856, 84.70847, 84.70862, 
    84.70847, 84.70947, 84.70878, 84.70992, 84.70975, 84.70982, 84.70992, 
    84.70964, 84.70936, 84.70935, 84.70882, 84.70859, 84.70944, 84.70774, 
    84.70851, 84.71022, 84.70994, 84.70989, 84.71, 84.70931, 84.70955, 
    84.70847, 84.70864, 84.70836, 84.7085, 84.70852, 84.70869, 84.70881, 
    84.70954, 84.70979, 84.70998, 84.70994, 84.70972, 84.70934, 84.70856, 
    84.70863, 84.70838, 84.7095, 84.70877, 84.70932, 84.7086, 84.70966, 
    84.70869, 84.70981, 84.70975, 84.70956, 84.70875, 84.70866, 84.70858, 
    84.70863, 84.70934, 84.70937, 84.70956, 84.70962, 84.70976, 84.70988, 
    84.70977, 84.70966, 84.70934, 84.70861, 84.70831, 84.70824, 84.70791, 
    84.70818, 84.70774, 84.70811, 84.70747, 84.70866, 84.70812, 84.70955, 
    84.70943, 84.7088, 84.70836, 84.7086, 84.70832, 84.70938, 84.70972, 
    84.7098, 84.70997, 84.7098, 84.70982, 84.70965, 84.7097, 84.70932, 
    84.70953, 84.70852, 84.70832, 84.70778, 84.70747, 84.70715, 84.70702, 
    84.70698, 84.70696 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004631352, 0.0004650756, 0.0004646982, 0.0004662633, 0.000465395, 
    0.0004664197, 0.0004635283, 0.0004651524, 0.0004641155, 0.0004633093, 
    0.0004692999, 0.0004663326, 0.0004723805, 0.0004704885, 0.0004752402, 
    0.0004720861, 0.000475876, 0.0004751488, 0.0004773365, 0.0004767097, 
    0.000479508, 0.0004776256, 0.000480958, 0.0004790583, 0.0004793555, 
    0.0004775633, 0.00046693, 0.000468931, 0.0004668114, 0.0004670967, 
    0.0004669685, 0.0004654128, 0.0004646289, 0.0004629863, 0.0004632844, 
    0.0004644907, 0.0004672246, 0.0004662963, 0.000468635, 0.0004685821, 
    0.0004711855, 0.0004700117, 0.0004743867, 0.0004731432, 0.0004767358, 
    0.0004758323, 0.0004766933, 0.0004764321, 0.0004766965, 0.0004753716, 
    0.0004759392, 0.0004747731, 0.0004702322, 0.0004715672, 0.0004675852, 
    0.0004651906, 0.0004635993, 0.0004624703, 0.0004626298, 0.0004629341, 
    0.0004644976, 0.0004659673, 0.0004670872, 0.0004678364, 0.0004685744, 
    0.0004708091, 0.0004719912, 0.0004746381, 0.0004741602, 0.0004749695, 
    0.0004757424, 0.0004770401, 0.0004768264, 0.0004773982, 0.0004749477, 
    0.0004765764, 0.0004738875, 0.000474623, 0.0004687764, 0.0004665469, 
    0.0004656, 0.0004647703, 0.0004627525, 0.000464146, 0.0004635966, 
    0.0004649032, 0.0004657334, 0.0004653226, 0.0004678568, 0.0004668715, 
    0.0004720612, 0.000469826, 0.0004756523, 0.0004742581, 0.0004759862, 
    0.0004751044, 0.0004766153, 0.0004752554, 0.0004776108, 0.0004781238, 
    0.0004777731, 0.0004791193, 0.0004751797, 0.0004766928, 0.0004653115, 
    0.0004653785, 0.0004656904, 0.0004643189, 0.000464235, 0.0004629778, 
    0.0004640962, 0.0004645726, 0.0004657813, 0.0004664964, 0.000467176, 
    0.0004686704, 0.0004703393, 0.0004726725, 0.0004743485, 0.0004754717, 
    0.0004747828, 0.0004753909, 0.0004747111, 0.0004743923, 0.0004779315, 
    0.0004759443, 0.0004789256, 0.0004787606, 0.0004774114, 0.000478779, 
    0.0004654254, 0.0004650399, 0.0004637018, 0.0004647489, 0.0004628408, 
    0.0004639089, 0.0004645231, 0.0004668923, 0.0004674125, 0.0004678952, 
    0.0004688482, 0.0004700714, 0.000472217, 0.0004740835, 0.0004757871, 
    0.0004756621, 0.0004757061, 0.0004760867, 0.0004751438, 0.0004762413, 
    0.0004764255, 0.0004759438, 0.0004787383, 0.00047794, 0.0004787568, 
    0.0004782369, 0.0004651651, 0.0004658135, 0.000465463, 0.000466122, 
    0.0004656577, 0.0004677219, 0.0004683407, 0.0004712357, 0.0004700474, 
    0.0004719383, 0.0004702393, 0.0004705404, 0.0004720002, 0.0004703309, 
    0.0004739806, 0.0004715065, 0.0004761014, 0.0004736314, 0.000476256, 
    0.0004757793, 0.0004765684, 0.0004772753, 0.0004781642, 0.0004798048, 
    0.0004794248, 0.0004807966, 0.0004667801, 0.0004676212, 0.000467547, 
    0.000468427, 0.0004690778, 0.0004704884, 0.0004727505, 0.0004718997, 
    0.0004734612, 0.0004737748, 0.0004714021, 0.000472859, 0.0004681835, 
    0.000468939, 0.000468489, 0.0004668457, 0.0004720955, 0.0004694015, 
    0.0004743755, 0.0004729163, 0.0004771743, 0.000475057, 0.0004792156, 
    0.0004809936, 0.0004826659, 0.0004846208, 0.00046808, 0.0004675084, 
    0.0004685315, 0.0004699473, 0.0004712602, 0.000473006, 0.0004731844, 
    0.0004735114, 0.0004743583, 0.0004750705, 0.0004736148, 0.0004752488, 
    0.0004691145, 0.0004723293, 0.0004672918, 0.000468809, 0.000469863, 
    0.0004694005, 0.0004718018, 0.0004723677, 0.0004746674, 0.0004734785, 
    0.0004805548, 0.0004774244, 0.0004861086, 0.0004836823, 0.0004673087, 
    0.0004680777, 0.0004707544, 0.0004694809, 0.0004731223, 0.0004740186, 
    0.0004747469, 0.0004756783, 0.0004757786, 0.0004763305, 0.0004754261, 
    0.0004762946, 0.0004730091, 0.0004744773, 0.0004704477, 0.0004714286, 
    0.0004709772, 0.0004704822, 0.0004720096, 0.0004736372, 0.0004736716, 
    0.0004741934, 0.0004756644, 0.000473136, 0.000480959, 0.0004761285, 
    0.0004689163, 0.0004703979, 0.0004706091, 0.0004700353, 0.0004739286, 
    0.000472518, 0.000476317, 0.0004752902, 0.0004769723, 0.0004761364, 
    0.0004760133, 0.0004749397, 0.0004742712, 0.0004725823, 0.0004712078, 
    0.0004701178, 0.0004703711, 0.0004715685, 0.0004737365, 0.0004757872, 
    0.000475338, 0.0004768437, 0.0004728571, 0.000474529, 0.0004738828, 
    0.0004755674, 0.000471877, 0.0004750213, 0.0004710732, 0.0004714192, 
    0.0004724898, 0.0004746434, 0.0004751193, 0.0004756281, 0.000475314, 
    0.0004737919, 0.0004735423, 0.0004724634, 0.0004721656, 0.0004713433, 
    0.0004706626, 0.0004712846, 0.0004719376, 0.000473792, 0.000475463, 
    0.0004772847, 0.0004777303, 0.000479859, 0.0004781265, 0.0004809857, 
    0.0004785553, 0.0004827618, 0.000475203, 0.0004784844, 0.0004725385, 
    0.000473179, 0.0004743378, 0.0004769949, 0.0004755601, 0.0004772379, 
    0.0004735325, 0.00047161, 0.0004711122, 0.0004701841, 0.0004711333, 
    0.0004710561, 0.0004719644, 0.0004716725, 0.0004738534, 0.0004726819, 
    0.0004760096, 0.0004772239, 0.0004806523, 0.0004827537, 0.0004848923, 
    0.0004858364, 0.0004861237, 0.0004862437 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.113897e-14, 3.122322e-14, 3.120686e-14, 3.127474e-14, 3.12371e-14, 
    3.128154e-14, 3.115607e-14, 3.122655e-14, 3.118157e-14, 3.114657e-14, 
    3.14063e-14, 3.127778e-14, 3.15397e-14, 3.145788e-14, 3.166328e-14, 
    3.152695e-14, 3.169076e-14, 3.165938e-14, 3.175384e-14, 3.172679e-14, 
    3.184741e-14, 3.176631e-14, 3.190991e-14, 3.182807e-14, 3.184087e-14, 
    3.176363e-14, 3.130368e-14, 3.13903e-14, 3.129854e-14, 3.13109e-14, 
    3.130536e-14, 3.123787e-14, 3.120382e-14, 3.113255e-14, 3.11455e-14, 
    3.119785e-14, 3.131646e-14, 3.127623e-14, 3.137763e-14, 3.137534e-14, 
    3.148805e-14, 3.143725e-14, 3.162646e-14, 3.157275e-14, 3.172792e-14, 
    3.168892e-14, 3.172608e-14, 3.171482e-14, 3.172623e-14, 3.166902e-14, 
    3.169353e-14, 3.164318e-14, 3.144676e-14, 3.150454e-14, 3.133209e-14, 
    3.122818e-14, 3.115916e-14, 3.111012e-14, 3.111706e-14, 3.113027e-14, 
    3.119816e-14, 3.126196e-14, 3.131054e-14, 3.134302e-14, 3.137501e-14, 
    3.147169e-14, 3.152288e-14, 3.163731e-14, 3.161669e-14, 3.165163e-14, 
    3.168504e-14, 3.174105e-14, 3.173184e-14, 3.17565e-14, 3.165073e-14, 
    3.172103e-14, 3.160495e-14, 3.16367e-14, 3.138361e-14, 3.128709e-14, 
    3.124595e-14, 3.121e-14, 3.112239e-14, 3.118289e-14, 3.115905e-14, 
    3.121579e-14, 3.125182e-14, 3.1234e-14, 3.134391e-14, 3.130119e-14, 
    3.152591e-14, 3.14292e-14, 3.168114e-14, 3.162092e-14, 3.169557e-14, 
    3.165749e-14, 3.172272e-14, 3.166402e-14, 3.176568e-14, 3.178779e-14, 
    3.177268e-14, 3.183074e-14, 3.166076e-14, 3.172607e-14, 3.12335e-14, 
    3.123641e-14, 3.124995e-14, 3.11904e-14, 3.118676e-14, 3.113219e-14, 
    3.118076e-14, 3.120143e-14, 3.125391e-14, 3.128492e-14, 3.13144e-14, 
    3.137917e-14, 3.145142e-14, 3.155238e-14, 3.162483e-14, 3.167336e-14, 
    3.164361e-14, 3.166988e-14, 3.164051e-14, 3.162675e-14, 3.17795e-14, 
    3.169376e-14, 3.182239e-14, 3.181529e-14, 3.175708e-14, 3.181609e-14, 
    3.123845e-14, 3.122173e-14, 3.116363e-14, 3.12091e-14, 3.112624e-14, 
    3.117262e-14, 3.119927e-14, 3.130207e-14, 3.132466e-14, 3.134557e-14, 
    3.138688e-14, 3.143985e-14, 3.153269e-14, 3.161337e-14, 3.168698e-14, 
    3.168159e-14, 3.168349e-14, 3.169992e-14, 3.165921e-14, 3.17066e-14, 
    3.171454e-14, 3.169376e-14, 3.181433e-14, 3.177991e-14, 3.181513e-14, 
    3.179272e-14, 3.122717e-14, 3.12553e-14, 3.12401e-14, 3.126868e-14, 
    3.124854e-14, 3.133803e-14, 3.136484e-14, 3.149021e-14, 3.14388e-14, 
    3.152062e-14, 3.144713e-14, 3.146015e-14, 3.152325e-14, 3.145111e-14, 
    3.160892e-14, 3.150192e-14, 3.170055e-14, 3.159381e-14, 3.170724e-14, 
    3.168666e-14, 3.172073e-14, 3.175122e-14, 3.178958e-14, 3.186028e-14, 
    3.184392e-14, 3.190302e-14, 3.129723e-14, 3.133368e-14, 3.133049e-14, 
    3.136863e-14, 3.139682e-14, 3.145791e-14, 3.155577e-14, 3.151899e-14, 
    3.158652e-14, 3.160006e-14, 3.149747e-14, 3.156046e-14, 3.135807e-14, 
    3.139079e-14, 3.137133e-14, 3.130009e-14, 3.152744e-14, 3.141083e-14, 
    3.162602e-14, 3.156298e-14, 3.174687e-14, 3.165544e-14, 3.183491e-14, 
    3.191145e-14, 3.198351e-14, 3.206753e-14, 3.135358e-14, 3.132882e-14, 
    3.137317e-14, 3.143444e-14, 3.149131e-14, 3.156682e-14, 3.157455e-14, 
    3.158868e-14, 3.162528e-14, 3.165604e-14, 3.159313e-14, 3.166375e-14, 
    3.139834e-14, 3.153756e-14, 3.131944e-14, 3.138516e-14, 3.143084e-14, 
    3.141082e-14, 3.151479e-14, 3.153927e-14, 3.163863e-14, 3.15873e-14, 
    3.189255e-14, 3.175763e-14, 3.21315e-14, 3.202719e-14, 3.132016e-14, 
    3.13535e-14, 3.146941e-14, 3.141428e-14, 3.157187e-14, 3.16106e-14, 
    3.164207e-14, 3.168227e-14, 3.168663e-14, 3.171044e-14, 3.167141e-14, 
    3.170891e-14, 3.156698e-14, 3.163043e-14, 3.145619e-14, 3.149862e-14, 
    3.147911e-14, 3.145769e-14, 3.152379e-14, 3.159412e-14, 3.159565e-14, 
    3.161816e-14, 3.168157e-14, 3.15725e-14, 3.190989e-14, 3.170164e-14, 
    3.138985e-14, 3.145395e-14, 3.146314e-14, 3.143831e-14, 3.160672e-14, 
    3.154573e-14, 3.170986e-14, 3.166554e-14, 3.173816e-14, 3.170208e-14, 
    3.169677e-14, 3.165041e-14, 3.162153e-14, 3.154852e-14, 3.148907e-14, 
    3.144192e-14, 3.145288e-14, 3.150468e-14, 3.159843e-14, 3.168701e-14, 
    3.16676e-14, 3.173264e-14, 3.156045e-14, 3.163267e-14, 3.160477e-14, 
    3.167754e-14, 3.1518e-14, 3.165379e-14, 3.148325e-14, 3.149822e-14, 
    3.154452e-14, 3.163755e-14, 3.165816e-14, 3.168012e-14, 3.166658e-14, 
    3.160081e-14, 3.159004e-14, 3.154341e-14, 3.153051e-14, 3.149496e-14, 
    3.146551e-14, 3.149241e-14, 3.152065e-14, 3.160085e-14, 3.167301e-14, 
    3.175165e-14, 3.177089e-14, 3.186257e-14, 3.178791e-14, 3.191104e-14, 
    3.180631e-14, 3.198755e-14, 3.166169e-14, 3.180329e-14, 3.154664e-14, 
    3.157434e-14, 3.162436e-14, 3.173908e-14, 3.16772e-14, 3.174958e-14, 
    3.158962e-14, 3.150645e-14, 3.148496e-14, 3.144478e-14, 3.148587e-14, 
    3.148253e-14, 3.152184e-14, 3.150922e-14, 3.160351e-14, 3.155288e-14, 
    3.169663e-14, 3.174902e-14, 3.189682e-14, 3.198727e-14, 3.207928e-14, 
    3.211984e-14, 3.213219e-14, 3.213735e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.035367e-14, 1.038171e-14, 1.037626e-14, 1.039886e-14, 1.038633e-14, 
    1.040112e-14, 1.035936e-14, 1.038282e-14, 1.036785e-14, 1.03562e-14, 
    1.044264e-14, 1.039987e-14, 1.048704e-14, 1.045981e-14, 1.052818e-14, 
    1.04828e-14, 1.053732e-14, 1.052688e-14, 1.055831e-14, 1.054931e-14, 
    1.058946e-14, 1.056247e-14, 1.061026e-14, 1.058302e-14, 1.058728e-14, 
    1.056158e-14, 1.040849e-14, 1.043732e-14, 1.040678e-14, 1.041089e-14, 
    1.040905e-14, 1.038659e-14, 1.037525e-14, 1.035153e-14, 1.035584e-14, 
    1.037327e-14, 1.041274e-14, 1.039936e-14, 1.04331e-14, 1.043234e-14, 
    1.046985e-14, 1.045295e-14, 1.051592e-14, 1.049804e-14, 1.054969e-14, 
    1.053671e-14, 1.054908e-14, 1.054533e-14, 1.054913e-14, 1.053008e-14, 
    1.053824e-14, 1.052149e-14, 1.045611e-14, 1.047534e-14, 1.041795e-14, 
    1.038336e-14, 1.036039e-14, 1.034407e-14, 1.034638e-14, 1.035078e-14, 
    1.037337e-14, 1.039461e-14, 1.041077e-14, 1.042158e-14, 1.043223e-14, 
    1.046441e-14, 1.048144e-14, 1.051953e-14, 1.051267e-14, 1.05243e-14, 
    1.053542e-14, 1.055406e-14, 1.055099e-14, 1.05592e-14, 1.0524e-14, 
    1.05474e-14, 1.050876e-14, 1.051933e-14, 1.043509e-14, 1.040297e-14, 
    1.038928e-14, 1.037731e-14, 1.034815e-14, 1.036829e-14, 1.036035e-14, 
    1.037924e-14, 1.039123e-14, 1.03853e-14, 1.042188e-14, 1.040766e-14, 
    1.048245e-14, 1.045027e-14, 1.053412e-14, 1.051408e-14, 1.053892e-14, 
    1.052625e-14, 1.054796e-14, 1.052842e-14, 1.056226e-14, 1.056962e-14, 
    1.056459e-14, 1.058391e-14, 1.052734e-14, 1.054907e-14, 1.038513e-14, 
    1.03861e-14, 1.039061e-14, 1.037079e-14, 1.036958e-14, 1.035141e-14, 
    1.036758e-14, 1.037446e-14, 1.039193e-14, 1.040225e-14, 1.041206e-14, 
    1.043361e-14, 1.045766e-14, 1.049126e-14, 1.051538e-14, 1.053153e-14, 
    1.052163e-14, 1.053037e-14, 1.05206e-14, 1.051602e-14, 1.056686e-14, 
    1.053832e-14, 1.058113e-14, 1.057877e-14, 1.05594e-14, 1.057903e-14, 
    1.038678e-14, 1.038122e-14, 1.036188e-14, 1.037701e-14, 1.034944e-14, 
    1.036487e-14, 1.037374e-14, 1.040795e-14, 1.041547e-14, 1.042243e-14, 
    1.043618e-14, 1.045381e-14, 1.048471e-14, 1.051156e-14, 1.053606e-14, 
    1.053427e-14, 1.05349e-14, 1.054037e-14, 1.052682e-14, 1.054259e-14, 
    1.054523e-14, 1.053832e-14, 1.057845e-14, 1.056699e-14, 1.057872e-14, 
    1.057126e-14, 1.038302e-14, 1.039239e-14, 1.038733e-14, 1.039684e-14, 
    1.039014e-14, 1.041992e-14, 1.042885e-14, 1.047057e-14, 1.045346e-14, 
    1.048069e-14, 1.045623e-14, 1.046057e-14, 1.048157e-14, 1.045756e-14, 
    1.051008e-14, 1.047447e-14, 1.054058e-14, 1.050505e-14, 1.05428e-14, 
    1.053596e-14, 1.05473e-14, 1.055744e-14, 1.057021e-14, 1.059374e-14, 
    1.05883e-14, 1.060797e-14, 1.040634e-14, 1.041847e-14, 1.041741e-14, 
    1.043011e-14, 1.043949e-14, 1.045982e-14, 1.049239e-14, 1.048015e-14, 
    1.050263e-14, 1.050713e-14, 1.047299e-14, 1.049395e-14, 1.042659e-14, 
    1.043748e-14, 1.0431e-14, 1.04073e-14, 1.048296e-14, 1.044415e-14, 
    1.051577e-14, 1.049479e-14, 1.0556e-14, 1.052557e-14, 1.05853e-14, 
    1.061077e-14, 1.063476e-14, 1.066272e-14, 1.04251e-14, 1.041686e-14, 
    1.043162e-14, 1.045201e-14, 1.047094e-14, 1.049607e-14, 1.049864e-14, 
    1.050335e-14, 1.051553e-14, 1.052577e-14, 1.050483e-14, 1.052833e-14, 
    1.043999e-14, 1.048633e-14, 1.041374e-14, 1.043561e-14, 1.045081e-14, 
    1.044415e-14, 1.047875e-14, 1.04869e-14, 1.051997e-14, 1.050289e-14, 
    1.060448e-14, 1.055958e-14, 1.068401e-14, 1.06493e-14, 1.041398e-14, 
    1.042507e-14, 1.046365e-14, 1.04453e-14, 1.049775e-14, 1.051064e-14, 
    1.052112e-14, 1.05345e-14, 1.053595e-14, 1.054387e-14, 1.053088e-14, 
    1.054336e-14, 1.049612e-14, 1.051724e-14, 1.045925e-14, 1.047337e-14, 
    1.046688e-14, 1.045975e-14, 1.048175e-14, 1.050516e-14, 1.050566e-14, 
    1.051316e-14, 1.053426e-14, 1.049796e-14, 1.061025e-14, 1.054094e-14, 
    1.043717e-14, 1.04585e-14, 1.046156e-14, 1.04533e-14, 1.050935e-14, 
    1.048905e-14, 1.054368e-14, 1.052893e-14, 1.05531e-14, 1.054109e-14, 
    1.053932e-14, 1.052389e-14, 1.051428e-14, 1.048998e-14, 1.047019e-14, 
    1.04545e-14, 1.045815e-14, 1.047539e-14, 1.050659e-14, 1.053607e-14, 
    1.052961e-14, 1.055126e-14, 1.049395e-14, 1.051799e-14, 1.05087e-14, 
    1.053292e-14, 1.047982e-14, 1.052502e-14, 1.046825e-14, 1.047324e-14, 
    1.048865e-14, 1.051961e-14, 1.052647e-14, 1.053378e-14, 1.052927e-14, 
    1.050738e-14, 1.05038e-14, 1.048828e-14, 1.048399e-14, 1.047215e-14, 
    1.046235e-14, 1.047131e-14, 1.04807e-14, 1.05074e-14, 1.053141e-14, 
    1.055759e-14, 1.056399e-14, 1.059451e-14, 1.056966e-14, 1.061064e-14, 
    1.057578e-14, 1.06361e-14, 1.052765e-14, 1.057477e-14, 1.048935e-14, 
    1.049857e-14, 1.051522e-14, 1.05534e-14, 1.053281e-14, 1.05569e-14, 
    1.050366e-14, 1.047598e-14, 1.046882e-14, 1.045545e-14, 1.046913e-14, 
    1.046802e-14, 1.04811e-14, 1.04769e-14, 1.050828e-14, 1.049143e-14, 
    1.053927e-14, 1.055671e-14, 1.06059e-14, 1.063601e-14, 1.066663e-14, 
    1.068014e-14, 1.068424e-14, 1.068596e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.36479e-11, -8.401602e-11, -8.394446e-11, -8.424138e-11, -8.407667e-11, 
    -8.427109e-11, -8.372253e-11, -8.403064e-11, -8.383395e-11, 
    -8.368103e-11, -8.48176e-11, -8.425462e-11, -8.540234e-11, -8.504331e-11, 
    -8.59452e-11, -8.534647e-11, -8.606592e-11, -8.592792e-11, -8.634325e-11, 
    -8.622426e-11, -8.675553e-11, -8.639817e-11, -8.703091e-11, 
    -8.667018e-11, -8.672662e-11, -8.638638e-11, -8.436791e-11, 
    -8.474751e-11, -8.434542e-11, -8.439955e-11, -8.437526e-11, 
    -8.408008e-11, -8.393132e-11, -8.361976e-11, -8.367632e-11, 
    -8.390515e-11, -8.442389e-11, -8.42478e-11, -8.469158e-11, -8.468156e-11, 
    -8.517562e-11, -8.495286e-11, -8.578324e-11, -8.554724e-11, 
    -8.622923e-11, -8.605772e-11, -8.622118e-11, -8.617161e-11, 
    -8.622182e-11, -8.597028e-11, -8.607805e-11, -8.58567e-11, -8.499458e-11, 
    -8.524795e-11, -8.449226e-11, -8.403788e-11, -8.373605e-11, 
    -8.352187e-11, -8.355215e-11, -8.360987e-11, -8.390649e-11, 
    -8.418536e-11, -8.439788e-11, -8.454005e-11, -8.468012e-11, 
    -8.510413e-11, -8.532852e-11, -8.583097e-11, -8.574029e-11, 
    -8.589391e-11, -8.604065e-11, -8.628704e-11, -8.624649e-11, 
    -8.635504e-11, -8.588985e-11, -8.619902e-11, -8.568864e-11, 
    -8.582823e-11, -8.471823e-11, -8.42953e-11, -8.411557e-11, -8.395822e-11, 
    -8.357543e-11, -8.383978e-11, -8.373557e-11, -8.398348e-11, 
    -8.414101e-11, -8.40631e-11, -8.454393e-11, -8.4357e-11, -8.534182e-11, 
    -8.491763e-11, -8.602354e-11, -8.57589e-11, -8.608697e-11, -8.591956e-11, 
    -8.62064e-11, -8.594825e-11, -8.639544e-11, -8.649281e-11, -8.642627e-11, 
    -8.668188e-11, -8.593394e-11, -8.622118e-11, -8.406091e-11, 
    -8.407362e-11, -8.413282e-11, -8.38726e-11, -8.385669e-11, -8.361821e-11, 
    -8.38304e-11, -8.392076e-11, -8.415013e-11, -8.428581e-11, -8.441479e-11, 
    -8.469837e-11, -8.501506e-11, -8.545791e-11, -8.577605e-11, 
    -8.598931e-11, -8.585854e-11, -8.5974e-11, -8.584494e-11, -8.578444e-11, 
    -8.645633e-11, -8.607906e-11, -8.664511e-11, -8.661379e-11, 
    -8.635762e-11, -8.661732e-11, -8.408254e-11, -8.400942e-11, 
    -8.375555e-11, -8.395423e-11, -8.359224e-11, -8.379487e-11, 
    -8.391138e-11, -8.436091e-11, -8.445967e-11, -8.455125e-11, 
    -8.473213e-11, -8.496426e-11, -8.537147e-11, -8.572577e-11, 
    -8.604919e-11, -8.602549e-11, -8.603383e-11, -8.610609e-11, 
    -8.592712e-11, -8.613547e-11, -8.617045e-11, -8.607901e-11, 
    -8.660959e-11, -8.645801e-11, -8.661313e-11, -8.651443e-11, 
    -8.403318e-11, -8.415622e-11, -8.408974e-11, -8.421476e-11, 
    -8.412668e-11, -8.451834e-11, -8.463576e-11, -8.518519e-11, 
    -8.495969e-11, -8.531856e-11, -8.499614e-11, -8.505328e-11, 
    -8.533028e-11, -8.501357e-11, -8.570624e-11, -8.523664e-11, -8.61089e-11, 
    -8.563997e-11, -8.613828e-11, -8.604779e-11, -8.619762e-11, -8.63318e-11, 
    -8.650061e-11, -8.68121e-11, -8.673997e-11, -8.700046e-11, -8.433965e-11, 
    -8.449923e-11, -8.448518e-11, -8.465218e-11, -8.477569e-11, 
    -8.504339e-11, -8.547274e-11, -8.531129e-11, -8.560769e-11, 
    -8.566719e-11, -8.521688e-11, -8.549337e-11, -8.460604e-11, 
    -8.474941e-11, -8.466404e-11, -8.435224e-11, -8.53485e-11, -8.483722e-11, 
    -8.578131e-11, -8.550435e-11, -8.631267e-11, -8.591068e-11, 
    -8.670027e-11, -8.703782e-11, -8.735548e-11, -8.772675e-11, 
    -8.458632e-11, -8.447789e-11, -8.467204e-11, -8.494067e-11, -8.51899e-11, 
    -8.552124e-11, -8.555514e-11, -8.561721e-11, -8.5778e-11, -8.591318e-11, 
    -8.563684e-11, -8.594707e-11, -8.478267e-11, -8.539287e-11, 
    -8.443689e-11, -8.472478e-11, -8.492484e-11, -8.483707e-11, 
    -8.529283e-11, -8.540025e-11, -8.583675e-11, -8.561111e-11, 
    -8.695452e-11, -8.636016e-11, -8.800941e-11, -8.754852e-11, -8.444e-11, 
    -8.458595e-11, -8.50939e-11, -8.485222e-11, -8.554336e-11, -8.571348e-11, 
    -8.585177e-11, -8.602857e-11, -8.604764e-11, -8.615239e-11, 
    -8.598074e-11, -8.614561e-11, -8.552194e-11, -8.580064e-11, 
    -8.503583e-11, -8.522198e-11, -8.513634e-11, -8.504241e-11, 
    -8.533232e-11, -8.56412e-11, -8.564779e-11, -8.574683e-11, -8.602595e-11, 
    -8.554615e-11, -8.703125e-11, -8.611412e-11, -8.474509e-11, 
    -8.502622e-11, -8.506636e-11, -8.495746e-11, -8.569643e-11, 
    -8.542868e-11, -8.614984e-11, -8.595493e-11, -8.627428e-11, 
    -8.611559e-11, -8.609224e-11, -8.588843e-11, -8.576154e-11, 
    -8.544095e-11, -8.518011e-11, -8.497326e-11, -8.502135e-11, 
    -8.524857e-11, -8.566009e-11, -8.604938e-11, -8.59641e-11, -8.625001e-11, 
    -8.549324e-11, -8.581057e-11, -8.568793e-11, -8.600772e-11, -8.5307e-11, 
    -8.590374e-11, -8.515447e-11, -8.522016e-11, -8.542336e-11, 
    -8.583211e-11, -8.592252e-11, -8.601908e-11, -8.59595e-11, -8.567053e-11, 
    -8.562319e-11, -8.541842e-11, -8.536188e-11, -8.520586e-11, 
    -8.507668e-11, -8.519471e-11, -8.531865e-11, -8.567065e-11, 
    -8.598787e-11, -8.633372e-11, -8.641834e-11, -8.682247e-11, 
    -8.649351e-11, -8.703636e-11, -8.657487e-11, -8.737373e-11, -8.59383e-11, 
    -8.656127e-11, -8.543261e-11, -8.55542e-11, -8.577413e-11, -8.627855e-11, 
    -8.600622e-11, -8.63247e-11, -8.562134e-11, -8.525642e-11, -8.516199e-11, 
    -8.498583e-11, -8.516602e-11, -8.515137e-11, -8.532378e-11, 
    -8.526838e-11, -8.568234e-11, -8.545997e-11, -8.609166e-11, 
    -8.632218e-11, -8.697316e-11, -8.737224e-11, -8.777846e-11, -8.79578e-11, 
    -8.801238e-11, -8.80352e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.016063e-12, -2.024934e-12, -2.023209e-12, -2.030364e-12, -2.026395e-12, 
    -2.03108e-12, -2.017861e-12, -2.025286e-12, -2.020546e-12, -2.016862e-12, 
    -2.044249e-12, -2.030683e-12, -2.058339e-12, -2.049687e-12, 
    -2.071419e-12, -2.056992e-12, -2.074329e-12, -2.071003e-12, 
    -2.081011e-12, -2.078144e-12, -2.090945e-12, -2.082335e-12, 
    -2.097581e-12, -2.088889e-12, -2.090249e-12, -2.08205e-12, -2.033413e-12, 
    -2.04256e-12, -2.032871e-12, -2.034175e-12, -2.03359e-12, -2.026477e-12, 
    -2.022892e-12, -2.015385e-12, -2.016748e-12, -2.022262e-12, 
    -2.034762e-12, -2.030518e-12, -2.041212e-12, -2.04097e-12, -2.052875e-12, 
    -2.047508e-12, -2.067517e-12, -2.06183e-12, -2.078264e-12, -2.074131e-12, 
    -2.078069e-12, -2.076875e-12, -2.078085e-12, -2.072024e-12, 
    -2.074621e-12, -2.069287e-12, -2.048513e-12, -2.054619e-12, 
    -2.036409e-12, -2.02546e-12, -2.018187e-12, -2.013026e-12, -2.013756e-12, 
    -2.015147e-12, -2.022294e-12, -2.029014e-12, -2.034135e-12, -2.03756e-12, 
    -2.040936e-12, -2.051153e-12, -2.05656e-12, -2.068667e-12, -2.066482e-12, 
    -2.070184e-12, -2.07372e-12, -2.079657e-12, -2.078679e-12, -2.081295e-12, 
    -2.070086e-12, -2.077536e-12, -2.065237e-12, -2.068601e-12, 
    -2.041854e-12, -2.031663e-12, -2.027332e-12, -2.023541e-12, 
    -2.014317e-12, -2.020687e-12, -2.018176e-12, -2.024149e-12, 
    -2.027945e-12, -2.026068e-12, -2.037654e-12, -2.03315e-12, -2.05688e-12, 
    -2.046659e-12, -2.073307e-12, -2.06693e-12, -2.074836e-12, -2.070802e-12, 
    -2.077714e-12, -2.071493e-12, -2.082269e-12, -2.084615e-12, 
    -2.083011e-12, -2.089171e-12, -2.071148e-12, -2.07807e-12, -2.026015e-12, 
    -2.026321e-12, -2.027748e-12, -2.021478e-12, -2.021094e-12, 
    -2.015348e-12, -2.020461e-12, -2.022638e-12, -2.028165e-12, 
    -2.031434e-12, -2.034542e-12, -2.041375e-12, -2.049007e-12, 
    -2.059678e-12, -2.067344e-12, -2.072483e-12, -2.069331e-12, 
    -2.072114e-12, -2.069004e-12, -2.067546e-12, -2.083736e-12, 
    -2.074645e-12, -2.088285e-12, -2.08753e-12, -2.081357e-12, -2.087615e-12, 
    -2.026536e-12, -2.024774e-12, -2.018657e-12, -2.023444e-12, 
    -2.014722e-12, -2.019604e-12, -2.022412e-12, -2.033244e-12, 
    -2.035624e-12, -2.037831e-12, -2.042189e-12, -2.047783e-12, 
    -2.057595e-12, -2.066132e-12, -2.073925e-12, -2.073354e-12, 
    -2.073555e-12, -2.075297e-12, -2.070984e-12, -2.076005e-12, 
    -2.076847e-12, -2.074644e-12, -2.087429e-12, -2.083777e-12, 
    -2.087514e-12, -2.085136e-12, -2.025347e-12, -2.028312e-12, -2.02671e-12, 
    -2.029722e-12, -2.0276e-12, -2.037037e-12, -2.039867e-12, -2.053106e-12, 
    -2.047673e-12, -2.05632e-12, -2.048551e-12, -2.049928e-12, -2.056602e-12, 
    -2.048971e-12, -2.065661e-12, -2.054346e-12, -2.075364e-12, 
    -2.064065e-12, -2.076072e-12, -2.073892e-12, -2.077502e-12, 
    -2.080735e-12, -2.084803e-12, -2.092309e-12, -2.090571e-12, 
    -2.096847e-12, -2.032732e-12, -2.036577e-12, -2.036238e-12, 
    -2.040263e-12, -2.043239e-12, -2.049689e-12, -2.060035e-12, 
    -2.056145e-12, -2.063287e-12, -2.064721e-12, -2.05387e-12, -2.060532e-12, 
    -2.039151e-12, -2.042605e-12, -2.040548e-12, -2.033035e-12, 
    -2.057041e-12, -2.044721e-12, -2.067471e-12, -2.060797e-12, 
    -2.080274e-12, -2.070588e-12, -2.089614e-12, -2.097748e-12, 
    -2.105402e-12, -2.114348e-12, -2.038676e-12, -2.036063e-12, 
    -2.040741e-12, -2.047214e-12, -2.05322e-12, -2.061204e-12, -2.06202e-12, 
    -2.063516e-12, -2.067391e-12, -2.070648e-12, -2.063989e-12, 
    -2.071465e-12, -2.043407e-12, -2.058111e-12, -2.035075e-12, 
    -2.042012e-12, -2.046833e-12, -2.044718e-12, -2.0557e-12, -2.058288e-12, 
    -2.068806e-12, -2.063369e-12, -2.09574e-12, -2.081418e-12, -2.121159e-12, 
    -2.110053e-12, -2.03515e-12, -2.038667e-12, -2.050906e-12, -2.045083e-12, 
    -2.061737e-12, -2.065836e-12, -2.069168e-12, -2.073428e-12, 
    -2.073888e-12, -2.076412e-12, -2.072276e-12, -2.076249e-12, 
    -2.061221e-12, -2.067936e-12, -2.049507e-12, -2.053993e-12, 
    -2.051929e-12, -2.049666e-12, -2.056652e-12, -2.064094e-12, 
    -2.064253e-12, -2.06664e-12, -2.073365e-12, -2.061804e-12, -2.097589e-12, 
    -2.07549e-12, -2.042501e-12, -2.049276e-12, -2.050243e-12, -2.047619e-12, 
    -2.065425e-12, -2.058973e-12, -2.076351e-12, -2.071654e-12, 
    -2.079349e-12, -2.075525e-12, -2.074963e-12, -2.070052e-12, 
    -2.066994e-12, -2.059269e-12, -2.052984e-12, -2.047999e-12, 
    -2.049158e-12, -2.054634e-12, -2.064549e-12, -2.07393e-12, -2.071875e-12, 
    -2.078764e-12, -2.060529e-12, -2.068176e-12, -2.06522e-12, -2.072926e-12, 
    -2.056041e-12, -2.07042e-12, -2.052366e-12, -2.053949e-12, -2.058845e-12, 
    -2.068694e-12, -2.070873e-12, -2.0732e-12, -2.071764e-12, -2.064801e-12, 
    -2.06366e-12, -2.058726e-12, -2.057364e-12, -2.053604e-12, -2.050492e-12, 
    -2.053335e-12, -2.056322e-12, -2.064804e-12, -2.072448e-12, 
    -2.080781e-12, -2.082821e-12, -2.092558e-12, -2.084632e-12, 
    -2.097712e-12, -2.086592e-12, -2.105842e-12, -2.071253e-12, 
    -2.086265e-12, -2.059068e-12, -2.061998e-12, -2.067298e-12, 
    -2.079452e-12, -2.07289e-12, -2.080564e-12, -2.063616e-12, -2.054822e-12, 
    -2.052547e-12, -2.048302e-12, -2.052644e-12, -2.052291e-12, 
    -2.056446e-12, -2.055111e-12, -2.065086e-12, -2.059727e-12, 
    -2.074949e-12, -2.080503e-12, -2.09619e-12, -2.105806e-12, -2.115594e-12, 
    -2.119915e-12, -2.121231e-12, -2.12178e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.363431e-15, 3.37254e-15, 3.370771e-15, 3.378111e-15, 3.374041e-15, 
    3.378846e-15, 3.36528e-15, 3.372901e-15, 3.368038e-15, 3.364254e-15, 
    3.392335e-15, 3.378439e-15, 3.406758e-15, 3.397911e-15, 3.42012e-15, 
    3.40538e-15, 3.42309e-15, 3.419698e-15, 3.429911e-15, 3.426986e-15, 
    3.440028e-15, 3.43126e-15, 3.446786e-15, 3.437937e-15, 3.439321e-15, 
    3.43097e-15, 3.38124e-15, 3.390605e-15, 3.380684e-15, 3.38202e-15, 
    3.381422e-15, 3.374124e-15, 3.370443e-15, 3.362737e-15, 3.364137e-15, 
    3.369798e-15, 3.382621e-15, 3.378272e-15, 3.389235e-15, 3.388988e-15, 
    3.401174e-15, 3.395681e-15, 3.416139e-15, 3.410331e-15, 3.427109e-15, 
    3.422891e-15, 3.42691e-15, 3.425692e-15, 3.426926e-15, 3.42074e-15, 
    3.423391e-15, 3.417947e-15, 3.39671e-15, 3.402956e-15, 3.384311e-15, 
    3.373076e-15, 3.365614e-15, 3.360313e-15, 3.361063e-15, 3.362491e-15, 
    3.369831e-15, 3.376729e-15, 3.381982e-15, 3.385493e-15, 3.388952e-15, 
    3.399405e-15, 3.404939e-15, 3.417311e-15, 3.415082e-15, 3.41886e-15, 
    3.422472e-15, 3.428528e-15, 3.427532e-15, 3.430199e-15, 3.418763e-15, 
    3.426364e-15, 3.413814e-15, 3.417246e-15, 3.389881e-15, 3.379446e-15, 
    3.374998e-15, 3.371111e-15, 3.361639e-15, 3.368181e-15, 3.365602e-15, 
    3.371737e-15, 3.375632e-15, 3.373707e-15, 3.385589e-15, 3.380971e-15, 
    3.405267e-15, 3.39481e-15, 3.422051e-15, 3.41554e-15, 3.423611e-15, 
    3.419494e-15, 3.426546e-15, 3.4202e-15, 3.431192e-15, 3.433582e-15, 
    3.431949e-15, 3.438226e-15, 3.419847e-15, 3.426909e-15, 3.373652e-15, 
    3.373966e-15, 3.37543e-15, 3.368992e-15, 3.368599e-15, 3.362698e-15, 
    3.36795e-15, 3.370184e-15, 3.375859e-15, 3.379212e-15, 3.382398e-15, 
    3.389401e-15, 3.397213e-15, 3.408129e-15, 3.415962e-15, 3.42121e-15, 
    3.417993e-15, 3.420833e-15, 3.417658e-15, 3.41617e-15, 3.432686e-15, 
    3.423415e-15, 3.437323e-15, 3.436555e-15, 3.430262e-15, 3.436642e-15, 
    3.374187e-15, 3.372379e-15, 3.366097e-15, 3.371014e-15, 3.362055e-15, 
    3.36707e-15, 3.369951e-15, 3.381065e-15, 3.383508e-15, 3.385769e-15, 
    3.390235e-15, 3.395963e-15, 3.406e-15, 3.414723e-15, 3.422682e-15, 
    3.4221e-15, 3.422305e-15, 3.424081e-15, 3.419679e-15, 3.424803e-15, 
    3.425662e-15, 3.423415e-15, 3.436452e-15, 3.43273e-15, 3.436538e-15, 
    3.434115e-15, 3.372967e-15, 3.376009e-15, 3.374365e-15, 3.377455e-15, 
    3.375277e-15, 3.384953e-15, 3.387852e-15, 3.401407e-15, 3.395849e-15, 
    3.404696e-15, 3.396749e-15, 3.398157e-15, 3.404979e-15, 3.397179e-15, 
    3.414242e-15, 3.402674e-15, 3.42415e-15, 3.412608e-15, 3.424872e-15, 
    3.422648e-15, 3.426331e-15, 3.429628e-15, 3.433776e-15, 3.44142e-15, 
    3.439651e-15, 3.446041e-15, 3.380542e-15, 3.384483e-15, 3.384138e-15, 
    3.388262e-15, 3.39131e-15, 3.397915e-15, 3.408496e-15, 3.404519e-15, 
    3.41182e-15, 3.413284e-15, 3.402193e-15, 3.409003e-15, 3.387121e-15, 
    3.390658e-15, 3.388554e-15, 3.380852e-15, 3.405433e-15, 3.392825e-15, 
    3.416091e-15, 3.409274e-15, 3.429158e-15, 3.419272e-15, 3.438676e-15, 
    3.446952e-15, 3.454744e-15, 3.463828e-15, 3.386635e-15, 3.383958e-15, 
    3.388752e-15, 3.395378e-15, 3.401526e-15, 3.40969e-15, 3.410526e-15, 
    3.412054e-15, 3.416011e-15, 3.419337e-15, 3.412535e-15, 3.420171e-15, 
    3.391474e-15, 3.406527e-15, 3.382944e-15, 3.390049e-15, 3.394988e-15, 
    3.392824e-15, 3.404065e-15, 3.406711e-15, 3.417454e-15, 3.411904e-15, 
    3.444909e-15, 3.430321e-15, 3.470745e-15, 3.459467e-15, 3.383022e-15, 
    3.386627e-15, 3.399158e-15, 3.393198e-15, 3.410236e-15, 3.414424e-15, 
    3.417826e-15, 3.422173e-15, 3.422644e-15, 3.425218e-15, 3.420999e-15, 
    3.425053e-15, 3.409707e-15, 3.416568e-15, 3.397729e-15, 3.402317e-15, 
    3.400207e-15, 3.397891e-15, 3.405038e-15, 3.412642e-15, 3.412807e-15, 
    3.415242e-15, 3.422097e-15, 3.410305e-15, 3.446784e-15, 3.424267e-15, 
    3.390556e-15, 3.397487e-15, 3.398481e-15, 3.395796e-15, 3.414004e-15, 
    3.40741e-15, 3.425156e-15, 3.420364e-15, 3.428216e-15, 3.424314e-15, 
    3.42374e-15, 3.418728e-15, 3.415605e-15, 3.407712e-15, 3.401285e-15, 
    3.396186e-15, 3.397372e-15, 3.402972e-15, 3.413107e-15, 3.422685e-15, 
    3.420587e-15, 3.427619e-15, 3.409001e-15, 3.41681e-15, 3.413793e-15, 
    3.421662e-15, 3.404412e-15, 3.419093e-15, 3.400654e-15, 3.402273e-15, 
    3.407279e-15, 3.417338e-15, 3.419567e-15, 3.42194e-15, 3.420476e-15, 
    3.413365e-15, 3.412201e-15, 3.407159e-15, 3.405764e-15, 3.401921e-15, 
    3.398736e-15, 3.401645e-15, 3.404698e-15, 3.41337e-15, 3.421172e-15, 
    3.429675e-15, 3.431755e-15, 3.441668e-15, 3.433595e-15, 3.446908e-15, 
    3.435584e-15, 3.45518e-15, 3.419948e-15, 3.435258e-15, 3.407508e-15, 
    3.410503e-15, 3.415912e-15, 3.428316e-15, 3.421625e-15, 3.429451e-15, 
    3.412155e-15, 3.403163e-15, 3.400839e-15, 3.396495e-15, 3.400939e-15, 
    3.400577e-15, 3.404827e-15, 3.403462e-15, 3.413657e-15, 3.408183e-15, 
    3.423725e-15, 3.42939e-15, 3.44537e-15, 3.45515e-15, 3.465098e-15, 
    3.469484e-15, 3.470819e-15, 3.471377e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.757486e-09, -8.795996e-09, -8.788509e-09, -8.819569e-09, -8.802339e-09, 
    -8.822678e-09, -8.765293e-09, -8.797524e-09, -8.776949e-09, 
    -8.760953e-09, -8.879847e-09, -8.820955e-09, -8.941015e-09, 
    -8.903458e-09, -8.997802e-09, -8.935171e-09, -9.01043e-09, -8.995993e-09, 
    -9.03944e-09, -9.026993e-09, -9.082567e-09, -9.045185e-09, -9.111373e-09, 
    -9.073639e-09, -9.079542e-09, -9.043952e-09, -8.832806e-09, 
    -8.872515e-09, -8.830453e-09, -8.836116e-09, -8.833575e-09, 
    -8.802695e-09, -8.787135e-09, -8.754543e-09, -8.76046e-09, -8.784397e-09, 
    -8.838662e-09, -8.820241e-09, -8.866664e-09, -8.865616e-09, 
    -8.917298e-09, -8.893996e-09, -8.98086e-09, -8.956172e-09, -9.027513e-09, 
    -9.009572e-09, -9.026671e-09, -9.021486e-09, -9.026738e-09, 
    -9.000425e-09, -9.011699e-09, -8.988544e-09, -8.89836e-09, -8.924865e-09, 
    -8.845814e-09, -8.798281e-09, -8.766707e-09, -8.744302e-09, -8.74747e-09, 
    -8.753508e-09, -8.784538e-09, -8.81371e-09, -8.835941e-09, -8.850813e-09, 
    -8.865465e-09, -8.90982e-09, -8.933293e-09, -8.985853e-09, -8.976366e-09, 
    -8.992436e-09, -9.007787e-09, -9.033561e-09, -9.029318e-09, 
    -9.040673e-09, -8.992012e-09, -9.024353e-09, -8.970964e-09, 
    -8.985566e-09, -8.869453e-09, -8.825211e-09, -8.806409e-09, 
    -8.789948e-09, -8.749906e-09, -8.777558e-09, -8.766658e-09, 
    -8.792591e-09, -8.80907e-09, -8.800919e-09, -8.851219e-09, -8.831664e-09, 
    -8.934684e-09, -8.890311e-09, -9.005997e-09, -8.978313e-09, 
    -9.012632e-09, -8.995119e-09, -9.025126e-09, -8.99812e-09, -9.044899e-09, 
    -9.055086e-09, -9.048125e-09, -9.074863e-09, -8.996624e-09, 
    -9.026671e-09, -8.800691e-09, -8.80202e-09, -8.808213e-09, -8.780992e-09, 
    -8.779327e-09, -8.75438e-09, -8.776578e-09, -8.786031e-09, -8.810025e-09, 
    -8.824218e-09, -8.837709e-09, -8.867374e-09, -8.900503e-09, 
    -8.946828e-09, -8.980108e-09, -9.002417e-09, -8.988737e-09, 
    -9.000814e-09, -8.987313e-09, -8.980986e-09, -9.051269e-09, 
    -9.011805e-09, -9.071017e-09, -9.06774e-09, -9.040943e-09, -9.06811e-09, 
    -8.802954e-09, -8.795304e-09, -8.768748e-09, -8.789531e-09, 
    -8.751664e-09, -8.772861e-09, -8.785048e-09, -8.832074e-09, 
    -8.842404e-09, -8.851985e-09, -8.870906e-09, -8.895189e-09, 
    -8.937786e-09, -8.974848e-09, -9.00868e-09, -9.006201e-09, -9.007073e-09, 
    -9.014632e-09, -8.99591e-09, -9.017706e-09, -9.021364e-09, -9.011799e-09, 
    -9.067302e-09, -9.051445e-09, -9.067671e-09, -9.057346e-09, 
    -8.797791e-09, -8.810662e-09, -8.803707e-09, -8.816786e-09, 
    -8.807572e-09, -8.848541e-09, -8.860825e-09, -8.9183e-09, -8.894711e-09, 
    -8.932251e-09, -8.898524e-09, -8.9045e-09, -8.933477e-09, -8.900346e-09, 
    -8.972805e-09, -8.923682e-09, -9.014926e-09, -8.965873e-09, -9.018e-09, 
    -9.008533e-09, -9.024206e-09, -9.038243e-09, -9.055901e-09, 
    -9.088485e-09, -9.08094e-09, -9.108188e-09, -8.829849e-09, -8.846543e-09, 
    -8.845073e-09, -8.862543e-09, -8.875463e-09, -8.903466e-09, 
    -8.948379e-09, -8.93149e-09, -8.962496e-09, -8.96872e-09, -8.921615e-09, 
    -8.950537e-09, -8.857715e-09, -8.872713e-09, -8.863783e-09, 
    -8.831166e-09, -8.935383e-09, -8.8819e-09, -8.980658e-09, -8.951686e-09, 
    -9.036242e-09, -8.994191e-09, -9.076786e-09, -9.112096e-09, 
    -9.145324e-09, -9.18416e-09, -8.855654e-09, -8.84431e-09, -8.86462e-09, 
    -8.892721e-09, -8.918792e-09, -8.953453e-09, -8.956999e-09, 
    -8.963492e-09, -8.980311e-09, -8.994452e-09, -8.965547e-09, 
    -8.997997e-09, -8.876193e-09, -8.940025e-09, -8.840022e-09, 
    -8.870137e-09, -8.891065e-09, -8.881884e-09, -8.929559e-09, 
    -8.940797e-09, -8.986458e-09, -8.962854e-09, -9.103382e-09, 
    -9.041209e-09, -9.213728e-09, -9.165517e-09, -8.840347e-09, 
    -8.855614e-09, -8.908749e-09, -8.883468e-09, -8.955766e-09, 
    -8.973562e-09, -8.988028e-09, -9.006522e-09, -9.008518e-09, 
    -9.019475e-09, -9.00152e-09, -9.018766e-09, -8.953527e-09, -8.98268e-09, 
    -8.902675e-09, -8.922148e-09, -8.91319e-09, -8.903363e-09, -8.93369e-09, 
    -8.966001e-09, -8.966691e-09, -8.977051e-09, -9.006248e-09, 
    -8.956059e-09, -9.111409e-09, -9.015471e-09, -8.872262e-09, 
    -8.901671e-09, -8.905869e-09, -8.894478e-09, -8.971778e-09, -8.94377e-09, 
    -9.019208e-09, -8.998819e-09, -9.032226e-09, -9.015626e-09, 
    -9.013183e-09, -8.991863e-09, -8.978589e-09, -8.945054e-09, 
    -8.917768e-09, -8.89613e-09, -8.901161e-09, -8.92493e-09, -8.967977e-09, 
    -9.0087e-09, -8.99978e-09, -9.029686e-09, -8.950524e-09, -8.983719e-09, 
    -8.97089e-09, -9.004342e-09, -8.931042e-09, -8.993465e-09, -8.915086e-09, 
    -8.921957e-09, -8.943214e-09, -8.985971e-09, -8.995429e-09, -9.00553e-09, 
    -8.999297e-09, -8.96907e-09, -8.964117e-09, -8.942697e-09, -8.936784e-09, 
    -8.920461e-09, -8.906949e-09, -8.919295e-09, -8.932261e-09, 
    -8.969082e-09, -9.002265e-09, -9.038443e-09, -9.047295e-09, 
    -9.089568e-09, -9.055158e-09, -9.111943e-09, -9.063668e-09, 
    -9.147233e-09, -8.99708e-09, -9.062246e-09, -8.944181e-09, -8.9569e-09, 
    -8.979907e-09, -9.032671e-09, -9.004185e-09, -9.0375e-09, -8.963923e-09, 
    -8.925751e-09, -8.915872e-09, -8.897445e-09, -8.916294e-09, 
    -8.914761e-09, -8.932797e-09, -8.927001e-09, -8.970304e-09, 
    -8.947044e-09, -9.013123e-09, -9.037236e-09, -9.105332e-09, 
    -9.147078e-09, -9.18957e-09, -9.208329e-09, -9.214039e-09, -9.216426e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039174e-10, -1.043745e-10, -1.042856e-10, -1.046543e-10, -1.044498e-10, 
    -1.046912e-10, -1.040101e-10, -1.043927e-10, -1.041484e-10, 
    -1.039585e-10, -1.053699e-10, -1.046708e-10, -1.06096e-10, -1.056502e-10, 
    -1.067701e-10, -1.060266e-10, -1.069201e-10, -1.067487e-10, 
    -1.072645e-10, -1.071167e-10, -1.077764e-10, -1.073326e-10, 
    -1.081184e-10, -1.076704e-10, -1.077405e-10, -1.07318e-10, -1.048115e-10, 
    -1.052829e-10, -1.047835e-10, -1.048508e-10, -1.048206e-10, -1.04454e-10, 
    -1.042693e-10, -1.038824e-10, -1.039527e-10, -1.042368e-10, -1.04881e-10, 
    -1.046623e-10, -1.052134e-10, -1.05201e-10, -1.058145e-10, -1.055378e-10, 
    -1.06569e-10, -1.062759e-10, -1.071229e-10, -1.069099e-10, -1.071129e-10, 
    -1.070513e-10, -1.071137e-10, -1.068013e-10, -1.069351e-10, 
    -1.066603e-10, -1.055897e-10, -1.059043e-10, -1.049659e-10, 
    -1.044016e-10, -1.040268e-10, -1.037609e-10, -1.037985e-10, 
    -1.038702e-10, -1.042385e-10, -1.045848e-10, -1.048487e-10, 
    -1.050252e-10, -1.051992e-10, -1.057257e-10, -1.060043e-10, 
    -1.066283e-10, -1.065157e-10, -1.067064e-10, -1.068887e-10, 
    -1.071946e-10, -1.071443e-10, -1.072791e-10, -1.067014e-10, 
    -1.070853e-10, -1.064515e-10, -1.066249e-10, -1.052465e-10, 
    -1.047213e-10, -1.044981e-10, -1.043027e-10, -1.038274e-10, 
    -1.041556e-10, -1.040262e-10, -1.043341e-10, -1.045297e-10, 
    -1.044329e-10, -1.0503e-10, -1.047979e-10, -1.060209e-10, -1.054941e-10, 
    -1.068674e-10, -1.065388e-10, -1.069462e-10, -1.067383e-10, 
    -1.070945e-10, -1.067739e-10, -1.073293e-10, -1.074502e-10, 
    -1.073676e-10, -1.07685e-10, -1.067562e-10, -1.071129e-10, -1.044302e-10, 
    -1.04446e-10, -1.045195e-10, -1.041964e-10, -1.041766e-10, -1.038805e-10, 
    -1.04144e-10, -1.042562e-10, -1.04541e-10, -1.047095e-10, -1.048697e-10, 
    -1.052218e-10, -1.056151e-10, -1.06165e-10, -1.065601e-10, -1.068249e-10, 
    -1.066625e-10, -1.068059e-10, -1.066456e-10, -1.065705e-10, 
    -1.074049e-10, -1.069364e-10, -1.076393e-10, -1.076004e-10, 
    -1.072823e-10, -1.076048e-10, -1.044571e-10, -1.043663e-10, -1.04051e-10, 
    -1.042978e-10, -1.038483e-10, -1.040999e-10, -1.042446e-10, 
    -1.048028e-10, -1.049254e-10, -1.050391e-10, -1.052637e-10, -1.05552e-10, 
    -1.060577e-10, -1.064976e-10, -1.068993e-10, -1.068699e-10, 
    -1.068802e-10, -1.069699e-10, -1.067477e-10, -1.070064e-10, 
    -1.070499e-10, -1.069363e-10, -1.075952e-10, -1.07407e-10, -1.075996e-10, 
    -1.07477e-10, -1.043958e-10, -1.045486e-10, -1.04466e-10, -1.046213e-10, 
    -1.045119e-10, -1.049983e-10, -1.051441e-10, -1.058264e-10, 
    -1.055463e-10, -1.05992e-10, -1.055916e-10, -1.056625e-10, -1.060065e-10, 
    -1.056132e-10, -1.064734e-10, -1.058902e-10, -1.069734e-10, 
    -1.063911e-10, -1.070099e-10, -1.068975e-10, -1.070836e-10, 
    -1.072502e-10, -1.074599e-10, -1.078467e-10, -1.077571e-10, 
    -1.080806e-10, -1.047764e-10, -1.049745e-10, -1.049571e-10, 
    -1.051645e-10, -1.053179e-10, -1.056503e-10, -1.061834e-10, 
    -1.059829e-10, -1.06351e-10, -1.064249e-10, -1.058657e-10, -1.062091e-10, 
    -1.051072e-10, -1.052852e-10, -1.051792e-10, -1.04792e-10, -1.060292e-10, 
    -1.053943e-10, -1.065666e-10, -1.062227e-10, -1.072265e-10, 
    -1.067273e-10, -1.077078e-10, -1.08127e-10, -1.085215e-10, -1.089825e-10, 
    -1.050827e-10, -1.04948e-10, -1.051891e-10, -1.055227e-10, -1.058322e-10, 
    -1.062437e-10, -1.062858e-10, -1.063628e-10, -1.065625e-10, 
    -1.067304e-10, -1.063872e-10, -1.067725e-10, -1.053265e-10, 
    -1.060843e-10, -1.048971e-10, -1.052546e-10, -1.055031e-10, 
    -1.053941e-10, -1.0596e-10, -1.060934e-10, -1.066355e-10, -1.063553e-10, 
    -1.080235e-10, -1.072855e-10, -1.093336e-10, -1.087612e-10, -1.04901e-10, 
    -1.050822e-10, -1.05713e-10, -1.054129e-10, -1.062711e-10, -1.064824e-10, 
    -1.066541e-10, -1.068737e-10, -1.068974e-10, -1.070274e-10, 
    -1.068143e-10, -1.07019e-10, -1.062445e-10, -1.065906e-10, -1.056409e-10, 
    -1.05872e-10, -1.057657e-10, -1.056491e-10, -1.060091e-10, -1.063926e-10, 
    -1.064008e-10, -1.065238e-10, -1.068704e-10, -1.062746e-10, 
    -1.081188e-10, -1.069799e-10, -1.052798e-10, -1.05629e-10, -1.056788e-10, 
    -1.055436e-10, -1.064612e-10, -1.061287e-10, -1.070243e-10, 
    -1.067822e-10, -1.071788e-10, -1.069817e-10, -1.069527e-10, 
    -1.066996e-10, -1.065421e-10, -1.06144e-10, -1.0582e-10, -1.055632e-10, 
    -1.056229e-10, -1.059051e-10, -1.064161e-10, -1.068995e-10, 
    -1.067936e-10, -1.071487e-10, -1.062089e-10, -1.06603e-10, -1.064507e-10, 
    -1.068478e-10, -1.059776e-10, -1.067187e-10, -1.057882e-10, 
    -1.058698e-10, -1.061221e-10, -1.066297e-10, -1.06742e-10, -1.068619e-10, 
    -1.067879e-10, -1.064291e-10, -1.063703e-10, -1.06116e-10, -1.060458e-10, 
    -1.05852e-10, -1.056916e-10, -1.058382e-10, -1.059921e-10, -1.064292e-10, 
    -1.068231e-10, -1.072526e-10, -1.073577e-10, -1.078596e-10, 
    -1.074511e-10, -1.081252e-10, -1.075521e-10, -1.085441e-10, 
    -1.067616e-10, -1.075352e-10, -1.061336e-10, -1.062846e-10, 
    -1.065577e-10, -1.071841e-10, -1.068459e-10, -1.072414e-10, -1.06368e-10, 
    -1.059148e-10, -1.057976e-10, -1.055788e-10, -1.058025e-10, 
    -1.057844e-10, -1.059985e-10, -1.059297e-10, -1.064437e-10, 
    -1.061676e-10, -1.06952e-10, -1.072383e-10, -1.080467e-10, -1.085423e-10, 
    -1.090468e-10, -1.092695e-10, -1.093373e-10, -1.093656e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.619456e-12, -8.657389e-12, -8.650015e-12, -8.68061e-12, -8.663638e-12, 
    -8.683673e-12, -8.627146e-12, -8.658896e-12, -8.638627e-12, 
    -8.622871e-12, -8.739987e-12, -8.681975e-12, -8.800241e-12, 
    -8.763244e-12, -8.85618e-12, -8.794484e-12, -8.868619e-12, -8.854399e-12, 
    -8.897197e-12, -8.884936e-12, -8.93968e-12, -8.902856e-12, -8.968056e-12, 
    -8.930886e-12, -8.9367e-12, -8.901642e-12, -8.693649e-12, -8.732765e-12, 
    -8.691332e-12, -8.69691e-12, -8.694406e-12, -8.663989e-12, -8.648661e-12, 
    -8.616556e-12, -8.622384e-12, -8.645964e-12, -8.699418e-12, 
    -8.681272e-12, -8.727001e-12, -8.725969e-12, -8.776879e-12, 
    -8.753925e-12, -8.839492e-12, -8.815172e-12, -8.885448e-12, 
    -8.867775e-12, -8.884618e-12, -8.87951e-12, -8.884685e-12, -8.858764e-12, 
    -8.869869e-12, -8.847061e-12, -8.758223e-12, -8.784333e-12, 
    -8.706463e-12, -8.659641e-12, -8.628539e-12, -8.606469e-12, -8.60959e-12, 
    -8.615537e-12, -8.646102e-12, -8.674839e-12, -8.696738e-12, 
    -8.711387e-12, -8.72582e-12, -8.769512e-12, -8.792634e-12, -8.84441e-12, 
    -8.835065e-12, -8.850895e-12, -8.866016e-12, -8.891405e-12, 
    -8.887226e-12, -8.898412e-12, -8.850476e-12, -8.882334e-12, 
    -8.829742e-12, -8.844127e-12, -8.729748e-12, -8.686167e-12, 
    -8.667646e-12, -8.651432e-12, -8.611988e-12, -8.639227e-12, 
    -8.628489e-12, -8.654035e-12, -8.670268e-12, -8.662239e-12, 
    -8.711787e-12, -8.692524e-12, -8.794005e-12, -8.750294e-12, 
    -8.864252e-12, -8.836982e-12, -8.870789e-12, -8.853538e-12, 
    -8.883096e-12, -8.856494e-12, -8.902574e-12, -8.912608e-12, 
    -8.905751e-12, -8.93209e-12, -8.855019e-12, -8.884618e-12, -8.662015e-12, 
    -8.663324e-12, -8.669424e-12, -8.64261e-12, -8.64097e-12, -8.616397e-12, 
    -8.638261e-12, -8.647572e-12, -8.671208e-12, -8.685189e-12, 
    -8.698479e-12, -8.7277e-12, -8.760334e-12, -8.805967e-12, -8.83875e-12, 
    -8.860726e-12, -8.84725e-12, -8.859147e-12, -8.845849e-12, -8.839615e-12, 
    -8.908849e-12, -8.869973e-12, -8.928303e-12, -8.925074e-12, 
    -8.898678e-12, -8.925439e-12, -8.664243e-12, -8.656708e-12, 
    -8.630549e-12, -8.651021e-12, -8.61372e-12, -8.6346e-12, -8.646605e-12, 
    -8.692927e-12, -8.703104e-12, -8.712541e-12, -8.73118e-12, -8.755099e-12, 
    -8.79706e-12, -8.833568e-12, -8.866896e-12, -8.864453e-12, -8.865313e-12, 
    -8.872758e-12, -8.854317e-12, -8.875786e-12, -8.87939e-12, -8.869968e-12, 
    -8.924642e-12, -8.909022e-12, -8.925006e-12, -8.914836e-12, 
    -8.659158e-12, -8.671836e-12, -8.664985e-12, -8.677867e-12, 
    -8.668792e-12, -8.709149e-12, -8.721249e-12, -8.777865e-12, 
    -8.754629e-12, -8.791608e-12, -8.758385e-12, -8.764272e-12, 
    -8.792816e-12, -8.76018e-12, -8.831556e-12, -8.783167e-12, -8.873048e-12, 
    -8.824728e-12, -8.876076e-12, -8.866751e-12, -8.88219e-12, -8.896018e-12, 
    -8.913413e-12, -8.945509e-12, -8.938077e-12, -8.964918e-12, 
    -8.690736e-12, -8.707181e-12, -8.705732e-12, -8.722942e-12, 
    -8.735669e-12, -8.763253e-12, -8.807496e-12, -8.790859e-12, 
    -8.821401e-12, -8.827532e-12, -8.78113e-12, -8.809621e-12, -8.718186e-12, 
    -8.73296e-12, -8.724163e-12, -8.692034e-12, -8.794693e-12, -8.742009e-12, 
    -8.839292e-12, -8.810752e-12, -8.894046e-12, -8.852623e-12, 
    -8.933985e-12, -8.968768e-12, -9.001502e-12, -9.039759e-12, 
    -8.716155e-12, -8.704981e-12, -8.724988e-12, -8.752669e-12, -8.77835e-12, 
    -8.812493e-12, -8.815986e-12, -8.822383e-12, -8.83895e-12, -8.85288e-12, 
    -8.824406e-12, -8.856372e-12, -8.736387e-12, -8.799266e-12, 
    -8.700758e-12, -8.730422e-12, -8.751037e-12, -8.741993e-12, 
    -8.788957e-12, -8.800026e-12, -8.845005e-12, -8.821753e-12, 
    -8.960184e-12, -8.898939e-12, -9.068885e-12, -9.021393e-12, 
    -8.701078e-12, -8.716116e-12, -8.768457e-12, -8.743554e-12, 
    -8.814772e-12, -8.832303e-12, -8.846553e-12, -8.86477e-12, -8.866736e-12, 
    -8.87753e-12, -8.859843e-12, -8.876831e-12, -8.812566e-12, -8.841284e-12, 
    -8.762474e-12, -8.781657e-12, -8.772831e-12, -8.763152e-12, 
    -8.793026e-12, -8.824854e-12, -8.825533e-12, -8.835739e-12, -8.8645e-12, 
    -8.815061e-12, -8.968091e-12, -8.873586e-12, -8.732516e-12, 
    -8.761484e-12, -8.76562e-12, -8.754399e-12, -8.830545e-12, -8.802955e-12, 
    -8.877267e-12, -8.857182e-12, -8.89009e-12, -8.873738e-12, -8.871332e-12, 
    -8.850329e-12, -8.837255e-12, -8.80422e-12, -8.777342e-12, -8.756026e-12, 
    -8.760982e-12, -8.784397e-12, -8.826801e-12, -8.866915e-12, 
    -8.858128e-12, -8.887589e-12, -8.809608e-12, -8.842307e-12, -8.82967e-12, 
    -8.862622e-12, -8.790416e-12, -8.851907e-12, -8.774699e-12, 
    -8.781469e-12, -8.802408e-12, -8.844526e-12, -8.853843e-12, 
    -8.863793e-12, -8.857652e-12, -8.827878e-12, -8.822999e-12, 
    -8.801898e-12, -8.796072e-12, -8.779994e-12, -8.766684e-12, 
    -8.778846e-12, -8.791618e-12, -8.827889e-12, -8.860576e-12, 
    -8.896214e-12, -8.904935e-12, -8.946577e-12, -8.91268e-12, -8.968618e-12, 
    -8.921063e-12, -9.003382e-12, -8.855469e-12, -8.919662e-12, -8.80336e-12, 
    -8.815889e-12, -8.838552e-12, -8.890529e-12, -8.862467e-12, 
    -8.895285e-12, -8.822807e-12, -8.785205e-12, -8.775474e-12, 
    -8.757322e-12, -8.77589e-12, -8.77438e-12, -8.792146e-12, -8.786437e-12, 
    -8.829094e-12, -8.80618e-12, -8.871272e-12, -8.895025e-12, -8.962106e-12, 
    -9.003229e-12, -9.045087e-12, -9.063567e-12, -9.069192e-12, -9.071543e-12 ;

 SMIN_NH4 =
  0.0004617865, 0.0004637153, 0.0004633402, 0.0004648959, 0.0004640328, 
    0.0004650514, 0.0004621772, 0.0004637917, 0.0004627609, 0.0004619596, 
    0.0004679143, 0.0004649649, 0.0004709763, 0.0004690958, 0.0004738186, 
    0.0004706837, 0.0004744505, 0.0004737278, 0.0004759021, 0.0004752791, 
    0.0004780603, 0.0004761894, 0.0004795013, 0.0004776133, 0.0004779087, 
    0.0004761275, 0.0004655586, 0.0004675476, 0.0004654407, 0.0004657244, 
    0.000465597, 0.0004640505, 0.0004632713, 0.0004616385, 0.0004619348, 
    0.0004631339, 0.0004658515, 0.0004649288, 0.0004672534, 0.0004672009, 
    0.0004697885, 0.0004686218, 0.0004729703, 0.0004717344, 0.000475305, 
    0.0004744071, 0.0004752628, 0.0004750032, 0.000475266, 0.0004739492, 
    0.0004745133, 0.0004733544, 0.0004688411, 0.000470168, 0.0004662099, 
    0.0004638296, 0.0004622479, 0.0004611255, 0.0004612841, 0.0004615866, 
    0.0004631408, 0.0004646017, 0.000465715, 0.0004664596, 0.0004671932, 
    0.0004694144, 0.0004705893, 0.0004732202, 0.0004727452, 0.0004735496, 
    0.0004743177, 0.0004756075, 0.0004753952, 0.0004759634, 0.0004735279, 
    0.0004751466, 0.0004724742, 0.0004732052, 0.000467394, 0.0004651779, 
    0.0004642366, 0.0004634119, 0.0004614061, 0.0004627913, 0.0004622452, 
    0.0004635439, 0.0004643692, 0.0004639609, 0.0004664799, 0.0004655005, 
    0.0004706589, 0.0004684372, 0.0004742282, 0.0004728425, 0.0004745601, 
    0.0004736836, 0.0004751853, 0.0004738337, 0.0004761747, 0.0004766845, 
    0.000476336, 0.000477674, 0.0004737584, 0.0004752623, 0.0004639498, 
    0.0004640164, 0.0004643265, 0.0004629632, 0.0004628797, 0.00046163, 
    0.0004627418, 0.0004632153, 0.0004644169, 0.0004651276, 0.0004658032, 
    0.0004672887, 0.0004689475, 0.0004712665, 0.0004729323, 0.0004740487, 
    0.000473364, 0.0004739684, 0.0004732927, 0.0004729758, 0.0004764934, 
    0.0004745184, 0.0004774814, 0.0004773174, 0.0004759765, 0.0004773357, 
    0.0004640631, 0.0004636798, 0.0004623497, 0.0004633906, 0.0004614938, 
    0.0004625556, 0.0004631661, 0.0004655211, 0.0004660382, 0.0004665181, 
    0.0004674654, 0.0004686812, 0.0004708138, 0.0004726689, 0.0004743621, 
    0.000474238, 0.0004742816, 0.0004746599, 0.0004737228, 0.0004748136, 
    0.0004749967, 0.0004745179, 0.0004772953, 0.0004765019, 0.0004773137, 
    0.000476797, 0.0004638043, 0.0004644489, 0.0004641004, 0.0004647555, 
    0.000464294, 0.0004663458, 0.0004669609, 0.0004698385, 0.0004686573, 
    0.0004705368, 0.000468848, 0.0004691473, 0.0004705983, 0.0004689391, 
    0.0004725666, 0.0004701076, 0.0004746745, 0.0004722196, 0.0004748282, 
    0.0004743544, 0.0004751387, 0.0004758412, 0.0004767247, 0.0004783552, 
    0.0004779775, 0.0004793408, 0.0004654097, 0.0004662457, 0.0004661719, 
    0.0004670467, 0.0004676936, 0.0004690956, 0.0004713441, 0.0004704985, 
    0.0004720505, 0.0004723621, 0.0004700039, 0.0004714519, 0.0004668046, 
    0.0004675556, 0.0004671083, 0.0004654749, 0.0004706931, 0.0004680153, 
    0.0004729592, 0.0004715088, 0.0004757409, 0.0004736365, 0.0004777696, 
    0.0004795366, 0.0004811986, 0.0004831414, 0.0004667018, 0.0004661336, 
    0.0004671506, 0.0004685578, 0.0004698628, 0.000471598, 0.0004717753, 
    0.0004721003, 0.0004729421, 0.0004736499, 0.0004722031, 0.0004738272, 
    0.00046773, 0.0004709254, 0.0004659183, 0.0004674264, 0.000468474, 
    0.0004680143, 0.000470401, 0.0004709635, 0.0004732492, 0.0004720676, 
    0.0004791005, 0.0004759894, 0.0004846199, 0.0004822087, 0.0004659351, 
    0.0004666995, 0.0004693601, 0.0004680942, 0.0004717135, 0.0004726044, 
    0.0004733283, 0.000474254, 0.0004743538, 0.0004749022, 0.0004740034, 
    0.0004748665, 0.0004716011, 0.0004730604, 0.0004690552, 0.0004700301, 
    0.0004695815, 0.0004690895, 0.0004706077, 0.0004722253, 0.0004722596, 
    0.0004727782, 0.0004742402, 0.0004717272, 0.0004795023, 0.0004747015, 
    0.0004675331, 0.0004690057, 0.0004692156, 0.0004686452, 0.000472515, 
    0.000471113, 0.0004748888, 0.0004738682, 0.0004755401, 0.0004747093, 
    0.000474587, 0.0004735199, 0.0004728555, 0.0004711768, 0.0004698107, 
    0.0004687273, 0.0004689791, 0.0004701692, 0.0004723241, 0.0004743622, 
    0.0004739157, 0.0004754123, 0.00047145, 0.0004731118, 0.0004724695, 
    0.0004741438, 0.0004704758, 0.0004736011, 0.0004696769, 0.0004700208, 
    0.000471085, 0.0004732255, 0.0004736985, 0.0004742041, 0.0004738919, 
    0.0004723791, 0.0004721311, 0.0004710587, 0.0004707626, 0.0004699454, 
    0.0004692688, 0.000469887, 0.0004705361, 0.0004723792, 0.0004740401, 
    0.0004758506, 0.0004762935, 0.0004784091, 0.0004766872, 0.0004795288, 
    0.0004771134, 0.0004812939, 0.0004737816, 0.0004770429, 0.0004711333, 
    0.0004717699, 0.0004729217, 0.0004755626, 0.0004741366, 0.000475804, 
    0.0004721213, 0.0004702105, 0.0004697157, 0.0004687931, 0.0004697367, 
    0.0004696599, 0.0004705628, 0.0004702725, 0.0004724403, 0.0004712759, 
    0.0004745833, 0.0004757901, 0.0004791974, 0.0004812859, 0.0004834111, 
    0.0004843493, 0.0004846348, 0.0004847542 ;

 SMIN_NH4_vr =
  0.003023245, 0.003028407, 0.003027397, 0.003031558, 0.003029246, 
    0.003031965, 0.003024275, 0.003028591, 0.003025832, 0.003023682, 
    0.003039597, 0.003031719, 0.003047752, 0.003042736, 0.003055305, 
    0.003046965, 0.00305698, 0.003055054, 0.003060828, 0.00305917, 
    0.003066547, 0.003061583, 0.003070358, 0.003065356, 0.003066135, 
    0.003061404, 0.003033325, 0.00303864, 0.003033004, 0.003033763, 
    0.003033418, 0.003029281, 0.003027197, 0.00302282, 0.00302361, 
    0.00302682, 0.003034082, 0.003031611, 0.003037815, 0.003037675, 
    0.00304457, 0.003041461, 0.003053037, 0.003049744, 0.003059235, 
    0.003056845, 0.003059117, 0.003058423, 0.003059117, 0.00305562, 
    0.003057112, 0.003054033, 0.00304208, 0.003045613, 0.003035054, 
    0.00302869, 0.003024452, 0.003021447, 0.003021865, 0.003022677, 
    0.003026833, 0.003030734, 0.003033708, 0.003035692, 0.003037646, 
    0.003043575, 0.0030467, 0.003053695, 0.00305243, 0.003054565, 
    0.003056604, 0.003060026, 0.003059461, 0.003060965, 0.003054491, 
    0.003058793, 0.003051683, 0.003053628, 0.003038217, 0.00303229, 
    0.003029775, 0.003027563, 0.00302219, 0.003025899, 0.003024434, 
    0.003027904, 0.003030109, 0.003029013, 0.003035743, 0.003033123, 
    0.00304688, 0.003040959, 0.003056371, 0.003052682, 0.003057244, 
    0.003054915, 0.003058899, 0.003055308, 0.00306152, 0.003062874, 
    0.003061942, 0.003065492, 0.00305509, 0.003059087, 0.003029001, 
    0.00302918, 0.003030005, 0.003026355, 0.00302613, 0.00302278, 
    0.003025752, 0.00302702, 0.003030228, 0.003032124, 0.003033925, 
    0.003037892, 0.003042314, 0.003048487, 0.003052918, 0.003055881, 
    0.003054059, 0.003055661, 0.003053864, 0.003053016, 0.003062358, 
    0.003057115, 0.003064972, 0.003064538, 0.003060977, 0.003064578, 
    0.003029299, 0.003028269, 0.003024709, 0.003027489, 0.003022409, 
    0.003025253, 0.003026883, 0.003033174, 0.00303455, 0.003035833, 
    0.003038357, 0.003041596, 0.003047278, 0.003052211, 0.00305671, 
    0.003056376, 0.003056491, 0.003057491, 0.003055, 0.003057894, 
    0.003058376, 0.003057105, 0.003064471, 0.003062367, 0.003064516, 
    0.003063141, 0.003028598, 0.003030317, 0.003029382, 0.003031134, 
    0.003029894, 0.003035378, 0.003037016, 0.003044686, 0.003041533, 
    0.003046543, 0.003042035, 0.003042834, 0.003046699, 0.00304227, 
    0.003051931, 0.00304538, 0.003057527, 0.003050998, 0.003057929, 
    0.003056665, 0.003058745, 0.003060611, 0.003062949, 0.003067275, 
    0.003066267, 0.00306988, 0.003032882, 0.003035111, 0.003034912, 
    0.003037243, 0.003038966, 0.003042705, 0.003048692, 0.003046435, 
    0.003050562, 0.003051393, 0.003045107, 0.003048965, 0.003036573, 
    0.003038573, 0.003037377, 0.003033011, 0.00304693, 0.003039788, 
    0.003052954, 0.00304909, 0.003060337, 0.003054748, 0.003065713, 
    0.003070398, 0.003074791, 0.003079925, 0.003036325, 0.003034803, 
    0.003037514, 0.003041271, 0.003044742, 0.003049363, 0.003049831, 
    0.003050691, 0.003052926, 0.003054809, 0.003050959, 0.003055272, 
    0.003039038, 0.003047547, 0.003034189, 0.003038218, 0.003041005, 
    0.003039779, 0.003046137, 0.00304763, 0.003053709, 0.003050566, 
    0.003069235, 0.003060984, 0.003083823, 0.003077454, 0.003034269, 
    0.003036306, 0.0030434, 0.003040025, 0.003049662, 0.003052033, 
    0.003053951, 0.003056413, 0.003056671, 0.003058129, 0.003055734, 
    0.003058028, 0.003049339, 0.003053222, 0.003042554, 0.003045148, 
    0.003043951, 0.003042635, 0.003046676, 0.003050985, 0.00305107, 
    0.003052446, 0.003056336, 0.003049643, 0.003070291, 0.003057551, 
    0.003038527, 0.003042453, 0.003043007, 0.003041486, 0.003051787, 
    0.003048056, 0.003058093, 0.003055377, 0.003059814, 0.003057609, 
    0.003057277, 0.003054442, 0.003052669, 0.003048203, 0.003044558, 
    0.00304167, 0.003042335, 0.003045508, 0.003051239, 0.003056658, 
    0.003055468, 0.003059438, 0.0030489, 0.003053322, 0.003051608, 
    0.003056059, 0.003046362, 0.003054684, 0.00304423, 0.003045142, 
    0.003047973, 0.003053671, 0.00305492, 0.003056265, 0.003055428, 
    0.003051407, 0.003050743, 0.003047883, 0.003047091, 0.003044914, 
    0.003043105, 0.003044753, 0.003046477, 0.003051383, 0.003055796, 
    0.0030606, 0.003061774, 0.003067384, 0.003062815, 0.003070347, 
    0.003063943, 0.003075011, 0.003055153, 0.003063814, 0.003048102, 
    0.003049792, 0.003052857, 0.00305987, 0.003056076, 0.003060507, 
    0.003050714, 0.003045623, 0.0030443, 0.003041842, 0.00304435, 
    0.003044146, 0.003046547, 0.003045769, 0.003051537, 0.003048438, 
    0.003057228, 0.003060435, 0.003069467, 0.003074991, 0.003080607, 
    0.00308308, 0.003083832, 0.003084144,
  0.00181005, 0.001816801, 0.001815489, 0.00182093, 0.001817912, 0.001821475, 
    0.001811419, 0.001817069, 0.001813462, 0.001810657, 0.001831478, 
    0.001821173, 0.001842159, 0.001835602, 0.00185206, 0.00184114, 
    0.001854259, 0.001851744, 0.001859308, 0.001857142, 0.001866807, 
    0.001860307, 0.00187181, 0.001865255, 0.001866281, 0.001860093, 
    0.001823247, 0.001830196, 0.001822835, 0.001823827, 0.001823382, 
    0.001817975, 0.001815249, 0.001809533, 0.001810571, 0.001814768, 
    0.001824273, 0.001821047, 0.001829171, 0.001828987, 0.001838019, 
    0.001833948, 0.001849107, 0.001844802, 0.001857232, 0.001854109, 
    0.001857086, 0.001856183, 0.001857097, 0.001852516, 0.001854479, 
    0.001850446, 0.001834711, 0.00183934, 0.001825524, 0.001817203, 
    0.001811667, 0.001807736, 0.001808292, 0.001809352, 0.001814793, 
    0.001819904, 0.001823796, 0.001826398, 0.001828961, 0.001836714, 
    0.001840812, 0.001849978, 0.001848324, 0.001851125, 0.001853798, 
    0.001858285, 0.001857546, 0.001859522, 0.00185105, 0.001856683, 
    0.001847382, 0.001849927, 0.001829661, 0.001821917, 0.001818626, 
    0.001815741, 0.001808719, 0.00181357, 0.001811658, 0.001816204, 
    0.001819091, 0.001817663, 0.001826469, 0.001823047, 0.001841055, 
    0.001833305, 0.001853486, 0.001848663, 0.001854642, 0.001851592, 
    0.001856817, 0.001852114, 0.001860257, 0.00186203, 0.001860819, 
    0.001865467, 0.001851854, 0.001857086, 0.001817623, 0.001817856, 
    0.001818941, 0.001814172, 0.001813879, 0.001809504, 0.001813397, 
    0.001815054, 0.001819258, 0.001821744, 0.001824105, 0.001829295, 
    0.001835086, 0.001843173, 0.001848976, 0.001852863, 0.001850479, 
    0.001852583, 0.001850231, 0.001849129, 0.001861366, 0.001854498, 
    0.001864799, 0.001864229, 0.00185957, 0.001864293, 0.00181802, 
    0.001816679, 0.001812024, 0.001815667, 0.001809028, 0.001812746, 
    0.001814883, 0.00182312, 0.001824927, 0.001826603, 0.001829912, 
    0.001834157, 0.001841595, 0.001848059, 0.001853953, 0.001853522, 
    0.001853674, 0.00185499, 0.001851729, 0.001855525, 0.001856162, 
    0.001854497, 0.001864153, 0.001861396, 0.001864217, 0.001862422, 
    0.001817115, 0.00181937, 0.001818151, 0.001820442, 0.001818829, 
    0.001826002, 0.00182815, 0.001838194, 0.001834073, 0.00184063, 
    0.001834739, 0.001835784, 0.001840845, 0.001835058, 0.001847704, 
    0.001839134, 0.001855041, 0.001846496, 0.001855576, 0.001853928, 
    0.001856657, 0.001859099, 0.001862171, 0.001867835, 0.001866524, 
    0.001871256, 0.001822729, 0.001825652, 0.001825394, 0.00182845, 
    0.001830709, 0.001835603, 0.001843443, 0.001840496, 0.001845905, 
    0.001846991, 0.001838772, 0.00184382, 0.001827606, 0.001830229, 
    0.001828667, 0.00182296, 0.001841176, 0.001831835, 0.001849072, 
    0.00184402, 0.001858751, 0.001851431, 0.001865802, 0.001871936, 
    0.0018777, 0.001884432, 0.001827245, 0.00182526, 0.001828813, 
    0.001833726, 0.00183828, 0.001844328, 0.001844947, 0.001846079, 
    0.001849011, 0.001851475, 0.001846438, 0.001852093, 0.001830839, 
    0.001841986, 0.00182451, 0.001829779, 0.001833437, 0.001831832, 
    0.001840159, 0.00184212, 0.001850083, 0.001845968, 0.001870423, 
    0.001859616, 0.00188955, 0.001881202, 0.001824567, 0.001827238, 
    0.001836526, 0.001832109, 0.001844732, 0.001847835, 0.001850356, 
    0.001853578, 0.001853925, 0.001855833, 0.001852706, 0.00185571, 
    0.001844341, 0.001849424, 0.001835464, 0.001838866, 0.001837301, 
    0.001835585, 0.00184088, 0.001846517, 0.001846637, 0.001848443, 
    0.001853533, 0.001844783, 0.001871819, 0.001855139, 0.001830149, 
    0.00183529, 0.001836023, 0.001834032, 0.001847524, 0.001842639, 
    0.001855787, 0.001852236, 0.001858052, 0.001855163, 0.001854738, 
    0.001851024, 0.001848711, 0.001842863, 0.001838101, 0.001834321, 
    0.0018352, 0.001839351, 0.001846862, 0.001853957, 0.001852404, 
    0.00185761, 0.001843817, 0.001849606, 0.001847369, 0.001853198, 
    0.001840418, 0.001851306, 0.001837632, 0.001838832, 0.001842542, 
    0.001849999, 0.001851645, 0.001853405, 0.001852319, 0.001847052, 
    0.001846188, 0.001842452, 0.00184142, 0.001838571, 0.001836211, 
    0.001838367, 0.001840631, 0.001847054, 0.001852837, 0.001859135, 
    0.001860674, 0.001868025, 0.001862043, 0.001871912, 0.001863525, 
    0.001878034, 0.001851935, 0.001863276, 0.001842711, 0.001844929, 
    0.001848942, 0.001858131, 0.001853171, 0.001858971, 0.001846154, 
    0.001839495, 0.00183777, 0.001834551, 0.001837843, 0.001837575, 
    0.001840724, 0.001839712, 0.001847267, 0.00184321, 0.001854727, 
    0.001858925, 0.001870761, 0.001878005, 0.001885367, 0.001888615, 
    0.001889603, 0.001890016,
  0.001646086, 0.00165329, 0.001651889, 0.001657697, 0.001654476, 
    0.001658278, 0.001647546, 0.001653576, 0.001649727, 0.001646734, 
    0.001668958, 0.001657956, 0.001680369, 0.001673364, 0.001690951, 
    0.00167928, 0.001693302, 0.001690614, 0.001698701, 0.001696385, 
    0.001706722, 0.00169977, 0.001712075, 0.001705062, 0.00170616, 
    0.001699541, 0.001660171, 0.00166759, 0.001659731, 0.001660789, 
    0.001660314, 0.001654543, 0.001651633, 0.001645534, 0.001646642, 
    0.00165112, 0.001661265, 0.001657822, 0.001666495, 0.001666299, 
    0.001675946, 0.001671598, 0.001687795, 0.001683194, 0.001696482, 
    0.001693142, 0.001696325, 0.00169536, 0.001696337, 0.001691439, 
    0.001693538, 0.001689226, 0.001672412, 0.001677357, 0.001662601, 
    0.001653718, 0.001647811, 0.001643618, 0.001644211, 0.001645341, 
    0.001651147, 0.001656601, 0.001660756, 0.001663535, 0.001666271, 
    0.001674552, 0.00167893, 0.001688725, 0.001686958, 0.001689952, 
    0.00169281, 0.001697607, 0.001696818, 0.001698931, 0.001689872, 
    0.001695894, 0.001685951, 0.001688672, 0.001667018, 0.001658751, 
    0.001655237, 0.001652159, 0.001644666, 0.001649841, 0.001647802, 
    0.001652653, 0.001655734, 0.00165421, 0.001663611, 0.001659957, 
    0.001679189, 0.00167091, 0.001692476, 0.00168732, 0.001693712, 
    0.001690451, 0.001696037, 0.00169101, 0.001699717, 0.001701612, 
    0.001700317, 0.001705289, 0.001690731, 0.001696325, 0.001654167, 
    0.001654416, 0.001655574, 0.001650484, 0.001650172, 0.001645504, 
    0.001649657, 0.001651426, 0.001655912, 0.001658566, 0.001661087, 
    0.001666628, 0.001672813, 0.001681453, 0.001687655, 0.00169181, 
    0.001689262, 0.001691511, 0.001688997, 0.001687818, 0.001700902, 
    0.001693558, 0.001704574, 0.001703965, 0.001698981, 0.001704034, 
    0.001654591, 0.00165316, 0.001648193, 0.00165208, 0.001644996, 
    0.001648962, 0.001651242, 0.001660034, 0.001661964, 0.001663754, 
    0.001667287, 0.00167182, 0.001679767, 0.001686675, 0.001692976, 
    0.001692514, 0.001692677, 0.001694084, 0.001690598, 0.001694656, 
    0.001695337, 0.001693557, 0.001703883, 0.001700934, 0.001703952, 
    0.001702032, 0.001653625, 0.001656032, 0.001654731, 0.001657177, 
    0.001655454, 0.001663111, 0.001665405, 0.001676133, 0.001671731, 
    0.001678735, 0.001672443, 0.001673558, 0.001678964, 0.001672783, 
    0.001686295, 0.001677137, 0.001694139, 0.001685003, 0.001694711, 
    0.001692949, 0.001695866, 0.001698478, 0.001701763, 0.001707822, 
    0.001706419, 0.001711483, 0.001659618, 0.001662738, 0.001662462, 
    0.001665726, 0.001668138, 0.001673365, 0.001681742, 0.001678593, 
    0.001684373, 0.001685533, 0.001676751, 0.001682144, 0.001664824, 
    0.001667625, 0.001665957, 0.001659864, 0.001679319, 0.00166934, 
    0.001687757, 0.001682358, 0.001698106, 0.001690278, 0.001705647, 
    0.00171221, 0.001718379, 0.001725586, 0.001664439, 0.00166232, 
    0.001666114, 0.00167136, 0.001676224, 0.001682688, 0.001683348, 
    0.001684559, 0.001687692, 0.001690327, 0.001684942, 0.001690987, 
    0.001668276, 0.001680185, 0.001661519, 0.001667144, 0.001671051, 
    0.001669337, 0.001678232, 0.001680328, 0.001688838, 0.001684439, 
    0.001710591, 0.001699031, 0.001731067, 0.001722127, 0.00166158, 
    0.001664432, 0.001674351, 0.001669633, 0.001683119, 0.001686435, 
    0.00168913, 0.001692574, 0.001692946, 0.001694986, 0.001691643, 
    0.001694854, 0.001682701, 0.001688134, 0.001673217, 0.00167685, 
    0.001675179, 0.001673346, 0.001679003, 0.001685027, 0.001685155, 
    0.001687085, 0.001692525, 0.001683173, 0.001712083, 0.001694242, 
    0.001667541, 0.001673031, 0.001673813, 0.001671688, 0.001686103, 
    0.001680883, 0.001694936, 0.00169114, 0.001697359, 0.001694269, 
    0.001693814, 0.001689844, 0.001687372, 0.001681122, 0.001676033, 
    0.001671996, 0.001672935, 0.001677369, 0.001685395, 0.00169298, 
    0.001691319, 0.001696886, 0.001682142, 0.001688328, 0.001685938, 
    0.001692168, 0.001678509, 0.001690144, 0.001675533, 0.001676815, 
    0.001680779, 0.001688748, 0.001690508, 0.00169239, 0.001691229, 
    0.001685598, 0.001684675, 0.001680682, 0.00167958, 0.001676536, 
    0.001674015, 0.001676318, 0.001678737, 0.0016856, 0.001691782, 
    0.001698516, 0.001700163, 0.001708024, 0.001701626, 0.001712183, 
    0.00170321, 0.001718735, 0.001690817, 0.001702945, 0.001680959, 
    0.00168333, 0.001687618, 0.001697442, 0.001692139, 0.001698341, 
    0.001684639, 0.001677523, 0.00167568, 0.001672241, 0.001675758, 
    0.001675472, 0.001678836, 0.001677755, 0.001685828, 0.001681493, 
    0.001693803, 0.001698291, 0.001710953, 0.001718705, 0.001726588, 
    0.001730066, 0.001731125, 0.001731567,
  0.001514891, 0.001522022, 0.001520635, 0.001526386, 0.001523196, 
    0.001526962, 0.001516336, 0.001522305, 0.001518495, 0.001515532, 
    0.001537543, 0.001526643, 0.001548858, 0.001541911, 0.001559359, 
    0.001547778, 0.001561694, 0.001559024, 0.001567055, 0.001564755, 
    0.001575025, 0.001568117, 0.001580346, 0.001573375, 0.001574466, 
    0.001567889, 0.001528836, 0.001536187, 0.001528401, 0.001529449, 
    0.001528978, 0.001523262, 0.001520381, 0.001514345, 0.001515441, 
    0.001519874, 0.00152992, 0.00152651, 0.001535102, 0.001534908, 
    0.001544471, 0.00154016, 0.001556227, 0.001551661, 0.001564851, 
    0.001561535, 0.001564695, 0.001563737, 0.001564708, 0.001559844, 
    0.001561928, 0.001557647, 0.001540968, 0.001545871, 0.001531244, 
    0.001522446, 0.001516598, 0.001512449, 0.001513035, 0.001514154, 
    0.0015199, 0.001525301, 0.001529416, 0.001532169, 0.00153488, 
    0.001543089, 0.00154743, 0.00155715, 0.001555396, 0.001558367, 
    0.001561205, 0.001565969, 0.001565184, 0.001567283, 0.001558288, 
    0.001564267, 0.001554396, 0.001557096, 0.00153562, 0.00152743, 
    0.00152395, 0.001520902, 0.001513486, 0.001518608, 0.001516589, 
    0.001521391, 0.001524442, 0.001522933, 0.001532244, 0.001528625, 
    0.001547688, 0.001539478, 0.001560874, 0.001555756, 0.0015621, 
    0.001558863, 0.00156441, 0.001559418, 0.001568064, 0.001569947, 
    0.00156866, 0.001573601, 0.001559141, 0.001564695, 0.001522891, 
    0.001523137, 0.001524283, 0.001519244, 0.001518935, 0.001514315, 
    0.001518426, 0.001520176, 0.001524619, 0.001527246, 0.001529744, 
    0.001535234, 0.001541364, 0.001549933, 0.001556087, 0.001560212, 
    0.001557683, 0.001559915, 0.00155742, 0.001556249, 0.001569242, 
    0.001561947, 0.00157289, 0.001572285, 0.001567333, 0.001572353, 
    0.00152331, 0.001521893, 0.001516976, 0.001520824, 0.001513812, 
    0.001517738, 0.001519995, 0.001528701, 0.001530613, 0.001532386, 
    0.001535887, 0.001540381, 0.001548261, 0.001555115, 0.00156137, 
    0.001560911, 0.001561073, 0.00156247, 0.001559009, 0.001563038, 
    0.001563714, 0.001561946, 0.001572204, 0.001569274, 0.001572272, 
    0.001570364, 0.001522354, 0.001524737, 0.001523449, 0.001525871, 
    0.001524165, 0.001531749, 0.001534022, 0.001544657, 0.001540292, 
    0.001547237, 0.001540998, 0.001542104, 0.001547465, 0.001541335, 
    0.001554738, 0.001545653, 0.001562524, 0.001553456, 0.001563092, 
    0.001561343, 0.00156424, 0.001566834, 0.001570097, 0.001576118, 
    0.001574724, 0.001579757, 0.001528289, 0.001531379, 0.001531107, 
    0.00153434, 0.001536731, 0.001541912, 0.00155022, 0.001547096, 
    0.00155283, 0.001553982, 0.001545269, 0.001550619, 0.001533447, 
    0.001536223, 0.00153457, 0.001528533, 0.001547817, 0.001537922, 
    0.001556189, 0.001550831, 0.001566464, 0.001558692, 0.001573956, 
    0.00158048, 0.001586616, 0.001593787, 0.001533065, 0.001530965, 
    0.001534724, 0.001539925, 0.001544748, 0.001551158, 0.001551814, 
    0.001553015, 0.001556125, 0.001558739, 0.001553395, 0.001559395, 
    0.001536867, 0.001548675, 0.001530172, 0.001535746, 0.001539618, 
    0.001537919, 0.001546739, 0.001548817, 0.001557262, 0.001552897, 
    0.001578871, 0.001567383, 0.001599243, 0.001590345, 0.001530232, 
    0.001533058, 0.00154289, 0.001538212, 0.001551586, 0.001554877, 
    0.001557552, 0.001560971, 0.00156134, 0.001563365, 0.001560046, 
    0.001563234, 0.001551172, 0.001556563, 0.001541766, 0.001545368, 
    0.001543711, 0.001541893, 0.001547503, 0.001553479, 0.001553606, 
    0.001555522, 0.001560922, 0.00155164, 0.001580354, 0.001562627, 
    0.001536138, 0.00154158, 0.001542357, 0.001540249, 0.001554547, 
    0.001549368, 0.001563316, 0.001559547, 0.001565722, 0.001562654, 
    0.001562202, 0.001558261, 0.001555807, 0.001549605, 0.001544558, 
    0.001540555, 0.001541486, 0.001545883, 0.001553845, 0.001561373, 
    0.001559725, 0.001565253, 0.001550617, 0.001556755, 0.001554383, 
    0.001560568, 0.001547013, 0.001558559, 0.001544062, 0.001545333, 
    0.001549265, 0.001557172, 0.00155892, 0.001560788, 0.001559635, 
    0.001554047, 0.001553131, 0.001549169, 0.001548075, 0.001545056, 
    0.001542556, 0.00154484, 0.001547239, 0.001554049, 0.001560184, 
    0.001566871, 0.001568507, 0.001576319, 0.001569961, 0.001580453, 
    0.001571535, 0.00158697, 0.001559226, 0.001571271, 0.001549443, 
    0.001551796, 0.001556051, 0.001565805, 0.001560539, 0.001566697, 
    0.001553095, 0.001546035, 0.001544207, 0.001540798, 0.001544285, 
    0.001544002, 0.001547338, 0.001546266, 0.001554275, 0.001549973, 
    0.001562191, 0.001566648, 0.00157923, 0.00158694, 0.001594784, 
    0.001598247, 0.001599301, 0.001599741,
  0.0013795, 0.001385892, 0.001384649, 0.001389807, 0.001386945, 0.001390323, 
    0.001380795, 0.001386146, 0.00138273, 0.001380075, 0.001399825, 
    0.001390037, 0.001409999, 0.00140375, 0.001419454, 0.001409026, 
    0.001421557, 0.001419152, 0.001426391, 0.001424317, 0.001433584, 
    0.001427349, 0.00143839, 0.001432094, 0.001433079, 0.001427144, 
    0.001392005, 0.001398606, 0.001391615, 0.001392556, 0.001392133, 
    0.001387005, 0.001384421, 0.001379011, 0.001379993, 0.001383967, 
    0.001392979, 0.001389918, 0.001397632, 0.001397457, 0.001406052, 
    0.001402176, 0.001416632, 0.001412521, 0.001424404, 0.001421414, 
    0.001424263, 0.001423399, 0.001424274, 0.00141989, 0.001421768, 
    0.001417911, 0.001402902, 0.001407311, 0.001394167, 0.001386272, 
    0.00138103, 0.001377312, 0.001377838, 0.00137884, 0.00138399, 
    0.001388833, 0.001392526, 0.001394997, 0.001397432, 0.001404809, 
    0.001408714, 0.001417463, 0.001415883, 0.00141856, 0.001421117, 
    0.001425412, 0.001424704, 0.001426597, 0.001418489, 0.001423877, 
    0.001414983, 0.001417415, 0.001398097, 0.001390744, 0.001387622, 
    0.001384888, 0.001378242, 0.001382831, 0.001381022, 0.001385326, 
    0.001388063, 0.001386709, 0.001395065, 0.001391816, 0.001408945, 
    0.001401563, 0.001420818, 0.001416207, 0.001421924, 0.001419006, 
    0.001424006, 0.001419506, 0.001427302, 0.001429, 0.001427839, 
    0.001432298, 0.001419257, 0.001424263, 0.001386671, 0.001386892, 
    0.00138792, 0.001383401, 0.001383125, 0.001378984, 0.001382668, 
    0.001384237, 0.001388221, 0.001390579, 0.00139282, 0.00139775, 
    0.001403259, 0.001410966, 0.001416506, 0.001420222, 0.001417943, 
    0.001419955, 0.001417706, 0.001416652, 0.001428364, 0.001421786, 
    0.001431657, 0.00143111, 0.001426642, 0.001431172, 0.001387047, 
    0.001385777, 0.001381369, 0.001384818, 0.001378534, 0.001382051, 
    0.001384075, 0.001391884, 0.0013936, 0.001395192, 0.001398337, 
    0.001402374, 0.001409461, 0.00141563, 0.001421265, 0.001420852, 
    0.001420998, 0.001422257, 0.001419138, 0.001422769, 0.001423379, 
    0.001421785, 0.001431037, 0.001428393, 0.001431098, 0.001429377, 
    0.00138619, 0.001388327, 0.001387172, 0.001389344, 0.001387814, 
    0.00139462, 0.001396662, 0.001406219, 0.001402295, 0.00140854, 
    0.001402929, 0.001403923, 0.001408745, 0.001403232, 0.001415291, 
    0.001407115, 0.001422306, 0.001414137, 0.001422818, 0.001421241, 
    0.001423852, 0.001426192, 0.001429136, 0.001434571, 0.001433312, 
    0.001437858, 0.001391514, 0.001394288, 0.001394043, 0.001396947, 
    0.001399095, 0.001403751, 0.001411224, 0.001408413, 0.001413573, 
    0.00141461, 0.00140677, 0.001411583, 0.001396145, 0.001398638, 
    0.001397153, 0.001391733, 0.001409061, 0.001400165, 0.001416598, 
    0.001411774, 0.001425858, 0.001418852, 0.001432619, 0.001438511, 
    0.001444058, 0.001450546, 0.001395802, 0.001393917, 0.001397292, 
    0.001401965, 0.0014063, 0.001412068, 0.001412658, 0.00141374, 0.00141654, 
    0.001418895, 0.001414082, 0.001419486, 0.001399217, 0.001409834, 
    0.001393205, 0.00139821, 0.001401689, 0.001400162, 0.001408092, 
    0.001409962, 0.001417564, 0.001413633, 0.001437057, 0.001426687, 
    0.001455488, 0.001447431, 0.001393258, 0.001395795, 0.00140463, 
    0.001400425, 0.001412453, 0.001415416, 0.001417825, 0.001420906, 
    0.001421238, 0.001423064, 0.001420072, 0.001422946, 0.001412081, 
    0.001416935, 0.001403619, 0.001406859, 0.001405368, 0.001403734, 
    0.001408779, 0.001414158, 0.001414272, 0.001415997, 0.001420862, 
    0.001412502, 0.001438398, 0.001422399, 0.001398562, 0.001403453, 
    0.001404151, 0.001402256, 0.001415119, 0.001410457, 0.00142302, 
    0.001419623, 0.001425189, 0.001422423, 0.001422016, 0.001418464, 
    0.001416253, 0.00141067, 0.00140613, 0.001402531, 0.001403367, 
    0.001407322, 0.001414487, 0.001421269, 0.001419783, 0.001424766, 
    0.001411581, 0.001417108, 0.001414971, 0.001420543, 0.001408338, 
    0.001418732, 0.001405684, 0.001406827, 0.001410364, 0.001417483, 
    0.001419058, 0.001420741, 0.001419702, 0.001414668, 0.001413844, 
    0.001410278, 0.001409294, 0.001406578, 0.00140433, 0.001406384, 
    0.001408542, 0.00141467, 0.001420197, 0.001426225, 0.001427701, 
    0.001434752, 0.001429013, 0.001438487, 0.001430433, 0.001444378, 
    0.001419334, 0.001430195, 0.001410525, 0.001412642, 0.001416473, 
    0.001425264, 0.001420516, 0.001426069, 0.001413811, 0.001407459, 
    0.001405815, 0.00140275, 0.001405885, 0.00140563, 0.00140863, 
    0.001407666, 0.001414874, 0.001411001, 0.001422006, 0.001426024, 
    0.001437382, 0.001444351, 0.001451449, 0.001454585, 0.001455539, 
    0.001455938,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.34871e-06, 1.360258e-06, 1.358009e-06, 1.367352e-06, 1.362165e-06, 
    1.368289e-06, 1.351046e-06, 1.360717e-06, 1.354539e-06, 1.349746e-06, 
    1.385578e-06, 1.367769e-06, 1.404196e-06, 1.392747e-06, 1.421594e-06, 
    1.402411e-06, 1.425478e-06, 1.421037e-06, 1.434419e-06, 1.430579e-06, 
    1.447767e-06, 1.436193e-06, 1.456716e-06, 1.444998e-06, 1.446828e-06, 
    1.435812e-06, 1.371343e-06, 1.383356e-06, 1.370633e-06, 1.372342e-06, 
    1.371575e-06, 1.362272e-06, 1.357596e-06, 1.347827e-06, 1.349598e-06, 
    1.356773e-06, 1.37311e-06, 1.367552e-06, 1.381578e-06, 1.381261e-06, 
    1.39696e-06, 1.38987e-06, 1.416391e-06, 1.408827e-06, 1.430739e-06, 
    1.425212e-06, 1.430479e-06, 1.42888e-06, 1.430499e-06, 1.422398e-06, 
    1.425866e-06, 1.418748e-06, 1.391199e-06, 1.399268e-06, 1.375271e-06, 
    1.360945e-06, 1.351469e-06, 1.344766e-06, 1.345712e-06, 1.347518e-06, 
    1.356815e-06, 1.365585e-06, 1.372288e-06, 1.376781e-06, 1.381215e-06, 
    1.394684e-06, 1.401837e-06, 1.417923e-06, 1.415012e-06, 1.419944e-06, 
    1.424663e-06, 1.432604e-06, 1.431295e-06, 1.434799e-06, 1.419812e-06, 
    1.429764e-06, 1.413354e-06, 1.417833e-06, 1.382427e-06, 1.369051e-06, 
    1.363389e-06, 1.35844e-06, 1.34644e-06, 1.354721e-06, 1.351454e-06, 
    1.359233e-06, 1.364188e-06, 1.361735e-06, 1.376903e-06, 1.370996e-06, 
    1.402262e-06, 1.388751e-06, 1.424112e-06, 1.415609e-06, 1.426153e-06, 
    1.420767e-06, 1.430002e-06, 1.421689e-06, 1.436104e-06, 1.439253e-06, 
    1.4371e-06, 1.445375e-06, 1.421228e-06, 1.430478e-06, 1.361668e-06, 
    1.362068e-06, 1.36393e-06, 1.355751e-06, 1.355251e-06, 1.347778e-06, 
    1.354426e-06, 1.357263e-06, 1.364475e-06, 1.36875e-06, 1.372821e-06, 
    1.381793e-06, 1.391848e-06, 1.40597e-06, 1.416159e-06, 1.42301e-06, 
    1.418807e-06, 1.422517e-06, 1.418369e-06, 1.416427e-06, 1.438072e-06, 
    1.425898e-06, 1.444183e-06, 1.443168e-06, 1.434881e-06, 1.443282e-06, 
    1.362348e-06, 1.360048e-06, 1.352079e-06, 1.358313e-06, 1.346965e-06, 
    1.353312e-06, 1.356968e-06, 1.37112e-06, 1.374239e-06, 1.377135e-06, 
    1.382863e-06, 1.390232e-06, 1.403207e-06, 1.414546e-06, 1.424936e-06, 
    1.424174e-06, 1.424442e-06, 1.426768e-06, 1.421009e-06, 1.427715e-06, 
    1.428842e-06, 1.425896e-06, 1.443032e-06, 1.438126e-06, 1.443146e-06, 
    1.43995e-06, 1.360795e-06, 1.364667e-06, 1.362574e-06, 1.366511e-06, 
    1.363736e-06, 1.376094e-06, 1.37981e-06, 1.397265e-06, 1.390087e-06, 
    1.401518e-06, 1.391245e-06, 1.393063e-06, 1.401893e-06, 1.391798e-06, 
    1.41392e-06, 1.398904e-06, 1.426859e-06, 1.411796e-06, 1.427805e-06, 
    1.42489e-06, 1.429717e-06, 1.434047e-06, 1.439503e-06, 1.4496e-06, 
    1.447258e-06, 1.455722e-06, 1.370449e-06, 1.37549e-06, 1.375045e-06, 
    1.380329e-06, 1.384244e-06, 1.392748e-06, 1.406443e-06, 1.401285e-06, 
    1.410761e-06, 1.412667e-06, 1.398273e-06, 1.407103e-06, 1.378867e-06, 
    1.38341e-06, 1.380704e-06, 1.370844e-06, 1.402473e-06, 1.386195e-06, 
    1.416326e-06, 1.407452e-06, 1.433429e-06, 1.420481e-06, 1.44597e-06, 
    1.456939e-06, 1.467297e-06, 1.479453e-06, 1.378245e-06, 1.374814e-06, 
    1.380958e-06, 1.389483e-06, 1.397414e-06, 1.407994e-06, 1.409079e-06, 
    1.411066e-06, 1.41622e-06, 1.420562e-06, 1.411695e-06, 1.421651e-06, 
    1.384466e-06, 1.40389e-06, 1.373517e-06, 1.382629e-06, 1.388977e-06, 
    1.38619e-06, 1.400694e-06, 1.404124e-06, 1.418105e-06, 1.410868e-06, 
    1.454228e-06, 1.434963e-06, 1.488739e-06, 1.473611e-06, 1.373617e-06, 
    1.378232e-06, 1.394356e-06, 1.386672e-06, 1.408701e-06, 1.414151e-06, 
    1.418588e-06, 1.424273e-06, 1.424886e-06, 1.42826e-06, 1.422733e-06, 
    1.428041e-06, 1.408015e-06, 1.416946e-06, 1.392505e-06, 1.398435e-06, 
    1.395705e-06, 1.392714e-06, 1.401954e-06, 1.411833e-06, 1.412043e-06, 
    1.415219e-06, 1.424189e-06, 1.408788e-06, 1.456726e-06, 1.427027e-06, 
    1.383273e-06, 1.392202e-06, 1.393479e-06, 1.390015e-06, 1.413604e-06, 
    1.405034e-06, 1.428177e-06, 1.421903e-06, 1.43219e-06, 1.427074e-06, 
    1.426321e-06, 1.419765e-06, 1.415691e-06, 1.405425e-06, 1.397099e-06, 
    1.390515e-06, 1.392044e-06, 1.399282e-06, 1.412438e-06, 1.42494e-06, 
    1.422197e-06, 1.431405e-06, 1.407095e-06, 1.417264e-06, 1.413329e-06, 
    1.423599e-06, 1.401148e-06, 1.420261e-06, 1.396283e-06, 1.398377e-06, 
    1.404863e-06, 1.417958e-06, 1.420861e-06, 1.423967e-06, 1.422049e-06, 
    1.412774e-06, 1.411256e-06, 1.404704e-06, 1.402898e-06, 1.39792e-06, 
    1.393804e-06, 1.397564e-06, 1.401518e-06, 1.412776e-06, 1.422961e-06, 
    1.434107e-06, 1.436841e-06, 1.449936e-06, 1.439273e-06, 1.456892e-06, 
    1.441908e-06, 1.467894e-06, 1.42137e-06, 1.441469e-06, 1.405158e-06, 
    1.409047e-06, 1.416096e-06, 1.432329e-06, 1.423552e-06, 1.433818e-06, 
    1.411197e-06, 1.399533e-06, 1.396522e-06, 1.390915e-06, 1.39665e-06, 
    1.396183e-06, 1.401681e-06, 1.399912e-06, 1.41315e-06, 1.406031e-06, 
    1.426301e-06, 1.433735e-06, 1.454832e-06, 1.467844e-06, 1.481147e-06, 
    1.48704e-06, 1.488835e-06, 1.489586e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.296261e-06, 8.332859e-06, 8.325721e-06, 8.355265e-06, 8.33886e-06, 
    8.358198e-06, 8.303632e-06, 8.334261e-06, 8.314692e-06, 8.299478e-06, 
    8.4126e-06, 8.356517e-06, 8.470882e-06, 8.435052e-06, 8.525057e-06, 
    8.46529e-06, 8.537108e-06, 8.5233e-06, 8.564803e-06, 8.552895e-06, 
    8.606034e-06, 8.570272e-06, 8.633576e-06, 8.597471e-06, 8.60311e-06, 
    8.569054e-06, 8.367845e-06, 8.405676e-06, 8.365591e-06, 8.370985e-06, 
    8.368553e-06, 8.339168e-06, 8.324378e-06, 8.293383e-06, 8.298994e-06, 
    8.321747e-06, 8.37335e-06, 8.355804e-06, 8.399978e-06, 8.398982e-06, 
    8.448213e-06, 8.426003e-06, 8.508841e-06, 8.485264e-06, 8.553382e-06, 
    8.536229e-06, 8.552563e-06, 8.547594e-06, 8.552604e-06, 8.52747e-06, 
    8.53822e-06, 8.516106e-06, 8.43026e-06, 8.455516e-06, 8.380198e-06, 
    8.334977e-06, 8.304943e-06, 8.28366e-06, 8.286651e-06, 8.292391e-06, 
    8.321865e-06, 8.349586e-06, 8.370732e-06, 8.384874e-06, 8.398814e-06, 
    8.441095e-06, 8.463457e-06, 8.513594e-06, 8.504528e-06, 8.519864e-06, 
    8.534515e-06, 8.559129e-06, 8.55507e-06, 8.565912e-06, 8.519409e-06, 
    8.550307e-06, 8.499297e-06, 8.513241e-06, 8.402722e-06, 8.360568e-06, 
    8.342694e-06, 8.327021e-06, 8.288959e-06, 8.315236e-06, 8.304866e-06, 
    8.329496e-06, 8.345163e-06, 8.337398e-06, 8.385253e-06, 8.366629e-06, 
    8.464771e-06, 8.422468e-06, 8.532816e-06, 8.506368e-06, 8.539129e-06, 
    8.522405e-06, 8.551053e-06, 8.525254e-06, 8.569933e-06, 8.579677e-06, 
    8.573002e-06, 8.59857e-06, 8.523774e-06, 8.552483e-06, 8.337231e-06, 
    8.338497e-06, 8.344374e-06, 8.318487e-06, 8.3169e-06, 8.293182e-06, 
    8.31426e-06, 8.323249e-06, 8.346048e-06, 8.359539e-06, 8.372366e-06, 
    8.40061e-06, 8.432165e-06, 8.476322e-06, 8.508073e-06, 8.52936e-06, 
    8.516293e-06, 8.527813e-06, 8.514918e-06, 8.508862e-06, 8.576005e-06, 
    8.53829e-06, 8.594868e-06, 8.591735e-06, 8.566107e-06, 8.592065e-06, 
    8.339368e-06, 8.33208e-06, 8.306838e-06, 8.326576e-06, 8.290584e-06, 
    8.310727e-06, 8.322303e-06, 8.367014e-06, 8.376827e-06, 8.385951e-06, 
    8.403956e-06, 8.427077e-06, 8.467687e-06, 8.503036e-06, 8.535333e-06, 
    8.532952e-06, 8.533782e-06, 8.540992e-06, 8.523106e-06, 8.543911e-06, 
    8.547398e-06, 8.53826e-06, 8.591292e-06, 8.576131e-06, 8.591635e-06, 
    8.581749e-06, 8.334435e-06, 8.346664e-06, 8.340038e-06, 8.352481e-06, 
    8.343701e-06, 8.38269e-06, 8.394375e-06, 8.449124e-06, 8.426623e-06, 
    8.462415e-06, 8.430238e-06, 8.435939e-06, 8.463569e-06, 8.431952e-06, 
    8.501067e-06, 8.454194e-06, 8.541264e-06, 8.494429e-06, 8.544183e-06, 
    8.535126e-06, 8.550088e-06, 8.563507e-06, 8.580368e-06, 8.61154e-06, 
    8.6043e-06, 8.630375e-06, 8.364907e-06, 8.380787e-06, 8.379378e-06, 
    8.395999e-06, 8.408296e-06, 8.434976e-06, 8.477795e-06, 8.461669e-06, 
    8.491236e-06, 8.49718e-06, 8.452224e-06, 8.479818e-06, 8.391338e-06, 
    8.405614e-06, 8.397098e-06, 8.366039e-06, 8.465322e-06, 8.414331e-06, 
    8.508501e-06, 8.480837e-06, 8.561571e-06, 8.521405e-06, 8.600321e-06, 
    8.634122e-06, 8.665914e-06, 8.703124e-06, 8.389448e-06, 8.378634e-06, 
    8.397959e-06, 8.424739e-06, 8.449563e-06, 8.482623e-06, 8.485993e-06, 
    8.492178e-06, 8.508217e-06, 8.521723e-06, 8.494124e-06, 8.525084e-06, 
    8.408931e-06, 8.469745e-06, 8.37445e-06, 8.403131e-06, 8.423043e-06, 
    8.414295e-06, 8.45972e-06, 8.470425e-06, 8.513995e-06, 8.49146e-06, 
    8.62576e-06, 8.56629e-06, 8.731447e-06, 8.68524e-06, 8.374854e-06, 
    8.389374e-06, 8.439988e-06, 8.415895e-06, 8.484804e-06, 8.501791e-06, 
    8.51558e-06, 8.533248e-06, 8.535133e-06, 8.545605e-06, 8.528432e-06, 
    8.544908e-06, 8.482605e-06, 8.510429e-06, 8.434102e-06, 8.452655e-06, 
    8.444107e-06, 8.434728e-06, 8.463631e-06, 8.494468e-06, 8.495106e-06, 
    8.504987e-06, 8.532891e-06, 8.484932e-06, 8.633428e-06, 8.541667e-06, 
    8.405217e-06, 8.433234e-06, 8.437216e-06, 8.426359e-06, 8.500065e-06, 
    8.473341e-06, 8.545348e-06, 8.525858e-06, 8.557761e-06, 8.541902e-06, 
    8.539552e-06, 8.51919e-06, 8.5065e-06, 8.474503e-06, 8.448464e-06, 
    8.427836e-06, 8.432613e-06, 8.455278e-06, 8.496329e-06, 8.535209e-06, 
    8.526679e-06, 8.555232e-06, 8.479635e-06, 8.511322e-06, 8.499058e-06, 
    8.530995e-06, 8.461209e-06, 8.520806e-06, 8.445983e-06, 8.452524e-06, 
    8.472787e-06, 8.513603e-06, 8.522604e-06, 8.532256e-06, 8.526281e-06, 
    8.497431e-06, 8.492691e-06, 8.472238e-06, 8.46659e-06, 8.451023e-06, 
    8.438124e-06, 8.449897e-06, 8.462246e-06, 8.497374e-06, 8.529046e-06, 
    8.563598e-06, 8.572053e-06, 8.61249e-06, 8.57957e-06, 8.633901e-06, 
    8.587711e-06, 8.667665e-06, 8.524223e-06, 8.586503e-06, 8.473708e-06, 
    8.48583e-06, 8.507794e-06, 8.558183e-06, 8.530945e-06, 8.562785e-06, 
    8.492499e-06, 8.456079e-06, 8.446641e-06, 8.42908e-06, 8.447027e-06, 
    8.445567e-06, 8.462753e-06, 8.457213e-06, 8.498517e-06, 8.476321e-06, 
    8.539387e-06, 8.562433e-06, 8.62755e-06, 8.667512e-06, 8.708214e-06, 
    8.726188e-06, 8.731659e-06, 8.733939e-06,
  4.945794e-06, 4.982928e-06, 4.9757e-06, 5.005711e-06, 4.989054e-06, 
    5.008717e-06, 4.953313e-06, 4.984406e-06, 4.964547e-06, 4.94913e-06, 
    5.064138e-06, 5.00705e-06, 5.123663e-06, 5.087079e-06, 5.179147e-06, 
    5.117965e-06, 5.191513e-06, 5.177374e-06, 5.219959e-06, 5.207747e-06, 
    5.262356e-06, 5.225599e-06, 5.290734e-06, 5.253567e-06, 5.259377e-06, 
    5.224389e-06, 5.018516e-06, 5.05702e-06, 5.016239e-06, 5.021722e-06, 
    5.019261e-06, 4.989399e-06, 4.974377e-06, 4.942957e-06, 4.948655e-06, 
    4.971733e-06, 5.024188e-06, 5.006358e-06, 5.051331e-06, 5.050314e-06, 
    5.100549e-06, 5.077878e-06, 5.162569e-06, 5.138448e-06, 5.208256e-06, 
    5.19067e-06, 5.207431e-06, 5.202346e-06, 5.207497e-06, 5.181712e-06, 
    5.192755e-06, 5.170084e-06, 5.082122e-06, 5.10792e-06, 5.031116e-06, 
    4.985139e-06, 4.954676e-06, 4.933102e-06, 4.93615e-06, 4.941963e-06, 
    4.971868e-06, 5.000042e-06, 5.021551e-06, 5.035959e-06, 5.050168e-06, 
    5.093275e-06, 5.116134e-06, 5.167454e-06, 5.158176e-06, 5.173894e-06, 
    5.188921e-06, 5.21419e-06, 5.210027e-06, 5.221171e-06, 5.173477e-06, 
    5.205159e-06, 5.152894e-06, 5.167171e-06, 5.054047e-06, 5.011165e-06, 
    4.99299e-06, 4.97709e-06, 4.938494e-06, 4.965137e-06, 4.954628e-06, 
    4.979639e-06, 4.995557e-06, 4.987681e-06, 5.036353e-06, 5.017411e-06, 
    5.11749e-06, 5.074297e-06, 5.187168e-06, 5.160079e-06, 5.193668e-06, 
    5.176518e-06, 5.205916e-06, 5.179455e-06, 5.225319e-06, 5.235326e-06, 
    5.228487e-06, 5.25477e-06, 5.17799e-06, 5.207432e-06, 4.987461e-06, 
    4.988745e-06, 4.994728e-06, 4.968449e-06, 4.966842e-06, 4.942802e-06, 
    4.964189e-06, 4.973308e-06, 4.996479e-06, 5.010205e-06, 5.023264e-06, 
    5.052021e-06, 5.084207e-06, 5.129331e-06, 5.161834e-06, 5.183661e-06, 
    5.170272e-06, 5.182093e-06, 5.16888e-06, 5.162691e-06, 5.231577e-06, 
    5.192858e-06, 5.250986e-06, 5.247764e-06, 5.221436e-06, 5.248127e-06, 
    4.989647e-06, 4.982258e-06, 4.956641e-06, 4.976685e-06, 4.940186e-06, 
    4.960606e-06, 4.972362e-06, 5.01781e-06, 5.027811e-06, 5.037096e-06, 
    5.055449e-06, 5.079037e-06, 5.120512e-06, 5.156692e-06, 5.189796e-06, 
    5.187368e-06, 5.188223e-06, 5.195628e-06, 5.177292e-06, 5.198641e-06, 
    5.202228e-06, 5.192852e-06, 5.247332e-06, 5.231748e-06, 5.247695e-06, 
    5.237545e-06, 4.984659e-06, 4.997095e-06, 4.990374e-06, 5.003016e-06, 
    4.99411e-06, 5.03376e-06, 5.04567e-06, 5.101527e-06, 5.078573e-06, 
    5.115117e-06, 5.08228e-06, 5.088094e-06, 5.116317e-06, 5.084052e-06, 
    5.154698e-06, 5.10677e-06, 5.195916e-06, 5.147927e-06, 5.198929e-06, 
    5.189652e-06, 5.205013e-06, 5.218785e-06, 5.236126e-06, 5.268179e-06, 
    5.26075e-06, 5.287592e-06, 5.015654e-06, 5.031823e-06, 5.030396e-06, 
    5.047334e-06, 5.059873e-06, 5.087087e-06, 5.130843e-06, 5.114372e-06, 
    5.144622e-06, 5.150703e-06, 5.104751e-06, 5.13295e-06, 5.042652e-06, 
    5.057206e-06, 5.048537e-06, 5.01693e-06, 5.118171e-06, 5.066126e-06, 
    5.162372e-06, 5.134069e-06, 5.216821e-06, 5.175612e-06, 5.256662e-06, 
    5.29145e-06, 5.324248e-06, 5.362679e-06, 5.040652e-06, 5.029657e-06, 
    5.049348e-06, 5.076641e-06, 5.102003e-06, 5.135795e-06, 5.139255e-06, 
    5.145596e-06, 5.162031e-06, 5.175865e-06, 5.147604e-06, 5.179335e-06, 
    5.060588e-06, 5.122695e-06, 5.025505e-06, 5.054706e-06, 5.07503e-06, 
    5.066108e-06, 5.112491e-06, 5.123445e-06, 5.168045e-06, 5.144971e-06, 
    5.282859e-06, 5.221699e-06, 5.391993e-06, 5.34422e-06, 5.025818e-06, 
    5.040613e-06, 5.092229e-06, 5.067647e-06, 5.138052e-06, 5.155435e-06, 
    5.169579e-06, 5.187684e-06, 5.189638e-06, 5.200376e-06, 5.182784e-06, 
    5.19968e-06, 5.135867e-06, 5.164349e-06, 5.086316e-06, 5.105272e-06, 
    5.096548e-06, 5.086986e-06, 5.116517e-06, 5.14805e-06, 5.14872e-06, 
    5.158846e-06, 5.187426e-06, 5.138337e-06, 5.290779e-06, 5.19646e-06, 
    5.056764e-06, 5.085343e-06, 5.089425e-06, 5.078345e-06, 5.153691e-06, 
    5.126346e-06, 5.200114e-06, 5.18014e-06, 5.212879e-06, 5.196602e-06, 
    5.194209e-06, 5.173331e-06, 5.160349e-06, 5.1276e-06, 5.101007e-06, 
    5.079951e-06, 5.084844e-06, 5.107982e-06, 5.149979e-06, 5.189817e-06, 
    5.181082e-06, 5.210389e-06, 5.132935e-06, 5.165366e-06, 5.152824e-06, 
    5.185547e-06, 5.113936e-06, 5.174908e-06, 5.098394e-06, 5.105085e-06, 
    5.125804e-06, 5.167571e-06, 5.176821e-06, 5.186712e-06, 5.180607e-06, 
    5.151046e-06, 5.146207e-06, 5.125299e-06, 5.119534e-06, 5.103628e-06, 
    5.090474e-06, 5.102493e-06, 5.115126e-06, 5.151057e-06, 5.183515e-06, 
    5.218982e-06, 5.227672e-06, 5.269252e-06, 5.235401e-06, 5.291306e-06, 
    5.243773e-06, 5.326144e-06, 5.178443e-06, 5.242369e-06, 5.126746e-06, 
    5.139158e-06, 5.161639e-06, 5.213321e-06, 5.185393e-06, 5.218058e-06, 
    5.146017e-06, 5.108783e-06, 5.09916e-06, 5.081231e-06, 5.09957e-06, 
    5.098078e-06, 5.115646e-06, 5.109998e-06, 5.152252e-06, 5.129539e-06, 
    5.19415e-06, 5.217798e-06, 5.284778e-06, 5.325985e-06, 5.368034e-06, 
    5.386635e-06, 5.392301e-06, 5.39467e-06,
  4.461278e-06, 4.500562e-06, 4.492913e-06, 4.524682e-06, 4.507047e-06, 
    4.527866e-06, 4.46923e-06, 4.502126e-06, 4.481114e-06, 4.464808e-06, 
    4.5866e-06, 4.526101e-06, 4.649783e-06, 4.610943e-06, 4.70876e-06, 
    4.643731e-06, 4.721916e-06, 4.706876e-06, 4.752196e-06, 4.739194e-06, 
    4.797359e-06, 4.758201e-06, 4.827619e-06, 4.787994e-06, 4.794186e-06, 
    4.756912e-06, 4.538247e-06, 4.579051e-06, 4.535835e-06, 4.541643e-06, 
    4.539036e-06, 4.507412e-06, 4.491512e-06, 4.45828e-06, 4.464305e-06, 
    4.488716e-06, 4.544255e-06, 4.525368e-06, 4.573025e-06, 4.571946e-06, 
    4.62524e-06, 4.60118e-06, 4.691131e-06, 4.665492e-06, 4.739737e-06, 
    4.72102e-06, 4.738857e-06, 4.733445e-06, 4.738928e-06, 4.71149e-06, 
    4.723238e-06, 4.699123e-06, 4.605683e-06, 4.633065e-06, 4.551596e-06, 
    4.502901e-06, 4.470671e-06, 4.447861e-06, 4.451083e-06, 4.457228e-06, 
    4.488858e-06, 4.51868e-06, 4.541463e-06, 4.556729e-06, 4.571791e-06, 
    4.617516e-06, 4.641786e-06, 4.696325e-06, 4.68646e-06, 4.703174e-06, 
    4.71916e-06, 4.746052e-06, 4.741621e-06, 4.753485e-06, 4.702731e-06, 
    4.736438e-06, 4.680846e-06, 4.696025e-06, 4.575899e-06, 4.53046e-06, 
    4.511212e-06, 4.494384e-06, 4.453561e-06, 4.481737e-06, 4.470621e-06, 
    4.497083e-06, 4.513931e-06, 4.505594e-06, 4.557146e-06, 4.537076e-06, 
    4.643226e-06, 4.59738e-06, 4.717294e-06, 4.688484e-06, 4.72421e-06, 
    4.705965e-06, 4.737245e-06, 4.70909e-06, 4.757902e-06, 4.76856e-06, 
    4.761276e-06, 4.789276e-06, 4.707531e-06, 4.738858e-06, 4.505361e-06, 
    4.506721e-06, 4.513055e-06, 4.48524e-06, 4.483541e-06, 4.458116e-06, 
    4.480735e-06, 4.490382e-06, 4.514908e-06, 4.529443e-06, 4.543277e-06, 
    4.573755e-06, 4.607894e-06, 4.655805e-06, 4.690349e-06, 4.713564e-06, 
    4.699323e-06, 4.711895e-06, 4.697842e-06, 4.691261e-06, 4.764566e-06, 
    4.723348e-06, 4.785245e-06, 4.781811e-06, 4.753767e-06, 4.782198e-06, 
    4.507675e-06, 4.499855e-06, 4.47275e-06, 4.493956e-06, 4.45535e-06, 
    4.476944e-06, 4.48938e-06, 4.537497e-06, 4.548095e-06, 4.557934e-06, 
    4.57739e-06, 4.60241e-06, 4.646437e-06, 4.684883e-06, 4.72009e-06, 
    4.717507e-06, 4.718416e-06, 4.726296e-06, 4.706788e-06, 4.729502e-06, 
    4.733319e-06, 4.723342e-06, 4.781351e-06, 4.764749e-06, 4.781738e-06, 
    4.770925e-06, 4.502396e-06, 4.515561e-06, 4.508445e-06, 4.52183e-06, 
    4.512399e-06, 4.554397e-06, 4.567021e-06, 4.626276e-06, 4.601917e-06, 
    4.640707e-06, 4.605851e-06, 4.61202e-06, 4.641979e-06, 4.607731e-06, 
    4.682761e-06, 4.631842e-06, 4.726603e-06, 4.675563e-06, 4.729809e-06, 
    4.719938e-06, 4.736284e-06, 4.750945e-06, 4.769412e-06, 4.803568e-06, 
    4.79565e-06, 4.824269e-06, 4.535215e-06, 4.552345e-06, 4.550834e-06, 
    4.568786e-06, 4.582082e-06, 4.610951e-06, 4.657412e-06, 4.639918e-06, 
    4.672053e-06, 4.678516e-06, 4.629702e-06, 4.65965e-06, 4.563823e-06, 
    4.579252e-06, 4.570062e-06, 4.536566e-06, 4.64395e-06, 4.588712e-06, 
    4.690922e-06, 4.66084e-06, 4.748853e-06, 4.705e-06, 4.791294e-06, 
    4.828382e-06, 4.863384e-06, 4.904427e-06, 4.561703e-06, 4.550051e-06, 
    4.570922e-06, 4.599866e-06, 4.626784e-06, 4.662673e-06, 4.66635e-06, 
    4.673088e-06, 4.69056e-06, 4.705271e-06, 4.675222e-06, 4.708962e-06, 
    4.582836e-06, 4.648756e-06, 4.54565e-06, 4.5766e-06, 4.598157e-06, 
    4.588694e-06, 4.63792e-06, 4.649554e-06, 4.696954e-06, 4.672425e-06, 
    4.819219e-06, 4.754046e-06, 4.935764e-06, 4.884707e-06, 4.545983e-06, 
    4.561663e-06, 4.616408e-06, 4.590326e-06, 4.665072e-06, 4.683547e-06, 
    4.698586e-06, 4.717842e-06, 4.719922e-06, 4.731348e-06, 4.71263e-06, 
    4.730608e-06, 4.662749e-06, 4.693024e-06, 4.610135e-06, 4.630254e-06, 
    4.620993e-06, 4.610845e-06, 4.642196e-06, 4.675695e-06, 4.676408e-06, 
    4.687172e-06, 4.717563e-06, 4.665375e-06, 4.827662e-06, 4.727176e-06, 
    4.578786e-06, 4.6091e-06, 4.613433e-06, 4.601676e-06, 4.681693e-06, 
    4.652635e-06, 4.731069e-06, 4.709818e-06, 4.744657e-06, 4.727332e-06, 
    4.724785e-06, 4.702576e-06, 4.688771e-06, 4.653966e-06, 4.625726e-06, 
    4.60338e-06, 4.608572e-06, 4.633132e-06, 4.677746e-06, 4.720112e-06, 
    4.710818e-06, 4.742006e-06, 4.659635e-06, 4.694105e-06, 4.68077e-06, 
    4.71557e-06, 4.639454e-06, 4.704248e-06, 4.622952e-06, 4.630056e-06, 
    4.652059e-06, 4.696448e-06, 4.706288e-06, 4.716809e-06, 4.710315e-06, 
    4.67888e-06, 4.673738e-06, 4.651523e-06, 4.645398e-06, 4.628509e-06, 
    4.614546e-06, 4.627303e-06, 4.640717e-06, 4.678893e-06, 4.713407e-06, 
    4.751154e-06, 4.760409e-06, 4.804709e-06, 4.768638e-06, 4.828225e-06, 
    4.777552e-06, 4.865402e-06, 4.708009e-06, 4.776059e-06, 4.65306e-06, 
    4.666248e-06, 4.690141e-06, 4.745126e-06, 4.715406e-06, 4.750169e-06, 
    4.673536e-06, 4.633981e-06, 4.623766e-06, 4.604738e-06, 4.624202e-06, 
    4.622617e-06, 4.641271e-06, 4.635273e-06, 4.680162e-06, 4.656028e-06, 
    4.724722e-06, 4.749893e-06, 4.821267e-06, 4.865235e-06, 4.910151e-06, 
    4.930035e-06, 4.936093e-06, 4.938627e-06,
  4.331464e-06, 4.372464e-06, 4.364479e-06, 4.397654e-06, 4.379235e-06, 
    4.40098e-06, 4.33976e-06, 4.374097e-06, 4.352161e-06, 4.335146e-06, 
    4.462378e-06, 4.399136e-06, 4.528507e-06, 4.487844e-06, 4.590315e-06, 
    4.52217e-06, 4.604113e-06, 4.588338e-06, 4.635883e-06, 4.622239e-06, 
    4.68331e-06, 4.642187e-06, 4.71511e-06, 4.673472e-06, 4.679976e-06, 
    4.640834e-06, 4.411826e-06, 4.454482e-06, 4.409305e-06, 4.415374e-06, 
    4.41265e-06, 4.379616e-06, 4.363016e-06, 4.328336e-06, 4.334622e-06, 
    4.360096e-06, 4.418105e-06, 4.39837e-06, 4.448179e-06, 4.447051e-06, 
    4.502809e-06, 4.477628e-06, 4.571832e-06, 4.544963e-06, 4.622808e-06, 
    4.603172e-06, 4.621885e-06, 4.616207e-06, 4.621959e-06, 4.593177e-06, 
    4.605499e-06, 4.58021e-06, 4.48234e-06, 4.511001e-06, 4.425776e-06, 
    4.374906e-06, 4.341264e-06, 4.317468e-06, 4.320829e-06, 4.327238e-06, 
    4.360246e-06, 4.391384e-06, 4.415186e-06, 4.431141e-06, 4.446888e-06, 
    4.494724e-06, 4.520133e-06, 4.577276e-06, 4.566935e-06, 4.584457e-06, 
    4.601221e-06, 4.629435e-06, 4.624786e-06, 4.637237e-06, 4.583992e-06, 
    4.619347e-06, 4.561051e-06, 4.576962e-06, 4.451186e-06, 4.40369e-06, 
    4.383584e-06, 4.366013e-06, 4.323414e-06, 4.352812e-06, 4.341211e-06, 
    4.368831e-06, 4.386424e-06, 4.377718e-06, 4.431578e-06, 4.410602e-06, 
    4.521641e-06, 4.473653e-06, 4.599264e-06, 4.569057e-06, 4.606518e-06, 
    4.587384e-06, 4.620194e-06, 4.59066e-06, 4.641874e-06, 4.653062e-06, 
    4.645415e-06, 4.674818e-06, 4.589026e-06, 4.621886e-06, 4.377475e-06, 
    4.378894e-06, 4.385508e-06, 4.356469e-06, 4.354695e-06, 4.328164e-06, 
    4.351766e-06, 4.361836e-06, 4.387444e-06, 4.402627e-06, 4.417082e-06, 
    4.448942e-06, 4.484655e-06, 4.534815e-06, 4.571012e-06, 4.595352e-06, 
    4.580419e-06, 4.593602e-06, 4.578867e-06, 4.571968e-06, 4.648869e-06, 
    4.605614e-06, 4.670584e-06, 4.666977e-06, 4.637533e-06, 4.667383e-06, 
    4.379891e-06, 4.371725e-06, 4.343434e-06, 4.365567e-06, 4.325279e-06, 
    4.34781e-06, 4.360791e-06, 4.411042e-06, 4.422117e-06, 4.432401e-06, 
    4.452743e-06, 4.478915e-06, 4.525003e-06, 4.565282e-06, 4.602197e-06, 
    4.599487e-06, 4.600441e-06, 4.608707e-06, 4.588247e-06, 4.612069e-06, 
    4.616074e-06, 4.605608e-06, 4.666494e-06, 4.649061e-06, 4.6669e-06, 
    4.655545e-06, 4.374378e-06, 4.388126e-06, 4.380695e-06, 4.394674e-06, 
    4.384824e-06, 4.428705e-06, 4.441901e-06, 4.503894e-06, 4.4784e-06, 
    4.519003e-06, 4.482516e-06, 4.488972e-06, 4.520335e-06, 4.484483e-06, 
    4.563059e-06, 4.509721e-06, 4.609028e-06, 4.555516e-06, 4.612391e-06, 
    4.602037e-06, 4.619185e-06, 4.63457e-06, 4.653957e-06, 4.689833e-06, 
    4.681513e-06, 4.711587e-06, 4.408657e-06, 4.426559e-06, 4.42498e-06, 
    4.443747e-06, 4.45765e-06, 4.487853e-06, 4.536498e-06, 4.518176e-06, 
    4.551837e-06, 4.55861e-06, 4.507479e-06, 4.538842e-06, 4.438558e-06, 
    4.454691e-06, 4.445081e-06, 4.410069e-06, 4.522398e-06, 4.464585e-06, 
    4.571612e-06, 4.540088e-06, 4.632375e-06, 4.586373e-06, 4.676937e-06, 
    4.715912e-06, 4.752721e-06, 4.79592e-06, 4.436342e-06, 4.424161e-06, 
    4.44598e-06, 4.476255e-06, 4.504425e-06, 4.542009e-06, 4.545861e-06, 
    4.552922e-06, 4.571233e-06, 4.586656e-06, 4.555158e-06, 4.590526e-06, 
    4.458441e-06, 4.527432e-06, 4.419563e-06, 4.451918e-06, 4.474467e-06, 
    4.464566e-06, 4.516083e-06, 4.528267e-06, 4.577935e-06, 4.552227e-06, 
    4.70628e-06, 4.637826e-06, 4.828927e-06, 4.775161e-06, 4.41991e-06, 
    4.436299e-06, 4.493564e-06, 4.466274e-06, 4.544522e-06, 4.563882e-06, 
    4.579646e-06, 4.599839e-06, 4.60202e-06, 4.614007e-06, 4.594373e-06, 
    4.61323e-06, 4.542089e-06, 4.573816e-06, 4.486998e-06, 4.508058e-06, 
    4.498363e-06, 4.487742e-06, 4.520561e-06, 4.555654e-06, 4.556401e-06, 
    4.567682e-06, 4.599548e-06, 4.54484e-06, 4.715157e-06, 4.609632e-06, 
    4.454203e-06, 4.485916e-06, 4.49045e-06, 4.478147e-06, 4.561939e-06, 
    4.531494e-06, 4.613714e-06, 4.591423e-06, 4.627972e-06, 4.609793e-06, 
    4.607122e-06, 4.58383e-06, 4.569357e-06, 4.532889e-06, 4.503317e-06, 
    4.47993e-06, 4.485363e-06, 4.51107e-06, 4.557803e-06, 4.60222e-06, 
    4.592473e-06, 4.625189e-06, 4.538826e-06, 4.574949e-06, 4.560973e-06, 
    4.597456e-06, 4.51769e-06, 4.585585e-06, 4.500414e-06, 4.50785e-06, 
    4.530891e-06, 4.577406e-06, 4.587722e-06, 4.598755e-06, 4.591945e-06, 
    4.558992e-06, 4.553602e-06, 4.530329e-06, 4.523915e-06, 4.506231e-06, 
    4.491616e-06, 4.504969e-06, 4.519013e-06, 4.559005e-06, 4.595188e-06, 
    4.63479e-06, 4.644504e-06, 4.691032e-06, 4.653145e-06, 4.715749e-06, 
    4.662506e-06, 4.754847e-06, 4.589529e-06, 4.660938e-06, 4.531939e-06, 
    4.545754e-06, 4.570795e-06, 4.628464e-06, 4.597284e-06, 4.633757e-06, 
    4.553391e-06, 4.51196e-06, 4.501265e-06, 4.481351e-06, 4.501721e-06, 
    4.500062e-06, 4.519592e-06, 4.513312e-06, 4.560335e-06, 4.535048e-06, 
    4.607056e-06, 4.633467e-06, 4.708433e-06, 4.75467e-06, 4.801947e-06, 
    4.822891e-06, 4.829274e-06, 4.831944e-06,
  4.364438e-06, 4.405079e-06, 4.397161e-06, 4.430065e-06, 4.411794e-06, 
    4.433366e-06, 4.372658e-06, 4.406699e-06, 4.38495e-06, 4.368085e-06, 
    4.494324e-06, 4.431536e-06, 4.56006e-06, 4.519627e-06, 4.621583e-06, 
    4.553757e-06, 4.635328e-06, 4.619614e-06, 4.666991e-06, 4.653389e-06, 
    4.7143e-06, 4.673276e-06, 4.746046e-06, 4.704481e-06, 4.710972e-06, 
    4.671926e-06, 4.444127e-06, 4.486481e-06, 4.441626e-06, 4.44765e-06, 
    4.444945e-06, 4.412172e-06, 4.395711e-06, 4.361337e-06, 4.367566e-06, 
    4.392816e-06, 4.450359e-06, 4.430776e-06, 4.480217e-06, 4.479097e-06, 
    4.534503e-06, 4.509473e-06, 4.603176e-06, 4.576431e-06, 4.653956e-06, 
    4.63439e-06, 4.653037e-06, 4.647378e-06, 4.653111e-06, 4.624434e-06, 
    4.636708e-06, 4.611518e-06, 4.514156e-06, 4.542649e-06, 4.457975e-06, 
    4.407503e-06, 4.374149e-06, 4.350571e-06, 4.353899e-06, 4.36025e-06, 
    4.392964e-06, 4.423845e-06, 4.447462e-06, 4.4633e-06, 4.478936e-06, 
    4.526467e-06, 4.551731e-06, 4.608597e-06, 4.598301e-06, 4.615748e-06, 
    4.632446e-06, 4.660563e-06, 4.655928e-06, 4.66834e-06, 4.615285e-06, 
    4.650508e-06, 4.592443e-06, 4.608284e-06, 4.483207e-06, 4.436054e-06, 
    4.416109e-06, 4.398683e-06, 4.356461e-06, 4.385594e-06, 4.374097e-06, 
    4.401476e-06, 4.418925e-06, 4.410289e-06, 4.463734e-06, 4.442913e-06, 
    4.553231e-06, 4.505524e-06, 4.630497e-06, 4.600413e-06, 4.637724e-06, 
    4.618662e-06, 4.651351e-06, 4.621926e-06, 4.672963e-06, 4.684121e-06, 
    4.676495e-06, 4.705824e-06, 4.620298e-06, 4.653039e-06, 4.410048e-06, 
    4.411456e-06, 4.418016e-06, 4.38922e-06, 4.387461e-06, 4.361167e-06, 
    4.384558e-06, 4.394541e-06, 4.419936e-06, 4.434999e-06, 4.449344e-06, 
    4.480977e-06, 4.516457e-06, 4.566336e-06, 4.60236e-06, 4.626599e-06, 
    4.611726e-06, 4.624856e-06, 4.61018e-06, 4.603311e-06, 4.67994e-06, 
    4.636824e-06, 4.701599e-06, 4.698001e-06, 4.668636e-06, 4.698406e-06, 
    4.412444e-06, 4.404346e-06, 4.376299e-06, 4.39824e-06, 4.358309e-06, 
    4.380637e-06, 4.393505e-06, 4.44335e-06, 4.454341e-06, 4.464551e-06, 
    4.484751e-06, 4.510753e-06, 4.556574e-06, 4.596655e-06, 4.633418e-06, 
    4.630719e-06, 4.631669e-06, 4.639904e-06, 4.619522e-06, 4.643255e-06, 
    4.647246e-06, 4.636817e-06, 4.697519e-06, 4.680131e-06, 4.697924e-06, 
    4.686597e-06, 4.406977e-06, 4.420612e-06, 4.413242e-06, 4.427109e-06, 
    4.417338e-06, 4.460882e-06, 4.473985e-06, 4.535583e-06, 4.510241e-06, 
    4.550606e-06, 4.514331e-06, 4.520748e-06, 4.551933e-06, 4.516286e-06, 
    4.594443e-06, 4.541377e-06, 4.640224e-06, 4.586936e-06, 4.643576e-06, 
    4.633258e-06, 4.650346e-06, 4.665682e-06, 4.685014e-06, 4.720809e-06, 
    4.712505e-06, 4.742528e-06, 4.440983e-06, 4.458752e-06, 4.457183e-06, 
    4.475816e-06, 4.489625e-06, 4.519635e-06, 4.568009e-06, 4.549783e-06, 
    4.583273e-06, 4.590013e-06, 4.539146e-06, 4.570342e-06, 4.470664e-06, 
    4.486687e-06, 4.477141e-06, 4.442385e-06, 4.553984e-06, 4.496515e-06, 
    4.602957e-06, 4.571581e-06, 4.663494e-06, 4.617656e-06, 4.707939e-06, 
    4.746848e-06, 4.783623e-06, 4.826823e-06, 4.468463e-06, 4.456371e-06, 
    4.478034e-06, 4.50811e-06, 4.53611e-06, 4.573492e-06, 4.577325e-06, 
    4.584352e-06, 4.602579e-06, 4.617938e-06, 4.586578e-06, 4.621792e-06, 
    4.490413e-06, 4.55899e-06, 4.451806e-06, 4.483933e-06, 4.506333e-06, 
    4.496496e-06, 4.547702e-06, 4.55982e-06, 4.609254e-06, 4.58366e-06, 
    4.73723e-06, 4.668929e-06, 4.859856e-06, 4.806057e-06, 4.452151e-06, 
    4.468421e-06, 4.525312e-06, 4.498192e-06, 4.575993e-06, 4.595261e-06, 
    4.610957e-06, 4.63107e-06, 4.633242e-06, 4.645186e-06, 4.625624e-06, 
    4.644411e-06, 4.573572e-06, 4.605151e-06, 4.518785e-06, 4.539722e-06, 
    4.530083e-06, 4.519525e-06, 4.552155e-06, 4.587072e-06, 4.587815e-06, 
    4.599045e-06, 4.630783e-06, 4.576309e-06, 4.746096e-06, 4.640829e-06, 
    4.4862e-06, 4.517711e-06, 4.522217e-06, 4.50999e-06, 4.593328e-06, 
    4.563031e-06, 4.644894e-06, 4.622686e-06, 4.659104e-06, 4.640987e-06, 
    4.638325e-06, 4.615123e-06, 4.600712e-06, 4.564418e-06, 4.535008e-06, 
    4.511761e-06, 4.51716e-06, 4.542717e-06, 4.589211e-06, 4.633441e-06, 
    4.623732e-06, 4.65633e-06, 4.570326e-06, 4.60628e-06, 4.592366e-06, 
    4.628695e-06, 4.549301e-06, 4.616874e-06, 4.532121e-06, 4.539515e-06, 
    4.562431e-06, 4.608728e-06, 4.618999e-06, 4.62999e-06, 4.623205e-06, 
    4.590394e-06, 4.585029e-06, 4.561872e-06, 4.555492e-06, 4.537904e-06, 
    4.523375e-06, 4.53665e-06, 4.550616e-06, 4.590406e-06, 4.626436e-06, 
    4.665901e-06, 4.675586e-06, 4.722008e-06, 4.684205e-06, 4.746687e-06, 
    4.693545e-06, 4.78575e-06, 4.6208e-06, 4.691979e-06, 4.563473e-06, 
    4.577219e-06, 4.602144e-06, 4.659596e-06, 4.628524e-06, 4.664872e-06, 
    4.584819e-06, 4.543603e-06, 4.532968e-06, 4.513173e-06, 4.533421e-06, 
    4.531772e-06, 4.551192e-06, 4.544946e-06, 4.59173e-06, 4.566566e-06, 
    4.63826e-06, 4.664583e-06, 4.739378e-06, 4.785571e-06, 4.832852e-06, 
    4.853813e-06, 4.860203e-06, 4.862876e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.777963, 5.777943, 5.777946, 5.77793, 5.777939, 5.777928, 5.777958, 
    5.777942, 5.777952, 5.777961, 5.777898, 5.777929, 5.777866, 5.777886, 
    5.777837, 5.77787, 5.77783, 5.777838, 5.777815, 5.777822, 5.777792, 
    5.777812, 5.777777, 5.777797, 5.777794, 5.777812, 5.777923, 5.777902, 
    5.777925, 5.777921, 5.777923, 5.777939, 5.777947, 5.777964, 5.777961, 
    5.777948, 5.77792, 5.77793, 5.777905, 5.777906, 5.777879, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.777831, 5.777822, 5.777824, 5.777822, 
    5.777835, 5.777829, 5.777842, 5.777889, 5.777875, 5.777916, 5.777941, 
    5.777958, 5.777969, 5.777968, 5.777965, 5.777948, 5.777933, 5.777922, 
    5.777914, 5.777906, 5.777883, 5.777871, 5.777843, 5.777848, 5.77784, 
    5.777832, 5.777818, 5.77782, 5.777814, 5.77784, 5.777822, 5.777851, 
    5.777843, 5.777904, 5.777927, 5.777937, 5.777946, 5.777966, 5.777952, 
    5.777958, 5.777944, 5.777936, 5.77794, 5.777914, 5.777924, 5.77787, 
    5.777893, 5.777833, 5.777847, 5.777829, 5.777838, 5.777822, 5.777836, 
    5.777812, 5.777807, 5.77781, 5.777796, 5.777837, 5.777822, 5.77794, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777953, 5.777947, 
    5.777935, 5.777927, 5.777921, 5.777905, 5.777888, 5.777864, 5.777846, 
    5.777834, 5.777842, 5.777835, 5.777842, 5.777845, 5.777809, 5.777829, 
    5.777798, 5.7778, 5.777814, 5.7778, 5.777939, 5.777943, 5.777956, 
    5.777946, 5.777966, 5.777955, 5.777948, 5.777924, 5.777918, 5.777913, 
    5.777903, 5.77789, 5.777868, 5.777849, 5.777831, 5.777832, 5.777832, 
    5.777828, 5.777838, 5.777826, 5.777824, 5.777829, 5.7778, 5.777809, 
    5.7778, 5.777805, 5.777942, 5.777935, 5.777938, 5.777932, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.777891, 5.777871, 5.777889, 5.777885, 
    5.77787, 5.777888, 5.77785, 5.777875, 5.777828, 5.777853, 5.777826, 
    5.777831, 5.777823, 5.777815, 5.777806, 5.777789, 5.777793, 5.777779, 
    5.777925, 5.777916, 5.777917, 5.777907, 5.777901, 5.777886, 5.777863, 
    5.777872, 5.777855, 5.777852, 5.777876, 5.777862, 5.77791, 5.777902, 
    5.777907, 5.777924, 5.777869, 5.777897, 5.777846, 5.777861, 5.777816, 
    5.777839, 5.777795, 5.777777, 5.77776, 5.777739, 5.777911, 5.777917, 
    5.777906, 5.777892, 5.777878, 5.77786, 5.777858, 5.777854, 5.777846, 
    5.777838, 5.777853, 5.777836, 5.7779, 5.777867, 5.777919, 5.777904, 
    5.777893, 5.777897, 5.777873, 5.777866, 5.777843, 5.777855, 5.777781, 
    5.777814, 5.777723, 5.777749, 5.777919, 5.777911, 5.777884, 5.777896, 
    5.777859, 5.777849, 5.777842, 5.777832, 5.777831, 5.777825, 5.777835, 
    5.777826, 5.77786, 5.777844, 5.777886, 5.777876, 5.777881, 5.777886, 
    5.77787, 5.777853, 5.777853, 5.777847, 5.777832, 5.777859, 5.777777, 
    5.777827, 5.777903, 5.777887, 5.777885, 5.777891, 5.77785, 5.777865, 
    5.777825, 5.777836, 5.777819, 5.777827, 5.777829, 5.77784, 5.777847, 
    5.777864, 5.777879, 5.77789, 5.777887, 5.777875, 5.777852, 5.777831, 
    5.777836, 5.77782, 5.777862, 5.777844, 5.777851, 5.777833, 5.777872, 
    5.777839, 5.77788, 5.777876, 5.777865, 5.777843, 5.777838, 5.777833, 
    5.777836, 5.777852, 5.777854, 5.777865, 5.777869, 5.777877, 5.777884, 
    5.777878, 5.777871, 5.777852, 5.777834, 5.777815, 5.777811, 5.777789, 
    5.777807, 5.777777, 5.777802, 5.777758, 5.777837, 5.777803, 5.777865, 
    5.777858, 5.777846, 5.777818, 5.777833, 5.777816, 5.777854, 5.777874, 
    5.77788, 5.777889, 5.777879, 5.77788, 5.777871, 5.777874, 5.777851, 
    5.777863, 5.777829, 5.777816, 5.777781, 5.777759, 5.777736, 5.777726, 
    5.777723, 5.777722 ;

 SOIL1C_TO_SOIL2C =
  3.180147e-08, 3.194125e-08, 3.191407e-08, 3.202681e-08, 3.196427e-08, 
    3.203809e-08, 3.182981e-08, 3.19468e-08, 3.187212e-08, 3.181405e-08, 
    3.224559e-08, 3.203184e-08, 3.246759e-08, 3.233128e-08, 3.267369e-08, 
    3.244638e-08, 3.271953e-08, 3.266713e-08, 3.282481e-08, 3.277964e-08, 
    3.298133e-08, 3.284566e-08, 3.308587e-08, 3.294893e-08, 3.297036e-08, 
    3.284119e-08, 3.207485e-08, 3.221898e-08, 3.206631e-08, 3.208687e-08, 
    3.207764e-08, 3.196557e-08, 3.190909e-08, 3.179079e-08, 3.181226e-08, 
    3.189915e-08, 3.209611e-08, 3.202925e-08, 3.219774e-08, 3.219394e-08, 
    3.238152e-08, 3.229694e-08, 3.261221e-08, 3.252261e-08, 3.278153e-08, 
    3.271641e-08, 3.277847e-08, 3.275965e-08, 3.277871e-08, 3.268322e-08, 
    3.272413e-08, 3.26401e-08, 3.231278e-08, 3.240898e-08, 3.212207e-08, 
    3.194954e-08, 3.183494e-08, 3.175362e-08, 3.176511e-08, 3.178703e-08, 
    3.189966e-08, 3.200554e-08, 3.208623e-08, 3.214021e-08, 3.219339e-08, 
    3.235438e-08, 3.243957e-08, 3.263033e-08, 3.25959e-08, 3.265422e-08, 
    3.270993e-08, 3.280347e-08, 3.278808e-08, 3.282929e-08, 3.265268e-08, 
    3.277006e-08, 3.257629e-08, 3.262929e-08, 3.220786e-08, 3.204729e-08, 
    3.197904e-08, 3.19193e-08, 3.177395e-08, 3.187433e-08, 3.183476e-08, 
    3.192889e-08, 3.19887e-08, 3.195912e-08, 3.214168e-08, 3.207071e-08, 
    3.244462e-08, 3.228357e-08, 3.270344e-08, 3.260297e-08, 3.272752e-08, 
    3.266396e-08, 3.277286e-08, 3.267485e-08, 3.284462e-08, 3.288159e-08, 
    3.285633e-08, 3.295337e-08, 3.266942e-08, 3.277847e-08, 3.195829e-08, 
    3.196311e-08, 3.198559e-08, 3.188679e-08, 3.188075e-08, 3.17902e-08, 
    3.187077e-08, 3.190507e-08, 3.199217e-08, 3.204368e-08, 3.209265e-08, 
    3.220032e-08, 3.232056e-08, 3.248869e-08, 3.260948e-08, 3.269044e-08, 
    3.264079e-08, 3.268463e-08, 3.263563e-08, 3.261266e-08, 3.286774e-08, 
    3.272451e-08, 3.293941e-08, 3.292752e-08, 3.283027e-08, 3.292886e-08, 
    3.19665e-08, 3.193874e-08, 3.184234e-08, 3.191778e-08, 3.178034e-08, 
    3.185728e-08, 3.190151e-08, 3.207219e-08, 3.210969e-08, 3.214446e-08, 
    3.221314e-08, 3.230127e-08, 3.245588e-08, 3.259039e-08, 3.271317e-08, 
    3.270418e-08, 3.270734e-08, 3.273478e-08, 3.266683e-08, 3.274593e-08, 
    3.275921e-08, 3.27245e-08, 3.292593e-08, 3.286838e-08, 3.292727e-08, 
    3.28898e-08, 3.194776e-08, 3.199448e-08, 3.196924e-08, 3.20167e-08, 
    3.198326e-08, 3.213196e-08, 3.217655e-08, 3.238515e-08, 3.229954e-08, 
    3.243579e-08, 3.231338e-08, 3.233507e-08, 3.244024e-08, 3.231999e-08, 
    3.258297e-08, 3.240469e-08, 3.273584e-08, 3.255782e-08, 3.2747e-08, 
    3.271265e-08, 3.276952e-08, 3.282047e-08, 3.288455e-08, 3.300281e-08, 
    3.297543e-08, 3.307431e-08, 3.206412e-08, 3.212471e-08, 3.211938e-08, 
    3.218279e-08, 3.222968e-08, 3.233131e-08, 3.249432e-08, 3.243303e-08, 
    3.254556e-08, 3.256815e-08, 3.239718e-08, 3.250216e-08, 3.216526e-08, 
    3.22197e-08, 3.218728e-08, 3.20689e-08, 3.244715e-08, 3.225304e-08, 
    3.261147e-08, 3.250632e-08, 3.28132e-08, 3.266059e-08, 3.296035e-08, 
    3.30885e-08, 3.320909e-08, 3.335003e-08, 3.215778e-08, 3.211661e-08, 
    3.219033e-08, 3.229232e-08, 3.238694e-08, 3.251274e-08, 3.252561e-08, 
    3.254917e-08, 3.261022e-08, 3.266154e-08, 3.255663e-08, 3.267441e-08, 
    3.223233e-08, 3.2464e-08, 3.210105e-08, 3.221034e-08, 3.22863e-08, 
    3.225298e-08, 3.242602e-08, 3.24668e-08, 3.263252e-08, 3.254685e-08, 
    3.305687e-08, 3.283123e-08, 3.345733e-08, 3.328237e-08, 3.210222e-08, 
    3.215764e-08, 3.235049e-08, 3.225873e-08, 3.252113e-08, 3.258572e-08, 
    3.263823e-08, 3.270534e-08, 3.271259e-08, 3.275236e-08, 3.268719e-08, 
    3.274978e-08, 3.2513e-08, 3.261881e-08, 3.232844e-08, 3.239912e-08, 
    3.236661e-08, 3.233094e-08, 3.244101e-08, 3.255828e-08, 3.256078e-08, 
    3.259838e-08, 3.270435e-08, 3.25222e-08, 3.3086e-08, 3.273782e-08, 
    3.221806e-08, 3.23248e-08, 3.234004e-08, 3.229869e-08, 3.257925e-08, 
    3.247759e-08, 3.275139e-08, 3.267739e-08, 3.279863e-08, 3.273838e-08, 
    3.272952e-08, 3.265214e-08, 3.260397e-08, 3.248226e-08, 3.238322e-08, 
    3.230469e-08, 3.232295e-08, 3.240921e-08, 3.256545e-08, 3.271325e-08, 
    3.268087e-08, 3.278942e-08, 3.250211e-08, 3.262258e-08, 3.257602e-08, 
    3.269743e-08, 3.24314e-08, 3.265795e-08, 3.237349e-08, 3.239843e-08, 
    3.247558e-08, 3.263076e-08, 3.266508e-08, 3.270175e-08, 3.267912e-08, 
    3.256942e-08, 3.255144e-08, 3.24737e-08, 3.245224e-08, 3.2393e-08, 
    3.234396e-08, 3.238877e-08, 3.243582e-08, 3.256946e-08, 3.268989e-08, 
    3.282119e-08, 3.285333e-08, 3.300674e-08, 3.288186e-08, 3.308794e-08, 
    3.291274e-08, 3.321601e-08, 3.267107e-08, 3.290758e-08, 3.247909e-08, 
    3.252525e-08, 3.260875e-08, 3.280025e-08, 3.269686e-08, 3.281777e-08, 
    3.255074e-08, 3.24122e-08, 3.237635e-08, 3.230946e-08, 3.237787e-08, 
    3.237231e-08, 3.243777e-08, 3.241673e-08, 3.25739e-08, 3.248948e-08, 
    3.27293e-08, 3.281681e-08, 3.306395e-08, 3.321545e-08, 3.336966e-08, 
    3.343774e-08, 3.345846e-08, 3.346712e-08 ;

 SOIL1C_TO_SOIL3C =
  3.771755e-10, 3.788339e-10, 3.785115e-10, 3.798491e-10, 3.791071e-10, 
    3.799829e-10, 3.775117e-10, 3.788997e-10, 3.780137e-10, 3.773248e-10, 
    3.824449e-10, 3.799087e-10, 3.85079e-10, 3.834616e-10, 3.875244e-10, 
    3.848273e-10, 3.880682e-10, 3.874465e-10, 3.893175e-10, 3.887815e-10, 
    3.911746e-10, 3.895649e-10, 3.924151e-10, 3.907902e-10, 3.910444e-10, 
    3.895118e-10, 3.804191e-10, 3.821291e-10, 3.803178e-10, 3.805616e-10, 
    3.804522e-10, 3.791224e-10, 3.784523e-10, 3.770488e-10, 3.773036e-10, 
    3.783344e-10, 3.806713e-10, 3.79878e-10, 3.818772e-10, 3.81832e-10, 
    3.840576e-10, 3.830542e-10, 3.867948e-10, 3.857317e-10, 3.888039e-10, 
    3.880312e-10, 3.887676e-10, 3.885443e-10, 3.887705e-10, 3.876374e-10, 
    3.881228e-10, 3.871257e-10, 3.832421e-10, 3.843835e-10, 3.809793e-10, 
    3.789323e-10, 3.775726e-10, 3.766078e-10, 3.767442e-10, 3.770042e-10, 
    3.783404e-10, 3.795967e-10, 3.805541e-10, 3.811945e-10, 3.818255e-10, 
    3.837356e-10, 3.847464e-10, 3.870098e-10, 3.866013e-10, 3.872933e-10, 
    3.879544e-10, 3.890643e-10, 3.888816e-10, 3.893706e-10, 3.87275e-10, 
    3.886678e-10, 3.863687e-10, 3.869975e-10, 3.819972e-10, 3.80092e-10, 
    3.792823e-10, 3.785735e-10, 3.768491e-10, 3.780399e-10, 3.775705e-10, 
    3.786873e-10, 3.793969e-10, 3.790459e-10, 3.81212e-10, 3.803699e-10, 
    3.848064e-10, 3.828955e-10, 3.878773e-10, 3.866852e-10, 3.88163e-10, 
    3.874089e-10, 3.88701e-10, 3.875381e-10, 3.895526e-10, 3.899912e-10, 
    3.896914e-10, 3.908429e-10, 3.874737e-10, 3.887676e-10, 3.790361e-10, 
    3.790933e-10, 3.7936e-10, 3.781878e-10, 3.781161e-10, 3.770418e-10, 
    3.779977e-10, 3.784048e-10, 3.79438e-10, 3.800492e-10, 3.806303e-10, 
    3.819077e-10, 3.833344e-10, 3.853293e-10, 3.867625e-10, 3.877231e-10, 
    3.87134e-10, 3.876541e-10, 3.870727e-10, 3.868002e-10, 3.898269e-10, 
    3.881274e-10, 3.906773e-10, 3.905362e-10, 3.893822e-10, 3.905521e-10, 
    3.791335e-10, 3.788041e-10, 3.776605e-10, 3.785555e-10, 3.769248e-10, 
    3.778376e-10, 3.783625e-10, 3.803876e-10, 3.808324e-10, 3.81245e-10, 
    3.820598e-10, 3.831055e-10, 3.849399e-10, 3.865359e-10, 3.879928e-10, 
    3.878861e-10, 3.879237e-10, 3.882492e-10, 3.874429e-10, 3.883815e-10, 
    3.885391e-10, 3.881272e-10, 3.905173e-10, 3.898344e-10, 3.905332e-10, 
    3.900886e-10, 3.789112e-10, 3.794655e-10, 3.79166e-10, 3.797292e-10, 
    3.793324e-10, 3.810967e-10, 3.816257e-10, 3.841008e-10, 3.83085e-10, 
    3.847016e-10, 3.832492e-10, 3.835065e-10, 3.847544e-10, 3.833276e-10, 
    3.86448e-10, 3.843325e-10, 3.882618e-10, 3.861494e-10, 3.883942e-10, 
    3.879865e-10, 3.886614e-10, 3.892659e-10, 3.900263e-10, 3.914295e-10, 
    3.911046e-10, 3.922779e-10, 3.802917e-10, 3.810107e-10, 3.809474e-10, 
    3.816997e-10, 3.822561e-10, 3.83462e-10, 3.853961e-10, 3.846688e-10, 
    3.86004e-10, 3.86272e-10, 3.842435e-10, 3.85489e-10, 3.814918e-10, 
    3.821377e-10, 3.817531e-10, 3.803485e-10, 3.848364e-10, 3.825333e-10, 
    3.867861e-10, 3.855385e-10, 3.891797e-10, 3.873689e-10, 3.909257e-10, 
    3.924462e-10, 3.938772e-10, 3.955495e-10, 3.81403e-10, 3.809145e-10, 
    3.817892e-10, 3.829993e-10, 3.84122e-10, 3.856146e-10, 3.857673e-10, 
    3.860469e-10, 3.867712e-10, 3.873802e-10, 3.861354e-10, 3.875328e-10, 
    3.822875e-10, 3.850363e-10, 3.807299e-10, 3.820267e-10, 3.829279e-10, 
    3.825326e-10, 3.845856e-10, 3.850696e-10, 3.870359e-10, 3.860194e-10, 
    3.92071e-10, 3.893936e-10, 3.968228e-10, 3.947467e-10, 3.807439e-10, 
    3.814013e-10, 3.836895e-10, 3.826008e-10, 3.857142e-10, 3.864806e-10, 
    3.871035e-10, 3.878999e-10, 3.879859e-10, 3.884577e-10, 3.876845e-10, 
    3.884272e-10, 3.856178e-10, 3.868732e-10, 3.834279e-10, 3.842665e-10, 
    3.838807e-10, 3.834576e-10, 3.847636e-10, 3.86155e-10, 3.861846e-10, 
    3.866308e-10, 3.878881e-10, 3.857268e-10, 3.924167e-10, 3.882853e-10, 
    3.821182e-10, 3.833847e-10, 3.835655e-10, 3.830749e-10, 3.864037e-10, 
    3.851976e-10, 3.884462e-10, 3.875682e-10, 3.890068e-10, 3.88292e-10, 
    3.881868e-10, 3.872687e-10, 3.86697e-10, 3.852529e-10, 3.840779e-10, 
    3.83146e-10, 3.833627e-10, 3.843863e-10, 3.862401e-10, 3.879937e-10, 
    3.876096e-10, 3.888975e-10, 3.854885e-10, 3.869179e-10, 3.863655e-10, 
    3.87806e-10, 3.846495e-10, 3.873376e-10, 3.839624e-10, 3.842583e-10, 
    3.851737e-10, 3.870149e-10, 3.874222e-10, 3.878572e-10, 3.875888e-10, 
    3.862871e-10, 3.860738e-10, 3.851514e-10, 3.848968e-10, 3.841938e-10, 
    3.836119e-10, 3.841436e-10, 3.84702e-10, 3.862876e-10, 3.877166e-10, 
    3.892745e-10, 3.896558e-10, 3.914762e-10, 3.899943e-10, 3.924397e-10, 
    3.903608e-10, 3.939594e-10, 3.874933e-10, 3.902996e-10, 3.852153e-10, 
    3.85763e-10, 3.867538e-10, 3.89026e-10, 3.877993e-10, 3.892339e-10, 
    3.860655e-10, 3.844216e-10, 3.839963e-10, 3.832027e-10, 3.840144e-10, 
    3.839484e-10, 3.847251e-10, 3.844755e-10, 3.863403e-10, 3.853386e-10, 
    3.881842e-10, 3.892226e-10, 3.92155e-10, 3.939526e-10, 3.957825e-10, 
    3.965903e-10, 3.968362e-10, 3.96939e-10 ;

 SOIL1C_vr =
  19.97935, 19.9793, 19.97931, 19.97927, 19.97929, 19.97926, 19.97934, 
    19.9793, 19.97932, 19.97935, 19.97918, 19.97926, 19.9791, 19.97915, 
    19.97902, 19.9791, 19.979, 19.97902, 19.97896, 19.97898, 19.9789, 
    19.97895, 19.97886, 19.97891, 19.9789, 19.97895, 19.97925, 19.97919, 
    19.97925, 19.97924, 19.97925, 19.97929, 19.97931, 19.97936, 19.97935, 
    19.97931, 19.97924, 19.97926, 19.9792, 19.9792, 19.97913, 19.97916, 
    19.97904, 19.97907, 19.97898, 19.979, 19.97898, 19.97898, 19.97898, 
    19.97901, 19.979, 19.97903, 19.97915, 19.97912, 19.97923, 19.97929, 
    19.97934, 19.97937, 19.97937, 19.97936, 19.97931, 19.97927, 19.97924, 
    19.97922, 19.9792, 19.97914, 19.9791, 19.97903, 19.97905, 19.97902, 
    19.979, 19.97897, 19.97897, 19.97896, 19.97902, 19.97898, 19.97905, 
    19.97903, 19.97919, 19.97926, 19.97928, 19.97931, 19.97936, 19.97932, 
    19.97934, 19.9793, 19.97928, 19.97929, 19.97922, 19.97925, 19.9791, 
    19.97917, 19.979, 19.97904, 19.97899, 19.97902, 19.97898, 19.97902, 
    19.97895, 19.97894, 19.97895, 19.97891, 19.97902, 19.97898, 19.97929, 
    19.97929, 19.97928, 19.97932, 19.97932, 19.97936, 19.97932, 19.97931, 
    19.97928, 19.97926, 19.97924, 19.9792, 19.97915, 19.97909, 19.97904, 
    19.97901, 19.97903, 19.97901, 19.97903, 19.97904, 19.97894, 19.979, 
    19.97891, 19.97892, 19.97896, 19.97892, 19.97929, 19.9793, 19.97934, 
    19.97931, 19.97936, 19.97933, 19.97931, 19.97925, 19.97923, 19.97922, 
    19.97919, 19.97916, 19.9791, 19.97905, 19.979, 19.979, 19.979, 19.97899, 
    19.97902, 19.97899, 19.97898, 19.979, 19.97892, 19.97894, 19.97892, 
    19.97893, 19.9793, 19.97928, 19.97929, 19.97927, 19.97928, 19.97923, 
    19.97921, 19.97913, 19.97916, 19.97911, 19.97915, 19.97915, 19.9791, 
    19.97915, 19.97905, 19.97912, 19.97899, 19.97906, 19.97899, 19.979, 
    19.97898, 19.97896, 19.97894, 19.97889, 19.9789, 19.97886, 19.97925, 
    19.97923, 19.97923, 19.9792, 19.97919, 19.97915, 19.97908, 19.97911, 
    19.97906, 19.97906, 19.97912, 19.97908, 19.97921, 19.97919, 19.9792, 
    19.97925, 19.9791, 19.97918, 19.97904, 19.97908, 19.97896, 19.97902, 
    19.97891, 19.97886, 19.97881, 19.97876, 19.97921, 19.97923, 19.9792, 
    19.97916, 19.97913, 19.97908, 19.97907, 19.97906, 19.97904, 19.97902, 
    19.97906, 19.97902, 19.97919, 19.9791, 19.97924, 19.97919, 19.97916, 
    19.97918, 19.97911, 19.9791, 19.97903, 19.97906, 19.97887, 19.97896, 
    19.97872, 19.97878, 19.97924, 19.97921, 19.97914, 19.97918, 19.97907, 
    19.97905, 19.97903, 19.979, 19.979, 19.97898, 19.97901, 19.97899, 
    19.97908, 19.97904, 19.97915, 19.97912, 19.97913, 19.97915, 19.9791, 
    19.97906, 19.97906, 19.97904, 19.979, 19.97907, 19.97886, 19.97899, 
    19.97919, 19.97915, 19.97915, 19.97916, 19.97905, 19.97909, 19.97899, 
    19.97902, 19.97897, 19.97899, 19.97899, 19.97902, 19.97904, 19.97909, 
    19.97913, 19.97916, 19.97915, 19.97912, 19.97906, 19.979, 19.97901, 
    19.97897, 19.97908, 19.97904, 19.97905, 19.97901, 19.97911, 19.97902, 
    19.97913, 19.97912, 19.97909, 19.97903, 19.97902, 19.97901, 19.97901, 
    19.97906, 19.97906, 19.97909, 19.9791, 19.97912, 19.97914, 19.97913, 
    19.97911, 19.97906, 19.97901, 19.97896, 19.97895, 19.97889, 19.97894, 
    19.97886, 19.97892, 19.97881, 19.97902, 19.97893, 19.97909, 19.97907, 
    19.97904, 19.97897, 19.97901, 19.97896, 19.97906, 19.97912, 19.97913, 
    19.97916, 19.97913, 19.97913, 19.97911, 19.97911, 19.97905, 19.97909, 
    19.97899, 19.97896, 19.97887, 19.97881, 19.97875, 19.97872, 19.97872, 
    19.97871,
  19.98101, 19.98094, 19.98095, 19.98089, 19.98092, 19.98089, 19.98099, 
    19.98093, 19.98097, 19.981, 19.98078, 19.98089, 19.98067, 19.98074, 
    19.98057, 19.98068, 19.98054, 19.98057, 19.98049, 19.98051, 19.98041, 
    19.98048, 19.98036, 19.98043, 19.98042, 19.98048, 19.98087, 19.98079, 
    19.98087, 19.98086, 19.98087, 19.98092, 19.98095, 19.98101, 19.981, 
    19.98096, 19.98086, 19.98089, 19.98081, 19.98081, 19.98071, 19.98076, 
    19.9806, 19.98064, 19.98051, 19.98054, 19.98051, 19.98052, 19.98051, 
    19.98056, 19.98054, 19.98058, 19.98075, 19.9807, 19.98084, 19.98093, 
    19.98099, 19.98103, 19.98103, 19.98101, 19.98096, 19.9809, 19.98086, 
    19.98083, 19.98081, 19.98073, 19.98068, 19.98059, 19.9806, 19.98058, 
    19.98055, 19.9805, 19.98051, 19.98049, 19.98058, 19.98052, 19.98061, 
    19.98059, 19.9808, 19.98088, 19.98092, 19.98095, 19.98102, 19.98097, 
    19.98099, 19.98094, 19.98091, 19.98093, 19.98083, 19.98087, 19.98068, 
    19.98076, 19.98055, 19.9806, 19.98054, 19.98057, 19.98051, 19.98056, 
    19.98048, 19.98046, 19.98047, 19.98042, 19.98057, 19.98051, 19.98093, 
    19.98092, 19.98091, 19.98096, 19.98097, 19.98101, 19.98097, 19.98096, 
    19.98091, 19.98088, 19.98086, 19.9808, 19.98074, 19.98066, 19.9806, 
    19.98056, 19.98058, 19.98056, 19.98059, 19.9806, 19.98047, 19.98054, 
    19.98043, 19.98044, 19.98049, 19.98044, 19.98092, 19.98094, 19.98099, 
    19.98095, 19.98102, 19.98098, 19.98096, 19.98087, 19.98085, 19.98083, 
    19.9808, 19.98075, 19.98067, 19.98061, 19.98055, 19.98055, 19.98055, 
    19.98053, 19.98057, 19.98053, 19.98052, 19.98054, 19.98044, 19.98047, 
    19.98044, 19.98046, 19.98093, 19.98091, 19.98092, 19.9809, 19.98092, 
    19.98084, 19.98082, 19.98071, 19.98075, 19.98069, 19.98075, 19.98074, 
    19.98068, 19.98074, 19.98061, 19.9807, 19.98053, 19.98062, 19.98053, 
    19.98055, 19.98052, 19.98049, 19.98046, 19.9804, 19.98041, 19.98036, 
    19.98087, 19.98084, 19.98085, 19.98081, 19.98079, 19.98074, 19.98066, 
    19.98069, 19.98063, 19.98062, 19.98071, 19.98065, 19.98082, 19.98079, 
    19.98081, 19.98087, 19.98068, 19.98078, 19.9806, 19.98065, 19.9805, 
    19.98057, 19.98042, 19.98036, 19.9803, 19.98022, 19.98083, 19.98085, 
    19.98081, 19.98076, 19.98071, 19.98065, 19.98064, 19.98063, 19.9806, 
    19.98057, 19.98063, 19.98056, 19.98079, 19.98067, 19.98086, 19.9808, 
    19.98076, 19.98078, 19.98069, 19.98067, 19.98059, 19.98063, 19.98037, 
    19.98049, 19.98017, 19.98026, 19.98085, 19.98083, 19.98073, 19.98078, 
    19.98064, 19.98061, 19.98058, 19.98055, 19.98055, 19.98053, 19.98056, 
    19.98053, 19.98065, 19.98059, 19.98074, 19.9807, 19.98072, 19.98074, 
    19.98068, 19.98062, 19.98062, 19.9806, 19.98055, 19.98064, 19.98036, 
    19.98053, 19.98079, 19.98074, 19.98073, 19.98075, 19.98061, 19.98067, 
    19.98053, 19.98056, 19.9805, 19.98053, 19.98054, 19.98058, 19.9806, 
    19.98066, 19.98071, 19.98075, 19.98074, 19.9807, 19.98062, 19.98055, 
    19.98056, 19.98051, 19.98065, 19.98059, 19.98061, 19.98055, 19.98069, 
    19.98057, 19.98072, 19.98071, 19.98067, 19.98059, 19.98057, 19.98055, 
    19.98056, 19.98062, 19.98063, 19.98067, 19.98068, 19.98071, 19.98073, 
    19.98071, 19.98069, 19.98062, 19.98056, 19.98049, 19.98047, 19.9804, 
    19.98046, 19.98036, 19.98044, 19.98029, 19.98057, 19.98045, 19.98066, 
    19.98064, 19.9806, 19.9805, 19.98055, 19.98049, 19.98063, 19.9807, 
    19.98071, 19.98075, 19.98071, 19.98072, 19.98068, 19.9807, 19.98062, 
    19.98066, 19.98054, 19.98049, 19.98037, 19.98029, 19.98022, 19.98018, 
    19.98017, 19.98017,
  19.98273, 19.98265, 19.98267, 19.98261, 19.98264, 19.9826, 19.98271, 
    19.98265, 19.98269, 19.98272, 19.98249, 19.9826, 19.98237, 19.98244, 
    19.98226, 19.98238, 19.98223, 19.98226, 19.98217, 19.9822, 19.98209, 
    19.98216, 19.98203, 19.98211, 19.9821, 19.98217, 19.98258, 19.9825, 
    19.98258, 19.98257, 19.98258, 19.98264, 19.98267, 19.98273, 19.98272, 
    19.98268, 19.98257, 19.9826, 19.98251, 19.98252, 19.98241, 19.98246, 
    19.98229, 19.98234, 19.9822, 19.98223, 19.9822, 19.98221, 19.9822, 
    19.98225, 19.98223, 19.98228, 19.98245, 19.9824, 19.98255, 19.98265, 
    19.98271, 19.98275, 19.98275, 19.98274, 19.98268, 19.98262, 19.98257, 
    19.98254, 19.98252, 19.98243, 19.98238, 19.98228, 19.9823, 19.98227, 
    19.98224, 19.98219, 19.98219, 19.98217, 19.98227, 19.9822, 19.98231, 
    19.98228, 19.98251, 19.9826, 19.98263, 19.98266, 19.98274, 19.98269, 
    19.98271, 19.98266, 19.98263, 19.98264, 19.98254, 19.98258, 19.98238, 
    19.98247, 19.98224, 19.98229, 19.98223, 19.98226, 19.9822, 19.98226, 
    19.98216, 19.98214, 19.98216, 19.98211, 19.98226, 19.9822, 19.98264, 
    19.98264, 19.98263, 19.98268, 19.98269, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.9826, 19.98257, 19.98251, 19.98245, 19.98236, 19.98229, 
    19.98225, 19.98227, 19.98225, 19.98228, 19.98229, 19.98215, 19.98223, 
    19.98211, 19.98212, 19.98217, 19.98212, 19.98264, 19.98265, 19.98271, 
    19.98266, 19.98274, 19.9827, 19.98267, 19.98258, 19.98256, 19.98254, 
    19.98251, 19.98246, 19.98237, 19.9823, 19.98223, 19.98224, 19.98224, 
    19.98222, 19.98226, 19.98222, 19.98221, 19.98223, 19.98212, 19.98215, 
    19.98212, 19.98214, 19.98265, 19.98262, 19.98264, 19.98261, 19.98263, 
    19.98255, 19.98252, 19.98241, 19.98246, 19.98238, 19.98245, 19.98244, 
    19.98238, 19.98245, 19.98231, 19.9824, 19.98222, 19.98232, 19.98222, 
    19.98223, 19.9822, 19.98218, 19.98214, 19.98208, 19.98209, 19.98204, 
    19.98259, 19.98255, 19.98256, 19.98252, 19.9825, 19.98244, 19.98235, 
    19.98239, 19.98232, 19.98231, 19.9824, 19.98235, 19.98253, 19.9825, 
    19.98252, 19.98258, 19.98238, 19.98248, 19.98229, 19.98235, 19.98218, 
    19.98226, 19.9821, 19.98203, 19.98197, 19.98189, 19.98253, 19.98256, 
    19.98252, 19.98246, 19.98241, 19.98234, 19.98234, 19.98232, 19.98229, 
    19.98226, 19.98232, 19.98226, 19.98249, 19.98237, 19.98256, 19.98251, 
    19.98247, 19.98248, 19.98239, 19.98237, 19.98228, 19.98232, 19.98205, 
    19.98217, 19.98183, 19.98193, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98234, 19.9823, 19.98228, 19.98224, 19.98223, 19.98221, 19.98225, 
    19.98222, 19.98234, 19.98229, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98232, 19.98232, 19.9823, 19.98224, 19.98234, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98244, 19.98246, 19.98231, 19.98236, 
    19.98221, 19.98225, 19.98219, 19.98222, 19.98223, 19.98227, 19.98229, 
    19.98236, 19.98241, 19.98246, 19.98244, 19.9824, 19.98232, 19.98223, 
    19.98225, 19.98219, 19.98235, 19.98228, 19.98231, 19.98224, 19.98239, 
    19.98227, 19.98242, 19.9824, 19.98236, 19.98228, 19.98226, 19.98224, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98238, 19.98241, 19.98243, 
    19.98241, 19.98238, 19.98231, 19.98225, 19.98218, 19.98216, 19.98208, 
    19.98214, 19.98203, 19.98213, 19.98196, 19.98226, 19.98213, 19.98236, 
    19.98234, 19.98229, 19.98219, 19.98224, 19.98218, 19.98232, 19.9824, 
    19.98242, 19.98245, 19.98242, 19.98242, 19.98238, 19.9824, 19.98231, 
    19.98236, 19.98223, 19.98218, 19.98205, 19.98196, 19.98188, 19.98184, 
    19.98183, 19.98183,
  19.9841, 19.98403, 19.98404, 19.98398, 19.98401, 19.98397, 19.98409, 
    19.98402, 19.98406, 19.9841, 19.98386, 19.98398, 19.98375, 19.98382, 
    19.98363, 19.98376, 19.98361, 19.98364, 19.98355, 19.98358, 19.98347, 
    19.98354, 19.98341, 19.98349, 19.98347, 19.98355, 19.98396, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98405, 19.98411, 19.9841, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98384, 
    19.98367, 19.98372, 19.98358, 19.98361, 19.98358, 19.98359, 19.98358, 
    19.98363, 19.98361, 19.98365, 19.98383, 19.98378, 19.98393, 19.98402, 
    19.98409, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98366, 19.98368, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98365, 19.98358, 19.98369, 
    19.98366, 19.98388, 19.98397, 19.98401, 19.98404, 19.98412, 19.98406, 
    19.98409, 19.98403, 19.984, 19.98402, 19.98392, 19.98396, 19.98376, 
    19.98384, 19.98362, 19.98367, 19.98361, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98354, 19.98348, 19.98364, 19.98358, 19.98402, 
    19.98402, 19.984, 19.98406, 19.98406, 19.98411, 19.98407, 19.98405, 
    19.984, 19.98397, 19.98395, 19.98389, 19.98382, 19.98373, 19.98367, 
    19.98363, 19.98365, 19.98363, 19.98365, 19.98367, 19.98353, 19.98361, 
    19.98349, 19.9835, 19.98355, 19.9835, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98396, 19.98394, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98362, 19.98362, 
    19.9836, 19.98364, 19.98359, 19.98359, 19.98361, 19.9835, 19.98353, 
    19.9835, 19.98352, 19.98402, 19.984, 19.98401, 19.98399, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98384, 19.98376, 19.98383, 19.98382, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.9837, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98346, 19.98347, 19.98342, 
    19.98396, 19.98393, 19.98393, 19.9839, 19.98387, 19.98382, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98373, 19.98391, 19.98388, 
    19.98389, 19.98396, 19.98376, 19.98386, 19.98367, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98335, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.9837, 19.98363, 19.98387, 19.98375, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98377, 19.98375, 19.98366, 19.9837, 19.98343, 
    19.98355, 19.98322, 19.98331, 19.98394, 19.98391, 19.98381, 19.98386, 
    19.98372, 19.98368, 19.98365, 19.98362, 19.98361, 19.98359, 19.98363, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98382, 
    19.98376, 19.9837, 19.98369, 19.98368, 19.98362, 19.98372, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98384, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98357, 19.9836, 19.9836, 19.98365, 19.98367, 
    19.98374, 19.98379, 19.98383, 19.98382, 19.98378, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98373, 19.98366, 19.98369, 19.98362, 19.98376, 
    19.98364, 19.9838, 19.98378, 19.98374, 19.98366, 19.98364, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98379, 19.98381, 
    19.98379, 19.98376, 19.98369, 19.98363, 19.98355, 19.98354, 19.98346, 
    19.98352, 19.98341, 19.98351, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98357, 19.98362, 19.98356, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.9838, 19.98376, 19.98377, 19.98369, 
    19.98373, 19.9836, 19.98356, 19.98343, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.98571, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98558, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98529, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98564, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98522, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98565, 19.98562, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98527, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98567, 19.98567, 19.98571, 19.98567, 19.98566, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98522, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98572, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98528, 
    19.98526, 19.98529, 19.98526, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98563, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98535, 19.98526, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98556, 19.98553, 19.9855, 19.98545, 19.98538, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98554, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.9853, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98548, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98522, 19.98492, 19.985, 19.98556, 19.98554, 19.98545, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98528, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98535, 19.98534, 19.98533, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98534, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98542, 19.98534, 19.98527, 
    19.98529, 19.98524, 19.98537, 19.98532, 19.98534, 19.98528, 19.98541, 
    19.9853, 19.98543, 19.98542, 19.98539, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98539, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98518, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98493, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222428, 0.7222433, 0.7222413, 0.7222424, 0.722241, 0.7222448, 
    0.7222427, 0.722244, 0.7222451, 0.7222373, 0.7222412, 0.7222333, 
    0.7222357, 0.7222296, 0.7222337, 0.7222288, 0.7222297, 0.7222269, 
    0.7222277, 0.7222241, 0.7222265, 0.7222221, 0.7222246, 0.7222242, 
    0.7222266, 0.7222404, 0.7222378, 0.7222406, 0.7222401, 0.7222403, 
    0.7222424, 0.7222434, 0.7222455, 0.7222452, 0.7222435, 0.72224, 
    0.7222412, 0.7222382, 0.7222382, 0.7222348, 0.7222364, 0.7222307, 
    0.7222323, 0.7222276, 0.7222288, 0.7222277, 0.7222281, 0.7222277, 
    0.7222294, 0.7222286, 0.7222302, 0.7222361, 0.7222344, 0.7222396, 
    0.7222427, 0.7222447, 0.7222462, 0.722246, 0.7222456, 0.7222435, 
    0.7222416, 0.7222402, 0.7222392, 0.7222382, 0.7222353, 0.7222338, 
    0.7222304, 0.722231, 0.72223, 0.7222289, 0.7222272, 0.7222275, 0.7222268, 
    0.72223, 0.7222278, 0.7222313, 0.7222304, 0.722238, 0.7222409, 0.7222421, 
    0.7222432, 0.7222458, 0.722244, 0.7222447, 0.722243, 0.7222419, 
    0.7222425, 0.7222392, 0.7222404, 0.7222337, 0.7222366, 0.7222291, 
    0.7222309, 0.7222286, 0.7222298, 0.7222278, 0.7222295, 0.7222265, 
    0.7222258, 0.7222263, 0.7222245, 0.7222297, 0.7222277, 0.7222425, 
    0.7222424, 0.722242, 0.7222438, 0.7222439, 0.7222455, 0.7222441, 
    0.7222434, 0.7222419, 0.7222409, 0.7222401, 0.7222381, 0.722236, 
    0.7222329, 0.7222307, 0.7222293, 0.7222302, 0.7222294, 0.7222303, 
    0.7222307, 0.7222261, 0.7222286, 0.7222248, 0.722225, 0.7222267, 
    0.722225, 0.7222424, 0.7222428, 0.7222446, 0.7222432, 0.7222457, 
    0.7222443, 0.7222435, 0.7222404, 0.7222397, 0.7222391, 0.7222379, 
    0.7222363, 0.7222335, 0.7222311, 0.7222289, 0.722229, 0.7222289, 
    0.7222285, 0.7222297, 0.7222283, 0.7222281, 0.7222286, 0.722225, 
    0.7222261, 0.722225, 0.7222257, 0.7222427, 0.7222418, 0.7222423, 
    0.7222415, 0.7222421, 0.7222394, 0.7222385, 0.7222348, 0.7222363, 
    0.7222339, 0.7222361, 0.7222357, 0.7222338, 0.722236, 0.7222312, 
    0.7222344, 0.7222285, 0.7222317, 0.7222282, 0.7222289, 0.7222279, 
    0.7222269, 0.7222258, 0.7222236, 0.7222241, 0.7222223, 0.7222406, 
    0.7222395, 0.7222396, 0.7222384, 0.7222376, 0.7222357, 0.7222328, 
    0.722234, 0.7222319, 0.7222315, 0.7222345, 0.7222327, 0.7222388, 
    0.7222378, 0.7222384, 0.7222405, 0.7222337, 0.7222372, 0.7222307, 
    0.7222326, 0.722227, 0.7222298, 0.7222244, 0.7222221, 0.7222199, 
    0.7222174, 0.7222389, 0.7222396, 0.7222383, 0.7222365, 0.7222348, 
    0.7222325, 0.7222323, 0.7222318, 0.7222307, 0.7222298, 0.7222317, 
    0.7222295, 0.7222375, 0.7222334, 0.7222399, 0.7222379, 0.7222366, 
    0.7222372, 0.7222341, 0.7222333, 0.7222303, 0.7222319, 0.7222227, 
    0.7222267, 0.7222154, 0.7222186, 0.7222399, 0.7222389, 0.7222354, 
    0.7222371, 0.7222323, 0.7222311, 0.7222302, 0.722229, 0.7222289, 
    0.7222282, 0.7222294, 0.7222282, 0.7222325, 0.7222306, 0.7222358, 
    0.7222345, 0.7222351, 0.7222357, 0.7222338, 0.7222317, 0.7222316, 
    0.7222309, 0.722229, 0.7222323, 0.7222221, 0.7222284, 0.7222378, 
    0.7222359, 0.7222356, 0.7222363, 0.7222313, 0.7222331, 0.7222282, 
    0.7222295, 0.7222273, 0.7222284, 0.7222286, 0.72223, 0.7222309, 
    0.7222331, 0.7222348, 0.7222362, 0.7222359, 0.7222344, 0.7222315, 
    0.7222289, 0.7222295, 0.7222275, 0.7222327, 0.7222305, 0.7222313, 
    0.7222291, 0.722234, 0.7222298, 0.722235, 0.7222345, 0.7222332, 
    0.7222304, 0.7222297, 0.7222291, 0.7222295, 0.7222314, 0.7222318, 
    0.7222332, 0.7222336, 0.7222347, 0.7222356, 0.7222347, 0.7222339, 
    0.7222314, 0.7222293, 0.7222269, 0.7222263, 0.7222236, 0.7222258, 
    0.7222221, 0.7222252, 0.7222198, 0.7222296, 0.7222254, 0.7222331, 
    0.7222323, 0.7222307, 0.7222273, 0.7222292, 0.722227, 0.7222318, 
    0.7222343, 0.722235, 0.7222362, 0.7222349, 0.722235, 0.7222338, 
    0.7222342, 0.7222314, 0.7222329, 0.7222286, 0.722227, 0.7222226, 
    0.7222198, 0.722217, 0.7222158, 0.7222154, 0.7222153 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  5.139921e-21, 1.027984e-20, 0, 4.111937e-20, -2.569961e-20, 0, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 1.541976e-20, 
    -3.083953e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, -1.541976e-20, 
    2.006177e-36, 5.139921e-21, 1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, 
    -2.055969e-20, -2.569961e-20, 1.541976e-20, -2.569961e-20, 2.569961e-20, 
    1.027984e-20, -1.541976e-20, 2.569961e-20, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, 2.055969e-20, 3.083953e-20, -1.027984e-20, -3.083953e-20, 
    1.027984e-20, 0, 1.027984e-20, 2.055969e-20, 3.083953e-20, 5.139921e-21, 
    5.139921e-21, 3.083953e-20, -5.139921e-21, -3.597945e-20, -5.139921e-21, 
    -2.569961e-20, 2.055969e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 3.597945e-20, 3.083953e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 1.541976e-20, 
    -3.597945e-20, -1.541976e-20, -4.625929e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 2.055969e-20, 1.541976e-20, 4.111937e-20, 
    -2.055969e-20, -2.569961e-20, 2.055969e-20, -2.569961e-20, -2.055969e-20, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 0, 
    -2.569961e-20, 2.569961e-20, 5.139921e-21, -2.006177e-36, -5.139921e-21, 
    -2.055969e-20, 5.139921e-21, 5.139921e-20, 5.139921e-21, -1.541976e-20, 
    1.027984e-20, -2.055969e-20, 2.055969e-20, -5.139921e-21, 2.055969e-20, 
    -1.541976e-20, -2.569961e-20, 3.597945e-20, 3.597945e-20, -1.027984e-20, 
    1.541976e-20, 5.653913e-20, -5.139921e-21, 3.083953e-20, -1.027984e-20, 
    -1.027984e-20, -3.597945e-20, 2.006177e-36, 0, 2.055969e-20, 
    -1.027984e-20, 1.541976e-20, -2.006177e-36, 1.027984e-20, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, 4.625929e-20, 5.139921e-21, 5.139921e-21, 
    1.541976e-20, 2.055969e-20, -2.006177e-36, -5.139921e-21, 3.083953e-20, 
    0, 2.055969e-20, -5.139921e-21, -3.083953e-20, -5.139921e-21, 
    -3.083953e-20, 1.541976e-20, 5.139921e-21, 2.569961e-20, -1.027984e-20, 
    3.083953e-20, 1.027984e-20, 1.541976e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 2.055969e-20, -4.625929e-20, -1.027984e-20, -2.006177e-36, 
    1.027984e-20, 2.569961e-20, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -3.597945e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -4.625929e-20, 2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 1.027984e-20, -1.027984e-20, 2.569961e-20, 
    -1.027984e-20, 2.569961e-20, 2.055969e-20, -5.139921e-21, -4.625929e-20, 
    -1.541976e-20, 5.139921e-21, -2.569961e-20, 2.006177e-36, -3.083953e-20, 
    5.139921e-21, 2.055969e-20, 1.027984e-20, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, -3.597945e-20, 1.541976e-20, 
    -2.055969e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, -1.541976e-20, 
    2.569961e-20, -2.055969e-20, -2.055969e-20, 0, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, -5.139921e-21, 0, 
    -5.139921e-21, 1.541976e-20, 0, 3.083953e-20, 2.055969e-20, 1.027984e-20, 
    2.055969e-20, 2.006177e-36, -1.027984e-20, -3.597945e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, 1.541976e-20, 
    -1.027984e-20, 0, -5.139921e-21, -3.597945e-20, -2.055969e-20, 
    2.569961e-20, 0, 5.139921e-21, 2.055969e-20, -5.139921e-21, 3.083953e-20, 
    -5.139921e-21, 1.027984e-20, -2.055969e-20, 1.027984e-20, 0, 
    2.055969e-20, 5.139921e-21, -2.055969e-20, -5.139921e-21, -1.541976e-20, 
    2.569961e-20, -3.083953e-20, -1.541976e-20, 2.055969e-20, 2.006177e-36, 
    -5.139921e-21, -2.055969e-20, 2.006177e-36, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, -3.083953e-20, -5.139921e-21, 
    2.055969e-20, -5.139921e-21, -1.027984e-20, 2.006177e-36, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, 3.597945e-20, 3.083953e-20, 5.139921e-21, 
    -3.083953e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, -3.083953e-20, 
    2.055969e-20, 5.139921e-21, 0, -5.139921e-20, -1.027984e-20, 
    -1.541976e-20, -1.541976e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, -2.006177e-36, 0, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    -2.569961e-20, -1.541976e-20, 2.055969e-20, 1.027984e-20, 0, 
    -1.541976e-20, -2.055969e-20, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -1.027984e-20, -5.139921e-21, 2.569961e-20, 
    -2.055969e-20, 2.055969e-20, -1.027984e-20, 2.055969e-20, 2.006177e-36, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21,
  2.055969e-20, -2.055969e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    1.541976e-20, -2.055969e-20, -1.541976e-20, 2.569961e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, -2.569961e-20, 
    1.027984e-20, -2.055969e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -3.083953e-20, 0, -1.027984e-20, 0, 1.541976e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -2.006177e-36, -5.139921e-21, -1.541976e-20, 
    -1.541976e-20, 2.006177e-36, -2.055969e-20, 2.006177e-36, 0, 0, 
    -1.541976e-20, -5.139921e-21, -1.541976e-20, 0, -2.569961e-20, 
    -2.055969e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -3.083953e-20, 0, -5.139921e-21, -1.027984e-20, 3.597945e-20, 
    1.027984e-20, 1.541976e-20, 2.006177e-36, 0, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 
    -2.055969e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 2.006177e-36, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, 
    1.541976e-20, -3.083953e-20, 3.083953e-20, -1.541976e-20, 0, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, -1.027984e-20, 2.569961e-20, 
    -5.139921e-21, -2.055969e-20, -2.569961e-20, -2.055969e-20, 1.541976e-20, 
    2.569961e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 2.006177e-36, 
    5.139921e-21, 1.541976e-20, 1.541976e-20, -2.055969e-20, -2.055969e-20, 
    -2.569961e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 0, 
    5.139921e-21, -5.139921e-21, -2.006177e-36, 2.569961e-20, 2.569961e-20, 
    1.541976e-20, -5.139921e-21, 2.055969e-20, -1.027984e-20, -2.569961e-20, 
    0, 5.139921e-21, -5.139921e-21, -1.541976e-20, 1.541976e-20, 
    2.569961e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, -2.055969e-20, 1.541976e-20, -2.006177e-36, 
    -1.027984e-20, 2.006177e-36, -1.027984e-20, -2.569961e-20, 0, 
    -3.597945e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    2.569961e-20, -1.027984e-20, 0, 1.541976e-20, 2.006177e-36, 1.027984e-20, 
    -3.083953e-20, -2.055969e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 0, 1.541976e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 2.569961e-20, -1.027984e-20, 0, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    0, -5.139921e-21, -3.083953e-20, 1.541976e-20, 1.541976e-20, 
    1.027984e-20, 0, 5.139921e-21, -5.139921e-21, -3.083953e-20, 
    -5.139921e-21, 1.027984e-20, 4.111937e-20, 5.139921e-21, -5.139921e-21, 
    0, 5.139921e-21, 1.541976e-20, 2.055969e-20, -2.569961e-20, 1.541976e-20, 
    1.541976e-20, 2.006177e-36, 1.027984e-20, -1.541976e-20, 0, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 2.569961e-20, -5.139921e-21, -1.027984e-20, 
    2.055969e-20, -5.139921e-21, 1.027984e-20, -3.597945e-20, 0, 
    5.139921e-21, -3.083953e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 1.541976e-20, -1.541976e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -2.569961e-20, -2.055969e-20, 0, 1.541976e-20, -2.055969e-20, 0, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    0, -3.083953e-20, 0, -5.139921e-21, 2.055969e-20, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -2.055969e-20, 1.541976e-20, 1.541976e-20, 
    0, -5.139921e-21, 0, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 2.055969e-20, 2.055969e-20, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 0, 2.569961e-20, 5.139921e-21, 2.569961e-20, 
    1.541976e-20, 0, 1.541976e-20, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, -4.111937e-20, -1.541976e-20, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, 0, 1.027984e-20, 
    -2.055969e-20, -1.541976e-20, 1.541976e-20, 0, 1.027984e-20, 
    -2.006177e-36, 2.006177e-36, 1.541976e-20, 2.569961e-20, 2.055969e-20, 0, 
    5.139921e-21, -5.139921e-21, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    2.055969e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 2.569961e-20, 
    -5.139921e-21, 2.006177e-36, 3.597945e-20, 2.055969e-20, -3.083953e-20, 
    -1.027984e-20, 3.083953e-20, 2.055969e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, 2.055969e-20, -1.541976e-20, 
    -2.569961e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 0, 2.569961e-20, 1.027984e-20, 
    -3.083953e-20, -1.027984e-20, 2.055969e-20, 0, 5.139921e-21, 1.027984e-20,
  -2.055969e-20, 1.541976e-20, -1.027984e-20, -2.006177e-36, 3.083953e-20, 
    1.027984e-20, -5.139921e-21, -3.597945e-20, -3.597945e-20, -2.055969e-20, 
    0, -5.139921e-21, 5.139921e-21, -2.569961e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    0, -3.597945e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 0, 1.027984e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, 
    2.569961e-20, -1.541976e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 0, 
    2.055969e-20, -5.139921e-21, 5.139921e-21, -5.139921e-21, 3.083953e-20, 
    -5.139921e-21, 0, -4.625929e-20, 1.027984e-20, 3.083953e-20, 
    5.139921e-21, -2.055969e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-20, 0, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -2.055969e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, 0, 3.083953e-20, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 0, -1.541976e-20, 0, 5.139921e-21, -5.139921e-21, 0, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 2.006177e-36, 0, 
    1.541976e-20, 5.139921e-21, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    -2.569961e-20, -1.541976e-20, -1.541976e-20, -4.625929e-20, 
    -2.569961e-20, 5.139921e-21, 1.541976e-20, -2.006177e-36, -1.541976e-20, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 0, 
    -3.083953e-20, -3.597945e-20, -1.541976e-20, 1.027984e-20, -5.139921e-21, 
    0, 5.139921e-21, 5.139921e-21, -1.541976e-20, 3.597945e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, 2.006177e-36, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -2.055969e-20, 
    -2.055969e-20, 1.027984e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-20, -1.027984e-20, 2.055969e-20, 
    -1.027984e-20, 0, -1.541976e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -3.083953e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -3.083953e-20, 2.569961e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 0, -1.541976e-20, -5.139921e-21, 
    1.541976e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -3.083953e-20, -3.083953e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, -3.083953e-20, -5.139921e-21, 1.541976e-20, 
    -2.569961e-20, -2.006177e-36, -1.541976e-20, -1.541976e-20, 
    -1.027984e-20, 0, 1.027984e-20, -2.569961e-20, 5.139921e-21, 
    2.006177e-36, 2.569961e-20, -1.027984e-20, -1.541976e-20, -3.083953e-20, 
    -1.541976e-20, 0, -1.027984e-20, -2.055969e-20, -2.055969e-20, 
    1.541976e-20, -1.541976e-20, -2.055969e-20, -1.541976e-20, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, -2.055969e-20, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 0, 0, -1.027984e-20, 0, 
    -3.083953e-20, 2.055969e-20, -5.139921e-21, -2.055969e-20, -2.569961e-20, 
    1.027984e-20, -5.139921e-21, -3.083953e-20, -1.027984e-20, -3.597945e-20, 
    -2.006177e-36, 5.139921e-21, -1.027984e-20, -5.139921e-21, 2.006177e-36, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 2.055969e-20, -1.027984e-20, 
    0, 0, -5.139921e-21, 0, 1.541976e-20, -1.027984e-20, 0, 3.083953e-20, 
    -3.083953e-20, 5.139921e-21, -3.597945e-20, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 2.055969e-20, 0, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, 0, -3.597945e-20, 
    -1.027984e-20, 0, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -3.083953e-20, -1.027984e-20, -1.541976e-20, -2.055969e-20, 
    -5.139921e-21, -3.083953e-20, 1.027984e-20, 0, -2.006177e-36, 
    5.139921e-21, -3.083953e-20, -1.541976e-20, -2.569961e-20, 2.569961e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -3.083953e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -2.006177e-36, 0, -1.027984e-20, 5.139921e-21, 0, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, -2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -2.006177e-36, 5.139921e-21, 2.055969e-20, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 3.597945e-20, -5.139921e-21, -1.541976e-20, -1.541976e-20, 
    2.055969e-20, -5.139921e-21, 2.055969e-20, -2.569961e-20, 0, 
    -1.027984e-20, 2.006177e-36, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 0, 2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21,
  5.139921e-21, 2.006177e-36, 2.569961e-20, 0, 1.027984e-20, 1.027984e-20, 
    2.055969e-20, 5.139921e-21, 2.055969e-20, 2.006177e-36, 0, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, -3.597945e-20, -2.006177e-36, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-20, -1.541976e-20, 2.055969e-20, 0, 0, -2.055969e-20, 
    5.139921e-21, 1.027984e-20, 3.083953e-20, -2.055969e-20, -1.541976e-20, 
    0, 1.027984e-20, 2.006177e-36, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, 3.597945e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 1.027984e-20, -3.597945e-20, -2.569961e-20, 
    5.139921e-21, -2.055969e-20, -2.055969e-20, 1.027984e-20, -3.083953e-20, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-20, 5.139921e-21, 
    5.139921e-21, 3.083953e-20, 4.625929e-20, 0, 2.055969e-20, 5.139921e-20, 
    -1.027984e-20, -2.006177e-36, -1.541976e-20, 2.569961e-20, 1.027984e-20, 
    2.055969e-20, -2.055969e-20, 2.006177e-36, 1.541976e-20, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -1.541976e-20, 3.083953e-20, 2.569961e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, -2.569961e-20, -2.569961e-20, 
    5.139921e-21, -4.111937e-20, -2.569961e-20, -2.055969e-20, 4.625929e-20, 
    2.569961e-20, -1.027984e-20, -1.541976e-20, -3.083953e-20, 2.055969e-20, 
    -3.597945e-20, 5.139921e-21, -1.027984e-20, 3.083953e-20, -5.139921e-21, 
    1.027984e-20, -2.055969e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    3.083953e-20, -1.541976e-20, 5.139921e-21, 2.006177e-36, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 1.541976e-20, 2.006177e-36, 0, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, -2.569961e-20, 5.139921e-21, 
    2.569961e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, -3.083953e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -3.083953e-20, 2.006177e-36, 
    0, -1.027984e-20, 2.055969e-20, -1.027984e-20, -2.055969e-20, 
    -2.055969e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, -4.625929e-20, 
    -2.006177e-36, 1.541976e-20, -2.055969e-20, 1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 1.027984e-20, -2.006177e-36, 2.569961e-20, 0, 
    -1.541976e-20, 1.027984e-20, 1.027984e-20, 2.055969e-20, -2.055969e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 2.055969e-20, 4.111937e-20, 
    5.139921e-21, -2.569961e-20, 1.027984e-20, 5.653913e-20, -2.006177e-36, 
    2.006177e-36, 1.027984e-20, -2.055969e-20, -5.139921e-21, -1.027984e-20, 
    2.569961e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -3.597945e-20, 1.027984e-20, 2.055969e-20, 1.027984e-20, 2.055969e-20, 
    1.541976e-20, 2.569961e-20, -5.139921e-21, -1.027984e-20, 3.083953e-20, 
    1.027984e-20, 3.083953e-20, -1.027984e-20, -2.055969e-20, 3.083953e-20, 
    3.083953e-20, 2.569961e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 5.139921e-21, -4.111937e-20, 5.139921e-21, 
    1.027984e-20, 2.006177e-36, -2.006177e-36, -3.083953e-20, 2.055969e-20, 
    3.083953e-20, -3.083953e-20, 4.111937e-20, 5.139921e-21, -2.055969e-20, 
    -1.027984e-20, -4.111937e-20, -3.083953e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 2.006177e-36, -5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -1.541976e-20, 1.541976e-20, 3.597945e-20, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 3.083953e-20, 
    2.055969e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -2.055969e-20, -2.569961e-20, -5.139921e-21, 2.569961e-20, 0, 0, 0, 
    -2.055969e-20, 3.083953e-20, -2.006177e-36, -5.139921e-21, -1.027984e-20, 
    3.083953e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 2.055969e-20, 
    -5.139921e-21, 2.569961e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.569961e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 2.055969e-20, 5.139921e-21, -4.111937e-20, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, -2.569961e-20, 5.139921e-21, 
    2.569961e-20, -2.569961e-20, -1.027984e-20, 2.569961e-20, 2.055969e-20, 
    1.027984e-20, -2.055969e-20, -3.083953e-20, 2.055969e-20, 1.027984e-20, 
    3.083953e-20, 1.027984e-20, -2.055969e-20, -1.541976e-20, -1.027984e-20, 
    4.111937e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 0, 
    -1.027984e-20, 2.006177e-36, -5.139921e-21, 3.597945e-20, 2.055969e-20, 
    5.139921e-21, 2.055969e-20, -1.027984e-20, 1.027984e-20, 0, 
    -2.055969e-20, 3.597945e-20,
  -5.139921e-21, 2.569961e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, 0, 1.541976e-20, -2.055969e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, -2.006177e-36, 
    -1.541976e-20, 2.569961e-20, 1.027984e-20, 2.055969e-20, 0, 0, 
    1.027984e-20, -2.006177e-36, 1.027984e-20, -2.006177e-36, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    -3.083953e-20, -5.139921e-21, -1.541976e-20, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-20, 1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-20, 2.055969e-20, 0, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    -1.027984e-20, 2.055969e-20, -5.139921e-21, 3.597945e-20, 2.006177e-36, 
    -1.541976e-20, 1.027984e-20, 5.139921e-21, 3.083953e-20, 1.541976e-20, 
    2.055969e-20, -2.055969e-20, 2.569961e-20, 1.027984e-20, 2.569961e-20, 
    2.569961e-20, 0, 4.625929e-20, 1.541976e-20, -2.569961e-20, 
    -1.541976e-20, -1.027984e-20, 0, -1.541976e-20, 0, -1.541976e-20, 
    1.027984e-20, 2.055969e-20, 1.027984e-20, 1.027984e-20, -2.569961e-20, 
    -5.139921e-21, -1.541976e-20, -1.541976e-20, -1.027984e-20, 1.027984e-20, 
    -2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, -2.569961e-20, 
    -5.139921e-21, -1.027984e-20, -3.597945e-20, -2.055969e-20, 1.541976e-20, 
    -3.597945e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, -2.006177e-36, 
    -1.027984e-20, 2.006177e-36, -1.541976e-20, -1.027984e-20, 0, 
    1.027984e-20, -1.541976e-20, 2.569961e-20, 1.541976e-20, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, 0, 2.055969e-20, -3.597945e-20, 5.139921e-21, 
    2.569961e-20, -1.541976e-20, -2.569961e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, -2.569961e-20, 5.139921e-21, -2.569961e-20, -1.027984e-20, 
    0, 0, 0, 1.027984e-20, 1.541976e-20, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 0, 
    -1.027984e-20, -2.055969e-20, -1.541976e-20, 3.083953e-20, -5.139921e-21, 
    -1.027984e-20, 4.111937e-20, 2.006177e-36, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, -2.006177e-36, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, -1.541976e-20, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, 0, 
    1.027984e-20, 1.541976e-20, 1.027984e-20, -5.653913e-20, 0, 
    -2.055969e-20, 2.055969e-20, 0, 1.027984e-20, 0, 1.027984e-20, 0, 
    5.139921e-21, 1.541976e-20, -2.055969e-20, -1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 1.027984e-20, 
    1.541976e-20, 5.139921e-21, -3.083953e-20, 3.083953e-20, 1.541976e-20, 
    1.541976e-20, 1.541976e-20, 1.541976e-20, 1.541976e-20, -2.006177e-36, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, 3.083953e-20, 2.055969e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, 1.541976e-20, 0, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 1.027984e-20, -4.625929e-20, 1.541976e-20, -1.541976e-20, 
    -1.027984e-20, 0, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.055969e-20, -1.027984e-20, -2.006177e-36, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 3.597945e-20, -3.083953e-20, 
    1.027984e-20, 1.541976e-20, 0, -5.139921e-21, -2.569961e-20, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 0, 2.006177e-36, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 0, 1.541976e-20, -2.055969e-20, 
    2.569961e-20, -5.139921e-21, -5.139921e-21, 2.569961e-20, 2.055969e-20, 
    1.541976e-20, -3.083953e-20, -2.006177e-36, -5.139921e-21, 3.597945e-20, 
    2.569961e-20, 5.139921e-21, 0, -5.139921e-21, -5.139921e-21, 
    -2.055969e-20, -4.625929e-20, -1.541976e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, -2.006177e-36, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    5.139921e-21, 0, -2.055969e-20, 2.006177e-36, -1.027984e-20, 0, 
    2.055969e-20, -2.055969e-20, 1.027984e-20, 1.541976e-20, -2.055969e-20, 
    1.027984e-20, -5.139921e-21, 3.083953e-20, 2.006177e-36, -2.569961e-20, 
    -4.111937e-20, -2.006177e-36, 5.139921e-21, 4.111937e-20, -1.027984e-20, 
    5.139921e-21, 0, 1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, -2.006177e-36, -1.027984e-20, 
    -1.541976e-20,
  8.598664e-29, 8.598635e-29, 8.598641e-29, 8.598618e-29, 8.59863e-29, 
    8.598615e-29, 8.598658e-29, 8.598634e-29, 8.598649e-29, 8.598662e-29, 
    8.598573e-29, 8.598617e-29, 8.598527e-29, 8.598556e-29, 8.598485e-29, 
    8.598532e-29, 8.598476e-29, 8.598486e-29, 8.598454e-29, 8.598463e-29, 
    8.598422e-29, 8.59845e-29, 8.5984e-29, 8.598429e-29, 8.598424e-29, 
    8.598451e-29, 8.598608e-29, 8.598578e-29, 8.59861e-29, 8.598606e-29, 
    8.598607e-29, 8.59863e-29, 8.598642e-29, 8.598666e-29, 8.598662e-29, 
    8.598644e-29, 8.598604e-29, 8.598617e-29, 8.598583e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598498e-29, 8.598516e-29, 8.598463e-29, 
    8.598476e-29, 8.598463e-29, 8.598468e-29, 8.598463e-29, 8.598483e-29, 
    8.598475e-29, 8.598492e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598674e-29, 8.598671e-29, 8.598667e-29, 
    8.598643e-29, 8.598622e-29, 8.598606e-29, 8.598595e-29, 8.598584e-29, 
    8.598551e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598478e-29, 8.598459e-29, 8.598462e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598505e-29, 8.598494e-29, 8.598581e-29, 8.598613e-29, 
    8.598627e-29, 8.59864e-29, 8.598669e-29, 8.598649e-29, 8.598657e-29, 
    8.598638e-29, 8.598625e-29, 8.598631e-29, 8.598594e-29, 8.598609e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.5985e-29, 8.598474e-29, 
    8.598487e-29, 8.598465e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598448e-29, 8.598427e-29, 8.598486e-29, 8.598463e-29, 8.598632e-29, 
    8.598631e-29, 8.598626e-29, 8.598646e-29, 8.598648e-29, 8.598666e-29, 
    8.598649e-29, 8.598643e-29, 8.598625e-29, 8.598614e-29, 8.598604e-29, 
    8.598582e-29, 8.598557e-29, 8.598523e-29, 8.598498e-29, 8.598482e-29, 
    8.598492e-29, 8.598483e-29, 8.598493e-29, 8.598498e-29, 8.598445e-29, 
    8.598475e-29, 8.59843e-29, 8.598433e-29, 8.598453e-29, 8.598433e-29, 
    8.59863e-29, 8.598636e-29, 8.598655e-29, 8.59864e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598609e-29, 8.598601e-29, 8.598593e-29, 
    8.59858e-29, 8.598562e-29, 8.59853e-29, 8.598502e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598473e-29, 8.598486e-29, 8.59847e-29, 
    8.598468e-29, 8.598475e-29, 8.598433e-29, 8.598445e-29, 8.598433e-29, 
    8.598441e-29, 8.598634e-29, 8.598624e-29, 8.59863e-29, 8.59862e-29, 
    8.598627e-29, 8.598596e-29, 8.598587e-29, 8.598544e-29, 8.598562e-29, 
    8.598534e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598504e-29, 8.598541e-29, 8.598473e-29, 8.598509e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598455e-29, 8.598442e-29, 8.598418e-29, 
    8.598423e-29, 8.598403e-29, 8.59861e-29, 8.598598e-29, 8.598599e-29, 
    8.598586e-29, 8.598576e-29, 8.598556e-29, 8.598522e-29, 8.598535e-29, 
    8.598512e-29, 8.598507e-29, 8.598542e-29, 8.59852e-29, 8.598589e-29, 
    8.598578e-29, 8.598585e-29, 8.598609e-29, 8.598532e-29, 8.598571e-29, 
    8.598498e-29, 8.598519e-29, 8.598456e-29, 8.598488e-29, 8.598426e-29, 
    8.5984e-29, 8.598375e-29, 8.598346e-29, 8.598591e-29, 8.5986e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598488e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598528e-29, 8.598603e-29, 8.59858e-29, 8.598565e-29, 
    8.598571e-29, 8.598536e-29, 8.598527e-29, 8.598494e-29, 8.598511e-29, 
    8.598406e-29, 8.598453e-29, 8.598324e-29, 8.59836e-29, 8.598603e-29, 
    8.598591e-29, 8.598551e-29, 8.59857e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598479e-29, 8.598477e-29, 8.598469e-29, 8.598482e-29, 
    8.59847e-29, 8.598518e-29, 8.598497e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598556e-29, 8.598533e-29, 8.598509e-29, 8.598508e-29, 
    8.598501e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598472e-29, 
    8.598578e-29, 8.598557e-29, 8.598554e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598469e-29, 8.598485e-29, 8.598459e-29, 8.598472e-29, 
    8.598474e-29, 8.598489e-29, 8.5985e-29, 8.598524e-29, 8.598545e-29, 
    8.598561e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598477e-29, 
    8.598483e-29, 8.598461e-29, 8.59852e-29, 8.598495e-29, 8.598505e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598547e-29, 8.598542e-29, 
    8.598525e-29, 8.598494e-29, 8.598487e-29, 8.598479e-29, 8.598484e-29, 
    8.598506e-29, 8.59851e-29, 8.598526e-29, 8.59853e-29, 8.598543e-29, 
    8.598553e-29, 8.598544e-29, 8.598534e-29, 8.598506e-29, 8.598482e-29, 
    8.598455e-29, 8.598448e-29, 8.598417e-29, 8.598442e-29, 8.5984e-29, 
    8.598436e-29, 8.598374e-29, 8.598486e-29, 8.598437e-29, 8.598525e-29, 
    8.598516e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598456e-29, 
    8.59851e-29, 8.598539e-29, 8.598546e-29, 8.59856e-29, 8.598546e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598506e-29, 8.598523e-29, 
    8.598474e-29, 8.598456e-29, 8.598405e-29, 8.598374e-29, 8.598342e-29, 
    8.598328e-29, 8.598324e-29, 8.598322e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.164853e-08, 1.169975e-08, 1.168979e-08, 1.17311e-08, 1.170818e-08, 
    1.173523e-08, 1.165891e-08, 1.170178e-08, 1.167441e-08, 1.165314e-08, 
    1.181126e-08, 1.173294e-08, 1.189261e-08, 1.184266e-08, 1.196814e-08, 
    1.188484e-08, 1.198493e-08, 1.196573e-08, 1.202351e-08, 1.200696e-08, 
    1.208087e-08, 1.203115e-08, 1.211918e-08, 1.2069e-08, 1.207685e-08, 
    1.202951e-08, 1.17487e-08, 1.180151e-08, 1.174557e-08, 1.17531e-08, 
    1.174972e-08, 1.170866e-08, 1.168796e-08, 1.164461e-08, 1.165248e-08, 
    1.168432e-08, 1.175649e-08, 1.173199e-08, 1.179373e-08, 1.179234e-08, 
    1.186107e-08, 1.183008e-08, 1.194561e-08, 1.191277e-08, 1.200765e-08, 
    1.198379e-08, 1.200653e-08, 1.199964e-08, 1.200662e-08, 1.197163e-08, 
    1.198662e-08, 1.195583e-08, 1.183589e-08, 1.187114e-08, 1.1766e-08, 
    1.170279e-08, 1.166079e-08, 1.163099e-08, 1.163521e-08, 1.164324e-08, 
    1.168451e-08, 1.17233e-08, 1.175287e-08, 1.177265e-08, 1.179214e-08, 
    1.185113e-08, 1.188234e-08, 1.195225e-08, 1.193963e-08, 1.1961e-08, 
    1.198142e-08, 1.201569e-08, 1.201005e-08, 1.202515e-08, 1.196044e-08, 
    1.200345e-08, 1.193244e-08, 1.195187e-08, 1.179744e-08, 1.17386e-08, 
    1.171359e-08, 1.16917e-08, 1.163845e-08, 1.167522e-08, 1.166073e-08, 
    1.169522e-08, 1.171713e-08, 1.170629e-08, 1.177319e-08, 1.174718e-08, 
    1.188419e-08, 1.182518e-08, 1.197904e-08, 1.194222e-08, 1.198786e-08, 
    1.196457e-08, 1.200448e-08, 1.196856e-08, 1.203077e-08, 1.204432e-08, 
    1.203506e-08, 1.207062e-08, 1.196657e-08, 1.200653e-08, 1.170599e-08, 
    1.170776e-08, 1.171599e-08, 1.167979e-08, 1.167758e-08, 1.16444e-08, 
    1.167392e-08, 1.168649e-08, 1.17184e-08, 1.173728e-08, 1.175522e-08, 
    1.179468e-08, 1.183874e-08, 1.190035e-08, 1.194461e-08, 1.197427e-08, 
    1.195608e-08, 1.197214e-08, 1.195419e-08, 1.194577e-08, 1.203925e-08, 
    1.198676e-08, 1.206551e-08, 1.206115e-08, 1.202551e-08, 1.206164e-08, 
    1.1709e-08, 1.169883e-08, 1.166351e-08, 1.169115e-08, 1.164079e-08, 
    1.166898e-08, 1.168519e-08, 1.174773e-08, 1.176147e-08, 1.177421e-08, 
    1.179937e-08, 1.183167e-08, 1.188832e-08, 1.193761e-08, 1.198261e-08, 
    1.197931e-08, 1.198047e-08, 1.199052e-08, 1.196562e-08, 1.199461e-08, 
    1.199947e-08, 1.198675e-08, 1.206057e-08, 1.203948e-08, 1.206106e-08, 
    1.204733e-08, 1.170213e-08, 1.171925e-08, 1.171e-08, 1.17274e-08, 
    1.171514e-08, 1.176963e-08, 1.178597e-08, 1.18624e-08, 1.183103e-08, 
    1.188096e-08, 1.18361e-08, 1.184405e-08, 1.188259e-08, 1.183853e-08, 
    1.193489e-08, 1.186956e-08, 1.199091e-08, 1.192567e-08, 1.1995e-08, 
    1.198241e-08, 1.200325e-08, 1.202192e-08, 1.204541e-08, 1.208874e-08, 
    1.207871e-08, 1.211494e-08, 1.174477e-08, 1.176697e-08, 1.176502e-08, 
    1.178825e-08, 1.180543e-08, 1.184268e-08, 1.190241e-08, 1.187995e-08, 
    1.192118e-08, 1.192946e-08, 1.186681e-08, 1.190528e-08, 1.178183e-08, 
    1.180178e-08, 1.17899e-08, 1.174652e-08, 1.188512e-08, 1.181399e-08, 
    1.194534e-08, 1.190681e-08, 1.201926e-08, 1.196334e-08, 1.207318e-08, 
    1.212014e-08, 1.216433e-08, 1.221598e-08, 1.177909e-08, 1.1764e-08, 
    1.179101e-08, 1.182839e-08, 1.186306e-08, 1.190916e-08, 1.191387e-08, 
    1.192251e-08, 1.194488e-08, 1.196368e-08, 1.192524e-08, 1.19684e-08, 
    1.18064e-08, 1.18913e-08, 1.17583e-08, 1.179835e-08, 1.182618e-08, 
    1.181397e-08, 1.187738e-08, 1.189232e-08, 1.195305e-08, 1.192166e-08, 
    1.210855e-08, 1.202587e-08, 1.22553e-08, 1.219119e-08, 1.175873e-08, 
    1.177904e-08, 1.18497e-08, 1.181608e-08, 1.191223e-08, 1.19359e-08, 
    1.195514e-08, 1.197974e-08, 1.198239e-08, 1.199696e-08, 1.197308e-08, 
    1.199602e-08, 1.190925e-08, 1.194803e-08, 1.184162e-08, 1.186752e-08, 
    1.185561e-08, 1.184254e-08, 1.188287e-08, 1.192585e-08, 1.192676e-08, 
    1.194054e-08, 1.197937e-08, 1.191262e-08, 1.211923e-08, 1.199164e-08, 
    1.180118e-08, 1.184029e-08, 1.184587e-08, 1.183072e-08, 1.193353e-08, 
    1.189628e-08, 1.199661e-08, 1.196949e-08, 1.201392e-08, 1.199184e-08, 
    1.198859e-08, 1.196024e-08, 1.194259e-08, 1.189799e-08, 1.18617e-08, 
    1.183292e-08, 1.183961e-08, 1.187122e-08, 1.192847e-08, 1.198263e-08, 
    1.197077e-08, 1.201054e-08, 1.190526e-08, 1.194941e-08, 1.193235e-08, 
    1.197684e-08, 1.187935e-08, 1.196237e-08, 1.185813e-08, 1.186727e-08, 
    1.189554e-08, 1.19524e-08, 1.196498e-08, 1.197842e-08, 1.197013e-08, 
    1.192993e-08, 1.192334e-08, 1.189485e-08, 1.188699e-08, 1.186528e-08, 
    1.184731e-08, 1.186373e-08, 1.188097e-08, 1.192994e-08, 1.197407e-08, 
    1.202219e-08, 1.203396e-08, 1.209018e-08, 1.204442e-08, 1.211994e-08, 
    1.205574e-08, 1.216687e-08, 1.196718e-08, 1.205384e-08, 1.189682e-08, 
    1.191374e-08, 1.194434e-08, 1.201451e-08, 1.197663e-08, 1.202093e-08, 
    1.192308e-08, 1.187231e-08, 1.185918e-08, 1.183467e-08, 1.185974e-08, 
    1.18577e-08, 1.188168e-08, 1.187398e-08, 1.193157e-08, 1.190063e-08, 
    1.198851e-08, 1.202058e-08, 1.211115e-08, 1.216666e-08, 1.222317e-08, 
    1.224812e-08, 1.225572e-08, 1.225889e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382061e-10, 1.388139e-10, 1.386958e-10, 1.391861e-10, 1.389141e-10, 
    1.392351e-10, 1.383293e-10, 1.388381e-10, 1.385133e-10, 1.382608e-10, 
    1.401376e-10, 1.39208e-10, 1.411032e-10, 1.405103e-10, 1.419996e-10, 
    1.410109e-10, 1.42199e-10, 1.419711e-10, 1.42657e-10, 1.424605e-10, 
    1.433378e-10, 1.427476e-10, 1.437925e-10, 1.431968e-10, 1.4329e-10, 
    1.427282e-10, 1.39395e-10, 1.400219e-10, 1.393579e-10, 1.394473e-10, 
    1.394072e-10, 1.389197e-10, 1.386741e-10, 1.381596e-10, 1.38253e-10, 
    1.386309e-10, 1.394875e-10, 1.391967e-10, 1.399295e-10, 1.39913e-10, 
    1.407288e-10, 1.40361e-10, 1.417322e-10, 1.413425e-10, 1.424687e-10, 
    1.421854e-10, 1.424554e-10, 1.423735e-10, 1.424564e-10, 1.42041e-10, 
    1.42219e-10, 1.418535e-10, 1.404298e-10, 1.408483e-10, 1.396004e-10, 
    1.3885e-10, 1.383516e-10, 1.379979e-10, 1.380479e-10, 1.381433e-10, 
    1.386331e-10, 1.390936e-10, 1.394445e-10, 1.396793e-10, 1.399106e-10, 
    1.406107e-10, 1.409813e-10, 1.41811e-10, 1.416613e-10, 1.419149e-10, 
    1.421573e-10, 1.425641e-10, 1.424972e-10, 1.426764e-10, 1.419082e-10, 
    1.424188e-10, 1.41576e-10, 1.418065e-10, 1.399735e-10, 1.392751e-10, 
    1.389783e-10, 1.387185e-10, 1.380864e-10, 1.385229e-10, 1.383508e-10, 
    1.387602e-10, 1.390203e-10, 1.388917e-10, 1.396857e-10, 1.39377e-10, 
    1.410033e-10, 1.403028e-10, 1.42129e-10, 1.41692e-10, 1.422337e-10, 
    1.419573e-10, 1.42431e-10, 1.420047e-10, 1.427431e-10, 1.429039e-10, 
    1.42794e-10, 1.432161e-10, 1.41981e-10, 1.424554e-10, 1.388881e-10, 
    1.389091e-10, 1.390068e-10, 1.385771e-10, 1.385508e-10, 1.38157e-10, 
    1.385074e-10, 1.386566e-10, 1.390354e-10, 1.392595e-10, 1.394724e-10, 
    1.399407e-10, 1.404637e-10, 1.41195e-10, 1.417203e-10, 1.420725e-10, 
    1.418565e-10, 1.420472e-10, 1.418341e-10, 1.417342e-10, 1.428437e-10, 
    1.422207e-10, 1.431554e-10, 1.431037e-10, 1.426807e-10, 1.431095e-10, 
    1.389238e-10, 1.38803e-10, 1.383838e-10, 1.387119e-10, 1.381141e-10, 
    1.384488e-10, 1.386411e-10, 1.393835e-10, 1.395465e-10, 1.396978e-10, 
    1.399965e-10, 1.403798e-10, 1.410522e-10, 1.416373e-10, 1.421714e-10, 
    1.421322e-10, 1.42146e-10, 1.422653e-10, 1.419698e-10, 1.423138e-10, 
    1.423716e-10, 1.422206e-10, 1.430968e-10, 1.428465e-10, 1.431026e-10, 
    1.429396e-10, 1.388423e-10, 1.390455e-10, 1.389357e-10, 1.391421e-10, 
    1.389967e-10, 1.396434e-10, 1.398373e-10, 1.407446e-10, 1.403722e-10, 
    1.409649e-10, 1.404324e-10, 1.405268e-10, 1.409842e-10, 1.404612e-10, 
    1.41605e-10, 1.408296e-10, 1.4227e-10, 1.414956e-10, 1.423185e-10, 
    1.421691e-10, 1.424165e-10, 1.426381e-10, 1.429168e-10, 1.434312e-10, 
    1.433121e-10, 1.437422e-10, 1.393483e-10, 1.396119e-10, 1.395887e-10, 
    1.398644e-10, 1.400684e-10, 1.405105e-10, 1.412195e-10, 1.409528e-10, 
    1.414423e-10, 1.415405e-10, 1.407969e-10, 1.412535e-10, 1.397882e-10, 
    1.40025e-10, 1.39884e-10, 1.393691e-10, 1.410143e-10, 1.4017e-10, 
    1.41729e-10, 1.412716e-10, 1.426065e-10, 1.419426e-10, 1.432465e-10, 
    1.438039e-10, 1.443285e-10, 1.449416e-10, 1.397557e-10, 1.395766e-10, 
    1.398972e-10, 1.403408e-10, 1.407524e-10, 1.412995e-10, 1.413555e-10, 
    1.41458e-10, 1.417235e-10, 1.419468e-10, 1.414904e-10, 1.420027e-10, 
    1.400799e-10, 1.410876e-10, 1.395089e-10, 1.399843e-10, 1.403147e-10, 
    1.401698e-10, 1.409224e-10, 1.410997e-10, 1.418206e-10, 1.414479e-10, 
    1.436664e-10, 1.426849e-10, 1.454084e-10, 1.446473e-10, 1.395141e-10, 
    1.397551e-10, 1.405939e-10, 1.401948e-10, 1.413361e-10, 1.41617e-10, 
    1.418454e-10, 1.421373e-10, 1.421688e-10, 1.423418e-10, 1.420583e-10, 
    1.423306e-10, 1.413007e-10, 1.417609e-10, 1.40498e-10, 1.408054e-10, 
    1.406639e-10, 1.405088e-10, 1.409876e-10, 1.414976e-10, 1.415085e-10, 
    1.416721e-10, 1.42133e-10, 1.413407e-10, 1.437931e-10, 1.422786e-10, 
    1.400179e-10, 1.404821e-10, 1.405484e-10, 1.403686e-10, 1.415888e-10, 
    1.411467e-10, 1.423376e-10, 1.420157e-10, 1.425431e-10, 1.42281e-10, 
    1.422425e-10, 1.419059e-10, 1.416963e-10, 1.41167e-10, 1.407362e-10, 
    1.403946e-10, 1.404741e-10, 1.408493e-10, 1.415288e-10, 1.421717e-10, 
    1.420309e-10, 1.42503e-10, 1.412533e-10, 1.417773e-10, 1.415748e-10, 
    1.421029e-10, 1.409458e-10, 1.419312e-10, 1.406939e-10, 1.408024e-10, 
    1.411379e-10, 1.418129e-10, 1.419622e-10, 1.421216e-10, 1.420232e-10, 
    1.415461e-10, 1.414679e-10, 1.411297e-10, 1.410364e-10, 1.407787e-10, 
    1.405654e-10, 1.407603e-10, 1.40965e-10, 1.415463e-10, 1.420701e-10, 
    1.426412e-10, 1.42781e-10, 1.434483e-10, 1.429051e-10, 1.438015e-10, 
    1.430394e-10, 1.443586e-10, 1.419882e-10, 1.43017e-10, 1.411532e-10, 
    1.41354e-10, 1.417171e-10, 1.425501e-10, 1.421004e-10, 1.426263e-10, 
    1.414648e-10, 1.408622e-10, 1.407063e-10, 1.404154e-10, 1.40713e-10, 
    1.406888e-10, 1.409735e-10, 1.40882e-10, 1.415656e-10, 1.411984e-10, 
    1.422415e-10, 1.426222e-10, 1.436972e-10, 1.443562e-10, 1.45027e-10, 
    1.453231e-10, 1.454133e-10, 1.45451e-10 ;

 SOIL1N_vr =
  2.497419, 2.497412, 2.497414, 2.497408, 2.497411, 2.497408, 2.497418, 
    2.497412, 2.497416, 2.497418, 2.497398, 2.497408, 2.497387, 2.497393, 
    2.497377, 2.497388, 2.497375, 2.497377, 2.49737, 2.497372, 2.497362, 
    2.497369, 2.497357, 2.497364, 2.497363, 2.497369, 2.497406, 2.497399, 
    2.497406, 2.497405, 2.497406, 2.497411, 2.497414, 2.49742, 2.497418, 
    2.497414, 2.497405, 2.497408, 2.4974, 2.4974, 2.497391, 2.497395, 
    2.49738, 2.497384, 2.497372, 2.497375, 2.497372, 2.497373, 2.497372, 
    2.497376, 2.497375, 2.497379, 2.497394, 2.49739, 2.497404, 2.497412, 
    2.497417, 2.497421, 2.497421, 2.49742, 2.497414, 2.497409, 2.497405, 
    2.497403, 2.4974, 2.497392, 2.497388, 2.497379, 2.497381, 2.497378, 
    2.497375, 2.497371, 2.497371, 2.49737, 2.497378, 2.497372, 2.497382, 
    2.497379, 2.497399, 2.497407, 2.49741, 2.497413, 2.49742, 2.497416, 
    2.497417, 2.497413, 2.49741, 2.497411, 2.497403, 2.497406, 2.497388, 
    2.497396, 2.497375, 2.49738, 2.497374, 2.497377, 2.497372, 2.497377, 
    2.497369, 2.497367, 2.497368, 2.497364, 2.497377, 2.497372, 2.497411, 
    2.497411, 2.49741, 2.497415, 2.497415, 2.49742, 2.497416, 2.497414, 
    2.49741, 2.497407, 2.497405, 2.4974, 2.497394, 2.497386, 2.49738, 
    2.497376, 2.497379, 2.497376, 2.497379, 2.49738, 2.497368, 2.497375, 
    2.497364, 2.497365, 2.49737, 2.497365, 2.497411, 2.497412, 2.497417, 
    2.497413, 2.49742, 2.497416, 2.497414, 2.497406, 2.497404, 2.497402, 
    2.497399, 2.497395, 2.497387, 2.497381, 2.497375, 2.497375, 2.497375, 
    2.497374, 2.497377, 2.497374, 2.497373, 2.497375, 2.497365, 2.497368, 
    2.497365, 2.497367, 2.497412, 2.49741, 2.497411, 2.497409, 2.49741, 
    2.497403, 2.497401, 2.497391, 2.497395, 2.497388, 2.497394, 2.497393, 
    2.497388, 2.497394, 2.497381, 2.49739, 2.497374, 2.497383, 2.497374, 
    2.497375, 2.497372, 2.49737, 2.497367, 2.497361, 2.497363, 2.497358, 
    2.497406, 2.497403, 2.497404, 2.497401, 2.497398, 2.497393, 2.497386, 
    2.497389, 2.497383, 2.497382, 2.49739, 2.497385, 2.497401, 2.497399, 
    2.4974, 2.497406, 2.497388, 2.497397, 2.49738, 2.497385, 2.49737, 
    2.497378, 2.497363, 2.497357, 2.497351, 2.497345, 2.497402, 2.497404, 
    2.4974, 2.497395, 2.497391, 2.497385, 2.497384, 2.497383, 2.49738, 
    2.497378, 2.497383, 2.497377, 2.497398, 2.497387, 2.497405, 2.497399, 
    2.497396, 2.497397, 2.497389, 2.497387, 2.497379, 2.497383, 2.497359, 
    2.49737, 2.497339, 2.497348, 2.497405, 2.497402, 2.497392, 2.497397, 
    2.497384, 2.497381, 2.497379, 2.497375, 2.497375, 2.497373, 2.497376, 
    2.497373, 2.497385, 2.49738, 2.497394, 2.49739, 2.497392, 2.497393, 
    2.497388, 2.497382, 2.497382, 2.49738, 2.497375, 2.497384, 2.497357, 
    2.497374, 2.497399, 2.497394, 2.497393, 2.497395, 2.497381, 2.497386, 
    2.497373, 2.497377, 2.497371, 2.497374, 2.497374, 2.497378, 2.49738, 
    2.497386, 2.497391, 2.497395, 2.497394, 2.49739, 2.497382, 2.497375, 
    2.497377, 2.497371, 2.497385, 2.49738, 2.497382, 2.497376, 2.497389, 
    2.497378, 2.497391, 2.49739, 2.497386, 2.497379, 2.497377, 2.497376, 
    2.497377, 2.497382, 2.497383, 2.497387, 2.497388, 2.497391, 2.497393, 
    2.497391, 2.497388, 2.497382, 2.497376, 2.49737, 2.497368, 2.497361, 
    2.497367, 2.497357, 2.497365, 2.497351, 2.497377, 2.497366, 2.497386, 
    2.497384, 2.49738, 2.497371, 2.497376, 2.49737, 2.497383, 2.49739, 
    2.497391, 2.497395, 2.497391, 2.497391, 2.497388, 2.497389, 2.497382, 
    2.497386, 2.497374, 2.49737, 2.497358, 2.497351, 2.497344, 2.49734, 
    2.497339, 2.497339,
  2.497626, 2.497617, 2.497619, 2.497612, 2.497616, 2.497611, 2.497624, 
    2.497617, 2.497622, 2.497625, 2.497598, 2.497611, 2.497584, 2.497592, 
    2.497571, 2.497585, 2.497568, 2.497571, 2.497561, 2.497564, 2.497551, 
    2.49756, 2.497545, 2.497553, 2.497552, 2.49756, 2.497609, 2.497599, 
    2.497609, 2.497608, 2.497608, 2.497616, 2.497619, 2.497627, 2.497625, 
    2.49762, 2.497607, 2.497612, 2.497601, 2.497601, 2.497589, 2.497595, 
    2.497575, 2.49758, 2.497564, 2.497568, 2.497564, 2.497565, 2.497564, 
    2.49757, 2.497567, 2.497573, 2.497593, 2.497587, 2.497606, 2.497617, 
    2.497624, 2.497629, 2.497628, 2.497627, 2.49762, 2.497613, 2.497608, 
    2.497604, 2.497601, 2.497591, 2.497586, 2.497573, 2.497576, 2.497572, 
    2.497568, 2.497562, 2.497563, 2.497561, 2.497572, 2.497565, 2.497577, 
    2.497573, 2.4976, 2.49761, 2.497615, 2.497618, 2.497628, 2.497621, 
    2.497624, 2.497618, 2.497614, 2.497616, 2.497604, 2.497609, 2.497585, 
    2.497595, 2.497569, 2.497575, 2.497567, 2.497571, 2.497564, 2.497571, 
    2.49756, 2.497558, 2.497559, 2.497553, 2.497571, 2.497564, 2.497616, 
    2.497616, 2.497614, 2.497621, 2.497621, 2.497627, 2.497622, 2.497619, 
    2.497614, 2.497611, 2.497607, 2.497601, 2.497593, 2.497582, 2.497575, 
    2.49757, 2.497573, 2.49757, 2.497573, 2.497575, 2.497558, 2.497567, 
    2.497554, 2.497555, 2.497561, 2.497555, 2.497615, 2.497617, 2.497623, 
    2.497618, 2.497627, 2.497622, 2.49762, 2.497609, 2.497606, 2.497604, 
    2.4976, 2.497594, 2.497584, 2.497576, 2.497568, 2.497569, 2.497569, 
    2.497567, 2.497571, 2.497566, 2.497565, 2.497567, 2.497555, 2.497558, 
    2.497555, 2.497557, 2.497617, 2.497614, 2.497615, 2.497612, 2.497614, 
    2.497605, 2.497602, 2.497589, 2.497594, 2.497586, 2.497593, 2.497592, 
    2.497585, 2.497593, 2.497576, 2.497588, 2.497567, 2.497578, 2.497566, 
    2.497568, 2.497565, 2.497561, 2.497557, 2.49755, 2.497552, 2.497545, 
    2.497609, 2.497605, 2.497606, 2.497602, 2.497599, 2.497592, 2.497582, 
    2.497586, 2.497579, 2.497577, 2.497588, 2.497581, 2.497603, 2.497599, 
    2.497602, 2.497609, 2.497585, 2.497597, 2.497575, 2.497581, 2.497562, 
    2.497571, 2.497553, 2.497545, 2.497537, 2.497528, 2.497603, 2.497606, 
    2.497601, 2.497595, 2.497589, 2.497581, 2.49758, 2.497579, 2.497575, 
    2.497571, 2.497578, 2.497571, 2.497599, 2.497584, 2.497607, 2.4976, 
    2.497595, 2.497597, 2.497586, 2.497584, 2.497573, 2.497579, 2.497546, 
    2.497561, 2.497521, 2.497532, 2.497607, 2.497603, 2.497591, 2.497597, 
    2.49758, 2.497576, 2.497573, 2.497569, 2.497568, 2.497566, 2.49757, 
    2.497566, 2.497581, 2.497574, 2.497592, 2.497588, 2.49759, 2.497592, 
    2.497585, 2.497578, 2.497578, 2.497576, 2.497569, 2.49758, 2.497545, 
    2.497567, 2.497599, 2.497593, 2.497592, 2.497594, 2.497577, 2.497583, 
    2.497566, 2.497571, 2.497563, 2.497566, 2.497567, 2.497572, 2.497575, 
    2.497583, 2.497589, 2.497594, 2.497593, 2.497587, 2.497577, 2.497568, 
    2.49757, 2.497563, 2.497581, 2.497574, 2.497577, 2.497569, 2.497586, 
    2.497572, 2.49759, 2.497588, 2.497583, 2.497573, 2.497571, 2.497569, 
    2.49757, 2.497577, 2.497578, 2.497583, 2.497585, 2.497588, 2.497591, 
    2.497589, 2.497586, 2.497577, 2.49757, 2.497561, 2.497559, 2.49755, 
    2.497558, 2.497545, 2.497555, 2.497536, 2.497571, 2.497556, 2.497583, 
    2.49758, 2.497575, 2.497563, 2.497569, 2.497561, 2.497578, 2.497587, 
    2.497589, 2.497594, 2.497589, 2.49759, 2.497586, 2.497587, 2.497577, 
    2.497582, 2.497567, 2.497562, 2.497546, 2.497536, 2.497527, 2.497523, 
    2.497521, 2.497521,
  2.497841, 2.497832, 2.497833, 2.497826, 2.49783, 2.497825, 2.497839, 
    2.497831, 2.497836, 2.49784, 2.497811, 2.497825, 2.497796, 2.497805, 
    2.497782, 2.497797, 2.497779, 2.497782, 2.497772, 2.497775, 2.497761, 
    2.49777, 2.497754, 2.497763, 2.497762, 2.497771, 2.497823, 2.497813, 
    2.497823, 2.497822, 2.497822, 2.49783, 2.497834, 2.497842, 2.49784, 
    2.497834, 2.497821, 2.497826, 2.497814, 2.497814, 2.497802, 2.497808, 
    2.497786, 2.497792, 2.497775, 2.497779, 2.497775, 2.497776, 2.497775, 
    2.497781, 2.497779, 2.497784, 2.497806, 2.4978, 2.497819, 2.497831, 
    2.497839, 2.497844, 2.497844, 2.497842, 2.497834, 2.497827, 2.497822, 
    2.497818, 2.497814, 2.497804, 2.497798, 2.497785, 2.497787, 2.497783, 
    2.49778, 2.497773, 2.497774, 2.497772, 2.497783, 2.497776, 2.497789, 
    2.497785, 2.497813, 2.497824, 2.497829, 2.497833, 2.497843, 2.497836, 
    2.497839, 2.497832, 2.497828, 2.49783, 2.497818, 2.497823, 2.497797, 
    2.497808, 2.49778, 2.497787, 2.497778, 2.497783, 2.497775, 2.497782, 
    2.497771, 2.497768, 2.49777, 2.497763, 2.497782, 2.497775, 2.49783, 
    2.49783, 2.497828, 2.497835, 2.497836, 2.497842, 2.497836, 2.497834, 
    2.497828, 2.497825, 2.497821, 2.497814, 2.497806, 2.497794, 2.497786, 
    2.497781, 2.497784, 2.497781, 2.497785, 2.497786, 2.497769, 2.497779, 
    2.497764, 2.497765, 2.497772, 2.497765, 2.49783, 2.497832, 2.497838, 
    2.497833, 2.497843, 2.497837, 2.497834, 2.497823, 2.49782, 2.497818, 
    2.497813, 2.497807, 2.497797, 2.497788, 2.497779, 2.49778, 2.49778, 
    2.497778, 2.497782, 2.497777, 2.497776, 2.497779, 2.497765, 2.497769, 
    2.497765, 2.497767, 2.497831, 2.497828, 2.49783, 2.497826, 2.497829, 
    2.497819, 2.497816, 2.497802, 2.497807, 2.497798, 2.497806, 2.497805, 
    2.497798, 2.497806, 2.497788, 2.4978, 2.497778, 2.49779, 2.497777, 
    2.497779, 2.497776, 2.497772, 2.497768, 2.49776, 2.497762, 2.497755, 
    2.497823, 2.497819, 2.497819, 2.497815, 2.497812, 2.497805, 2.497794, 
    2.497798, 2.497791, 2.497789, 2.497801, 2.497794, 2.497816, 2.497813, 
    2.497815, 2.497823, 2.497797, 2.49781, 2.497786, 2.497793, 2.497773, 
    2.497783, 2.497763, 2.497754, 2.497746, 2.497736, 2.497817, 2.49782, 
    2.497815, 2.497808, 2.497801, 2.497793, 2.497792, 2.49779, 2.497786, 
    2.497783, 2.49779, 2.497782, 2.497812, 2.497796, 2.497821, 2.497813, 
    2.497808, 2.49781, 2.497799, 2.497796, 2.497785, 2.497791, 2.497756, 
    2.497771, 2.497729, 2.497741, 2.497821, 2.497817, 2.497804, 2.49781, 
    2.497792, 2.497788, 2.497784, 2.49778, 2.497779, 2.497777, 2.497781, 
    2.497777, 2.497793, 2.497786, 2.497805, 2.497801, 2.497803, 2.497805, 
    2.497798, 2.49779, 2.49779, 2.497787, 2.49778, 2.497792, 2.497754, 
    2.497778, 2.497813, 2.497806, 2.497805, 2.497807, 2.497788, 2.497795, 
    2.497777, 2.497782, 2.497774, 2.497778, 2.497778, 2.497783, 2.497787, 
    2.497795, 2.497802, 2.497807, 2.497806, 2.4978, 2.497789, 2.497779, 
    2.497782, 2.497774, 2.497794, 2.497786, 2.497789, 2.49778, 2.497798, 
    2.497783, 2.497802, 2.497801, 2.497795, 2.497785, 2.497783, 2.49778, 
    2.497782, 2.497789, 2.49779, 2.497796, 2.497797, 2.497801, 2.497804, 
    2.497801, 2.497798, 2.497789, 2.497781, 2.497772, 2.49777, 2.49776, 
    2.497768, 2.497754, 2.497766, 2.497746, 2.497782, 2.497766, 2.497795, 
    2.497792, 2.497786, 2.497773, 2.497781, 2.497772, 2.49779, 2.4978, 
    2.497802, 2.497807, 2.497802, 2.497802, 2.497798, 2.497799, 2.497789, 
    2.497794, 2.497778, 2.497772, 2.497756, 2.497746, 2.497735, 2.49773, 
    2.497729, 2.497729,
  2.498013, 2.498003, 2.498005, 2.497998, 2.498002, 2.497997, 2.498011, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.49797, 2.497951, 2.497955, 2.497944, 2.497947, 2.497934, 
    2.497943, 2.497927, 2.497936, 2.497934, 2.497943, 2.497994, 2.497985, 
    2.497995, 2.497994, 2.497994, 2.498002, 2.498006, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497998, 2.497986, 2.497987, 2.497974, 2.49798, 
    2.497958, 2.497964, 2.497947, 2.497952, 2.497947, 2.497949, 2.497947, 
    2.497954, 2.497951, 2.497957, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.498011, 2.498016, 2.498015, 2.498014, 2.498006, 2.497999, 2.497994, 
    2.49799, 2.497987, 2.497976, 2.49797, 2.497957, 2.49796, 2.497956, 
    2.497952, 2.497946, 2.497947, 2.497944, 2.497956, 2.497948, 2.497961, 
    2.497957, 2.497986, 2.497996, 2.498001, 2.498005, 2.498015, 2.498008, 
    2.498011, 2.498004, 2.498, 2.498002, 2.49799, 2.497995, 2.49797, 2.49798, 
    2.497952, 2.497959, 2.497951, 2.497955, 2.497948, 2.497954, 2.497943, 
    2.49794, 2.497942, 2.497936, 2.497955, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498008, 2.498013, 2.498008, 2.498006, 2.498, 2.497997, 
    2.497993, 2.497986, 2.497978, 2.497967, 2.497959, 2.497953, 2.497957, 
    2.497954, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497944, 2.497937, 2.498002, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497995, 2.497992, 2.49799, 2.497985, 2.497979, 
    2.497969, 2.49796, 2.497952, 2.497952, 2.497952, 2.49795, 2.497955, 
    2.497949, 2.497949, 2.497951, 2.497937, 2.497941, 2.497937, 2.49794, 
    2.498003, 2.498, 2.498002, 2.497998, 2.498001, 2.497991, 2.497988, 
    2.497974, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497978, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497952, 2.497948, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497992, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497963, 
    2.497961, 2.497973, 2.497966, 2.497988, 2.497985, 2.497987, 2.497995, 
    2.497969, 2.497983, 2.497958, 2.497966, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497989, 2.497992, 2.497987, 2.49798, 
    2.497973, 2.497965, 2.497964, 2.497963, 2.497959, 2.497955, 2.497962, 
    2.497954, 2.497984, 2.497968, 2.497993, 2.497985, 2.49798, 2.497983, 
    2.497971, 2.497968, 2.497957, 2.497963, 2.497929, 2.497944, 2.497902, 
    2.497914, 2.497993, 2.497989, 2.497976, 2.497982, 2.497965, 2.49796, 
    2.497957, 2.497952, 2.497952, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497958, 2.497977, 2.497973, 2.497975, 2.497977, 2.49797, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497927, 2.49795, 2.497985, 
    2.497978, 2.497977, 2.497979, 2.497961, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.497951, 2.497956, 2.497959, 2.497967, 2.497974, 
    2.497979, 2.497978, 2.497972, 2.497962, 2.497952, 2.497954, 2.497947, 
    2.497966, 2.497958, 2.497961, 2.497953, 2.497971, 2.497955, 2.497974, 
    2.497973, 2.497967, 2.497957, 2.497955, 2.497952, 2.497954, 2.497961, 
    2.497962, 2.497968, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497932, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497939, 2.497967, 2.497964, 2.497959, 
    2.497946, 2.497953, 2.497945, 2.497962, 2.497972, 2.497974, 2.497979, 
    2.497974, 2.497974, 2.49797, 2.497972, 2.497961, 2.497967, 2.497951, 
    2.497945, 2.497928, 2.497918, 2.497908, 2.497903, 2.497902, 2.497901,
  2.498213, 2.498205, 2.498207, 2.4982, 2.498204, 2.498199, 2.498212, 
    2.498205, 2.498209, 2.498213, 2.498187, 2.498199, 2.498174, 2.498182, 
    2.498161, 2.498175, 2.498159, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498144, 2.498151, 2.498197, 2.498188, 
    2.498198, 2.498196, 2.498197, 2.498204, 2.498207, 2.498214, 2.498213, 
    2.498207, 2.498196, 2.4982, 2.49819, 2.49819, 2.498179, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498163, 
    2.498159, 2.498154, 2.498154, 2.498152, 2.498163, 2.498156, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498206, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498185, 2.49816, 2.498166, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498145, 2.498162, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498209, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498164, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498204, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498189, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498184, 2.498175, 2.498183, 2.498182, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498156, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.498191, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498172, 2.498192, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498137, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498169, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498174, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498115, 2.498125, 2.498195, 2.498192, 2.498181, 2.498186, 
    2.49817, 2.498167, 2.498163, 2.498159, 2.498159, 2.498157, 2.498161, 
    2.498157, 2.498171, 2.498165, 2.498182, 2.498178, 2.49818, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498158, 2.498188, 2.498182, 2.498181, 2.498184, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498158, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498179, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498172, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.49816, 
    2.498161, 2.498168, 2.498169, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498168, 2.49816, 2.498152, 2.498151, 2.498142, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498162, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498153, 2.498169, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.138676e-08, 6.165671e-08, 6.160423e-08, 6.182197e-08, 6.170119e-08, 
    6.184376e-08, 6.144149e-08, 6.166744e-08, 6.15232e-08, 6.141106e-08, 
    6.224452e-08, 6.183168e-08, 6.267332e-08, 6.241004e-08, 6.30714e-08, 
    6.263235e-08, 6.315993e-08, 6.305873e-08, 6.33633e-08, 6.327605e-08, 
    6.366562e-08, 6.340358e-08, 6.386756e-08, 6.360304e-08, 6.364442e-08, 
    6.339493e-08, 6.191476e-08, 6.219313e-08, 6.189827e-08, 6.193796e-08, 
    6.192015e-08, 6.170368e-08, 6.15946e-08, 6.136612e-08, 6.14076e-08, 
    6.157541e-08, 6.195581e-08, 6.182668e-08, 6.215211e-08, 6.214476e-08, 
    6.250706e-08, 6.234371e-08, 6.295264e-08, 6.277958e-08, 6.327969e-08, 
    6.315392e-08, 6.327378e-08, 6.323744e-08, 6.327426e-08, 6.308979e-08, 
    6.316883e-08, 6.300651e-08, 6.23743e-08, 6.256011e-08, 6.200595e-08, 
    6.167274e-08, 6.14514e-08, 6.129434e-08, 6.131655e-08, 6.135888e-08, 
    6.157639e-08, 6.17809e-08, 6.193674e-08, 6.204099e-08, 6.214371e-08, 
    6.245464e-08, 6.261919e-08, 6.298765e-08, 6.292114e-08, 6.30338e-08, 
    6.314141e-08, 6.332208e-08, 6.329234e-08, 6.337194e-08, 6.303082e-08, 
    6.325753e-08, 6.288327e-08, 6.298563e-08, 6.217166e-08, 6.186151e-08, 
    6.172971e-08, 6.161432e-08, 6.133362e-08, 6.152747e-08, 6.145105e-08, 
    6.163285e-08, 6.174837e-08, 6.169123e-08, 6.204384e-08, 6.190675e-08, 
    6.262894e-08, 6.231787e-08, 6.312885e-08, 6.293479e-08, 6.317536e-08, 
    6.30526e-08, 6.326295e-08, 6.307364e-08, 6.340156e-08, 6.347297e-08, 
    6.342418e-08, 6.361162e-08, 6.306315e-08, 6.327378e-08, 6.168963e-08, 
    6.169895e-08, 6.174236e-08, 6.155154e-08, 6.153986e-08, 6.136499e-08, 
    6.152059e-08, 6.158686e-08, 6.175506e-08, 6.185456e-08, 6.194914e-08, 
    6.215708e-08, 6.238933e-08, 6.271407e-08, 6.294737e-08, 6.310376e-08, 
    6.300786e-08, 6.309252e-08, 6.299788e-08, 6.295353e-08, 6.344622e-08, 
    6.316957e-08, 6.358466e-08, 6.356169e-08, 6.337384e-08, 6.356428e-08, 
    6.170549e-08, 6.165187e-08, 6.146571e-08, 6.16114e-08, 6.134594e-08, 
    6.149453e-08, 6.157997e-08, 6.190962e-08, 6.198205e-08, 6.204921e-08, 
    6.218185e-08, 6.235207e-08, 6.265068e-08, 6.291049e-08, 6.314767e-08, 
    6.313029e-08, 6.31364e-08, 6.318939e-08, 6.305815e-08, 6.321093e-08, 
    6.323658e-08, 6.316953e-08, 6.355862e-08, 6.344746e-08, 6.35612e-08, 
    6.348883e-08, 6.16693e-08, 6.175953e-08, 6.171077e-08, 6.180245e-08, 
    6.173786e-08, 6.202507e-08, 6.211118e-08, 6.251408e-08, 6.234873e-08, 
    6.261189e-08, 6.237546e-08, 6.241735e-08, 6.262048e-08, 6.238822e-08, 
    6.289618e-08, 6.255181e-08, 6.319145e-08, 6.284758e-08, 6.321299e-08, 
    6.314664e-08, 6.325651e-08, 6.33549e-08, 6.347869e-08, 6.370711e-08, 
    6.365422e-08, 6.384523e-08, 6.189403e-08, 6.201106e-08, 6.200075e-08, 
    6.212322e-08, 6.221379e-08, 6.241009e-08, 6.272494e-08, 6.260655e-08, 
    6.28239e-08, 6.286754e-08, 6.253732e-08, 6.274008e-08, 6.208938e-08, 
    6.219452e-08, 6.213192e-08, 6.190326e-08, 6.263384e-08, 6.225891e-08, 
    6.295123e-08, 6.274812e-08, 6.334088e-08, 6.304609e-08, 6.36251e-08, 
    6.387263e-08, 6.410557e-08, 6.437782e-08, 6.207492e-08, 6.199541e-08, 
    6.213779e-08, 6.233478e-08, 6.251754e-08, 6.276051e-08, 6.278537e-08, 
    6.283089e-08, 6.294879e-08, 6.304793e-08, 6.284529e-08, 6.307278e-08, 
    6.221891e-08, 6.266638e-08, 6.196535e-08, 6.217645e-08, 6.232316e-08, 
    6.22588e-08, 6.259302e-08, 6.267179e-08, 6.299189e-08, 6.282641e-08, 
    6.381155e-08, 6.33757e-08, 6.458509e-08, 6.424712e-08, 6.196763e-08, 
    6.207465e-08, 6.244714e-08, 6.22699e-08, 6.277673e-08, 6.290148e-08, 
    6.300289e-08, 6.313254e-08, 6.314653e-08, 6.322334e-08, 6.309747e-08, 
    6.321837e-08, 6.276103e-08, 6.296541e-08, 6.240455e-08, 6.254106e-08, 
    6.247826e-08, 6.240938e-08, 6.262198e-08, 6.284848e-08, 6.285331e-08, 
    6.292594e-08, 6.313062e-08, 6.277878e-08, 6.386782e-08, 6.319527e-08, 
    6.219135e-08, 6.239751e-08, 6.242694e-08, 6.234709e-08, 6.288898e-08, 
    6.269264e-08, 6.322147e-08, 6.307854e-08, 6.331273e-08, 6.319635e-08, 
    6.317924e-08, 6.302977e-08, 6.293672e-08, 6.270164e-08, 6.251035e-08, 
    6.235867e-08, 6.239394e-08, 6.256057e-08, 6.286233e-08, 6.31478e-08, 
    6.308527e-08, 6.329493e-08, 6.273998e-08, 6.297268e-08, 6.288275e-08, 
    6.311726e-08, 6.260341e-08, 6.3041e-08, 6.249155e-08, 6.253973e-08, 
    6.268873e-08, 6.298848e-08, 6.305478e-08, 6.312558e-08, 6.308189e-08, 
    6.286999e-08, 6.283527e-08, 6.268511e-08, 6.264366e-08, 6.252924e-08, 
    6.243451e-08, 6.252106e-08, 6.261195e-08, 6.287008e-08, 6.31027e-08, 
    6.335631e-08, 6.341837e-08, 6.371471e-08, 6.347349e-08, 6.387156e-08, 
    6.353314e-08, 6.411896e-08, 6.306635e-08, 6.352317e-08, 6.269551e-08, 
    6.278468e-08, 6.294596e-08, 6.331585e-08, 6.311615e-08, 6.33497e-08, 
    6.283391e-08, 6.256631e-08, 6.249707e-08, 6.23679e-08, 6.250002e-08, 
    6.248928e-08, 6.261571e-08, 6.257508e-08, 6.287865e-08, 6.271559e-08, 
    6.317881e-08, 6.334785e-08, 6.382522e-08, 6.411786e-08, 6.441574e-08, 
    6.454725e-08, 6.458728e-08, 6.460402e-08 ;

 SOIL1_HR_S3 =
  7.284729e-10, 7.316777e-10, 7.310547e-10, 7.336395e-10, 7.322056e-10, 
    7.338982e-10, 7.291227e-10, 7.318049e-10, 7.300926e-10, 7.287614e-10, 
    7.38656e-10, 7.337548e-10, 7.437466e-10, 7.406208e-10, 7.484727e-10, 
    7.432602e-10, 7.495237e-10, 7.483222e-10, 7.519381e-10, 7.509022e-10, 
    7.555275e-10, 7.524162e-10, 7.57925e-10, 7.547844e-10, 7.552758e-10, 
    7.523137e-10, 7.34741e-10, 7.380458e-10, 7.345453e-10, 7.350165e-10, 
    7.348051e-10, 7.322353e-10, 7.309403e-10, 7.28228e-10, 7.287204e-10, 
    7.307125e-10, 7.352284e-10, 7.336954e-10, 7.375588e-10, 7.374716e-10, 
    7.417728e-10, 7.398335e-10, 7.470627e-10, 7.45008e-10, 7.509455e-10, 
    7.494523e-10, 7.508754e-10, 7.504438e-10, 7.50881e-10, 7.48691e-10, 
    7.496293e-10, 7.477022e-10, 7.401967e-10, 7.424025e-10, 7.358236e-10, 
    7.31868e-10, 7.292403e-10, 7.273758e-10, 7.276394e-10, 7.281419e-10, 
    7.307241e-10, 7.331519e-10, 7.35002e-10, 7.362396e-10, 7.37459e-10, 
    7.411504e-10, 7.431039e-10, 7.474782e-10, 7.466887e-10, 7.480261e-10, 
    7.493037e-10, 7.514488e-10, 7.510957e-10, 7.520408e-10, 7.479908e-10, 
    7.506825e-10, 7.462391e-10, 7.474544e-10, 7.377909e-10, 7.341089e-10, 
    7.325442e-10, 7.311745e-10, 7.278421e-10, 7.301433e-10, 7.292362e-10, 
    7.313943e-10, 7.327657e-10, 7.320874e-10, 7.362735e-10, 7.346461e-10, 
    7.432197e-10, 7.395268e-10, 7.491547e-10, 7.468507e-10, 7.497069e-10, 
    7.482495e-10, 7.507467e-10, 7.484992e-10, 7.523925e-10, 7.532402e-10, 
    7.526609e-10, 7.548863e-10, 7.483746e-10, 7.508754e-10, 7.320685e-10, 
    7.321791e-10, 7.326944e-10, 7.304291e-10, 7.302905e-10, 7.282145e-10, 
    7.300617e-10, 7.308484e-10, 7.328452e-10, 7.340263e-10, 7.351492e-10, 
    7.376179e-10, 7.40375e-10, 7.442304e-10, 7.470001e-10, 7.488568e-10, 
    7.477183e-10, 7.487234e-10, 7.475998e-10, 7.470731e-10, 7.529226e-10, 
    7.496381e-10, 7.545662e-10, 7.542935e-10, 7.520632e-10, 7.543242e-10, 
    7.322568e-10, 7.316202e-10, 7.294101e-10, 7.311396e-10, 7.279884e-10, 
    7.297524e-10, 7.307667e-10, 7.346802e-10, 7.355399e-10, 7.363372e-10, 
    7.379118e-10, 7.399327e-10, 7.434778e-10, 7.465623e-10, 7.49378e-10, 
    7.491717e-10, 7.492443e-10, 7.498734e-10, 7.483152e-10, 7.501292e-10, 
    7.504337e-10, 7.496376e-10, 7.54257e-10, 7.529373e-10, 7.542877e-10, 
    7.534284e-10, 7.318271e-10, 7.328982e-10, 7.323194e-10, 7.334078e-10, 
    7.326411e-10, 7.360506e-10, 7.370728e-10, 7.418561e-10, 7.39893e-10, 
    7.430172e-10, 7.402103e-10, 7.407077e-10, 7.431193e-10, 7.40362e-10, 
    7.463923e-10, 7.423041e-10, 7.498979e-10, 7.458154e-10, 7.501537e-10, 
    7.493658e-10, 7.506702e-10, 7.518385e-10, 7.533081e-10, 7.5602e-10, 
    7.55392e-10, 7.576599e-10, 7.34495e-10, 7.358844e-10, 7.35762e-10, 
    7.372158e-10, 7.382912e-10, 7.406216e-10, 7.443595e-10, 7.429539e-10, 
    7.455343e-10, 7.460523e-10, 7.42132e-10, 7.445391e-10, 7.368141e-10, 
    7.380623e-10, 7.373191e-10, 7.346047e-10, 7.432778e-10, 7.388268e-10, 
    7.470459e-10, 7.446346e-10, 7.516719e-10, 7.481722e-10, 7.550464e-10, 
    7.579852e-10, 7.607508e-10, 7.639832e-10, 7.366425e-10, 7.356985e-10, 
    7.373888e-10, 7.397274e-10, 7.418971e-10, 7.447817e-10, 7.450768e-10, 
    7.456172e-10, 7.47017e-10, 7.48194e-10, 7.457882e-10, 7.48489e-10, 
    7.383519e-10, 7.436642e-10, 7.353417e-10, 7.378478e-10, 7.395895e-10, 
    7.388254e-10, 7.427932e-10, 7.437284e-10, 7.475286e-10, 7.455641e-10, 
    7.572599e-10, 7.520853e-10, 7.664441e-10, 7.624315e-10, 7.353687e-10, 
    7.366392e-10, 7.410613e-10, 7.389573e-10, 7.449742e-10, 7.464553e-10, 
    7.476593e-10, 7.491984e-10, 7.493646e-10, 7.502765e-10, 7.487821e-10, 
    7.502174e-10, 7.447878e-10, 7.472142e-10, 7.405558e-10, 7.421764e-10, 
    7.414309e-10, 7.406131e-10, 7.43137e-10, 7.458261e-10, 7.458834e-10, 
    7.467457e-10, 7.491757e-10, 7.449986e-10, 7.57928e-10, 7.499433e-10, 
    7.380247e-10, 7.404721e-10, 7.408216e-10, 7.398736e-10, 7.463068e-10, 
    7.439759e-10, 7.502542e-10, 7.485574e-10, 7.513377e-10, 7.499561e-10, 
    7.497529e-10, 7.479784e-10, 7.468737e-10, 7.440827e-10, 7.418118e-10, 
    7.400111e-10, 7.404298e-10, 7.424079e-10, 7.459905e-10, 7.493797e-10, 
    7.486373e-10, 7.511264e-10, 7.44538e-10, 7.473007e-10, 7.462329e-10, 
    7.49017e-10, 7.429165e-10, 7.481117e-10, 7.415886e-10, 7.421606e-10, 
    7.439296e-10, 7.474881e-10, 7.482752e-10, 7.491159e-10, 7.485971e-10, 
    7.460815e-10, 7.456693e-10, 7.438866e-10, 7.433944e-10, 7.42036e-10, 
    7.409114e-10, 7.41939e-10, 7.43018e-10, 7.460825e-10, 7.488442e-10, 
    7.518551e-10, 7.525919e-10, 7.561102e-10, 7.532463e-10, 7.579725e-10, 
    7.539546e-10, 7.609097e-10, 7.484126e-10, 7.538362e-10, 7.440101e-10, 
    7.450686e-10, 7.469834e-10, 7.513748e-10, 7.490039e-10, 7.517766e-10, 
    7.456532e-10, 7.424762e-10, 7.416541e-10, 7.401205e-10, 7.416892e-10, 
    7.415616e-10, 7.430627e-10, 7.425803e-10, 7.461842e-10, 7.442483e-10, 
    7.497478e-10, 7.517547e-10, 7.574222e-10, 7.608967e-10, 7.644334e-10, 
    7.659948e-10, 7.664701e-10, 7.666687e-10 ;

 SOIL2C =
  5.784044, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784102, 5.784096, 5.784097, 5.784091, 5.784057, 5.784063, 
    5.784057, 5.784057, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.78407, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784084, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784057, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784088, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784052, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784051, 5.78406, 5.784057, 5.784073, 
    5.784066, 5.784085, 5.784081, 5.784086, 5.784083, 5.784089, 5.784084, 
    5.784091, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784051, 
    5.784052, 5.784053, 5.784048, 5.784048, 5.784044, 5.784048, 5.784049, 
    5.784053, 5.784055, 5.784058, 5.784062, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784084, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784095, 5.784091, 5.784095, 5.784052, 5.78405, 5.784046, 
    5.78405, 5.784043, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.78408, 5.784086, 5.784085, 5.784085, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784095, 5.784093, 
    5.784095, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784087, 
    5.784086, 5.784088, 5.784091, 5.784093, 5.784099, 5.784098, 5.784102, 
    5.784056, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.784079, 5.784071, 5.784076, 5.784061, 5.784063, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784076, 5.78409, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784114, 5.78406, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784077, 5.784078, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784074, 5.784058, 5.784063, 
    5.784066, 5.784065, 5.784073, 5.784075, 5.784082, 5.784078, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.78406, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784085, 5.784086, 5.784088, 5.784085, 
    5.784087, 5.784077, 5.784081, 5.784068, 5.784071, 5.78407, 5.784069, 
    5.784073, 5.784079, 5.784079, 5.784081, 5.784085, 5.784077, 5.784102, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784067, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.784089, 5.784076, 5.784081, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784083, 5.784085, 
    5.784084, 5.784079, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.784079, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784094, 5.784075, 
    5.784077, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.78407, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784087, 5.784091, 5.784101, 5.784109, 5.784115, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086051e-09, 1.090831e-09, 1.089902e-09, 1.093757e-09, 1.091618e-09, 
    1.094143e-09, 1.08702e-09, 1.091021e-09, 1.088467e-09, 1.086482e-09, 
    1.101238e-09, 1.093929e-09, 1.10883e-09, 1.104169e-09, 1.115879e-09, 
    1.108105e-09, 1.117446e-09, 1.115654e-09, 1.121047e-09, 1.119502e-09, 
    1.1264e-09, 1.12176e-09, 1.129975e-09, 1.125292e-09, 1.126024e-09, 
    1.121607e-09, 1.0954e-09, 1.100328e-09, 1.095108e-09, 1.095811e-09, 
    1.095495e-09, 1.091663e-09, 1.089731e-09, 1.085686e-09, 1.08642e-09, 
    1.089391e-09, 1.096127e-09, 1.09384e-09, 1.099602e-09, 1.099472e-09, 
    1.105887e-09, 1.102994e-09, 1.113776e-09, 1.110712e-09, 1.119566e-09, 
    1.11734e-09, 1.119462e-09, 1.118818e-09, 1.11947e-09, 1.116204e-09, 
    1.117604e-09, 1.11473e-09, 1.103536e-09, 1.106826e-09, 1.097014e-09, 
    1.091115e-09, 1.087196e-09, 1.084415e-09, 1.084808e-09, 1.085558e-09, 
    1.089409e-09, 1.09303e-09, 1.095789e-09, 1.097635e-09, 1.099453e-09, 
    1.104958e-09, 1.107872e-09, 1.114396e-09, 1.113218e-09, 1.115213e-09, 
    1.117118e-09, 1.120317e-09, 1.11979e-09, 1.1212e-09, 1.11516e-09, 
    1.119174e-09, 1.112548e-09, 1.11436e-09, 1.099948e-09, 1.094457e-09, 
    1.092123e-09, 1.09008e-09, 1.085111e-09, 1.088543e-09, 1.08719e-09, 
    1.090408e-09, 1.092454e-09, 1.091442e-09, 1.097685e-09, 1.095258e-09, 
    1.108045e-09, 1.102537e-09, 1.116896e-09, 1.11346e-09, 1.117719e-09, 
    1.115546e-09, 1.11927e-09, 1.115918e-09, 1.121724e-09, 1.122989e-09, 
    1.122125e-09, 1.125443e-09, 1.115732e-09, 1.119462e-09, 1.091414e-09, 
    1.091579e-09, 1.092347e-09, 1.088969e-09, 1.088762e-09, 1.085666e-09, 
    1.088421e-09, 1.089594e-09, 1.092572e-09, 1.094334e-09, 1.096008e-09, 
    1.09969e-09, 1.103802e-09, 1.109552e-09, 1.113683e-09, 1.116451e-09, 
    1.114754e-09, 1.116253e-09, 1.114577e-09, 1.113792e-09, 1.122515e-09, 
    1.117617e-09, 1.124966e-09, 1.124559e-09, 1.121233e-09, 1.124605e-09, 
    1.091695e-09, 1.090745e-09, 1.087449e-09, 1.090029e-09, 1.085329e-09, 
    1.08796e-09, 1.089472e-09, 1.095309e-09, 1.096591e-09, 1.09778e-09, 
    1.100129e-09, 1.103143e-09, 1.10843e-09, 1.11303e-09, 1.117229e-09, 
    1.116921e-09, 1.117029e-09, 1.117968e-09, 1.115644e-09, 1.118349e-09, 
    1.118803e-09, 1.117616e-09, 1.124505e-09, 1.122537e-09, 1.124551e-09, 
    1.123269e-09, 1.091054e-09, 1.092651e-09, 1.091788e-09, 1.093411e-09, 
    1.092268e-09, 1.097353e-09, 1.098877e-09, 1.106011e-09, 1.103083e-09, 
    1.107743e-09, 1.103556e-09, 1.104298e-09, 1.107895e-09, 1.103783e-09, 
    1.112776e-09, 1.106679e-09, 1.118004e-09, 1.111916e-09, 1.118386e-09, 
    1.117211e-09, 1.119156e-09, 1.120898e-09, 1.12309e-09, 1.127134e-09, 
    1.126198e-09, 1.12958e-09, 1.095033e-09, 1.097105e-09, 1.096922e-09, 
    1.099091e-09, 1.100694e-09, 1.10417e-09, 1.109744e-09, 1.107648e-09, 
    1.111496e-09, 1.112269e-09, 1.106422e-09, 1.110012e-09, 1.098492e-09, 
    1.100353e-09, 1.099245e-09, 1.095196e-09, 1.108131e-09, 1.101493e-09, 
    1.113751e-09, 1.110155e-09, 1.12065e-09, 1.115431e-09, 1.125682e-09, 
    1.130065e-09, 1.134189e-09, 1.13901e-09, 1.098236e-09, 1.096828e-09, 
    1.099349e-09, 1.102836e-09, 1.106072e-09, 1.110374e-09, 1.110814e-09, 
    1.11162e-09, 1.113708e-09, 1.115463e-09, 1.111875e-09, 1.115903e-09, 
    1.100785e-09, 1.108707e-09, 1.096295e-09, 1.100033e-09, 1.102631e-09, 
    1.101491e-09, 1.107408e-09, 1.108803e-09, 1.114471e-09, 1.111541e-09, 
    1.128983e-09, 1.121266e-09, 1.14268e-09, 1.136696e-09, 1.096336e-09, 
    1.098231e-09, 1.104826e-09, 1.101688e-09, 1.110661e-09, 1.11287e-09, 
    1.114666e-09, 1.116961e-09, 1.117209e-09, 1.118569e-09, 1.11634e-09, 
    1.118481e-09, 1.110383e-09, 1.114002e-09, 1.104072e-09, 1.106489e-09, 
    1.105377e-09, 1.104157e-09, 1.107921e-09, 1.111932e-09, 1.112017e-09, 
    1.113303e-09, 1.116927e-09, 1.110698e-09, 1.12998e-09, 1.118072e-09, 
    1.100297e-09, 1.103947e-09, 1.104468e-09, 1.103054e-09, 1.112649e-09, 
    1.109172e-09, 1.118536e-09, 1.116005e-09, 1.120151e-09, 1.118091e-09, 
    1.117788e-09, 1.115142e-09, 1.113494e-09, 1.109332e-09, 1.105945e-09, 
    1.103259e-09, 1.103884e-09, 1.106834e-09, 1.112177e-09, 1.117231e-09, 
    1.116124e-09, 1.119836e-09, 1.110011e-09, 1.114131e-09, 1.112538e-09, 
    1.11669e-09, 1.107592e-09, 1.11534e-09, 1.105612e-09, 1.106465e-09, 
    1.109103e-09, 1.11441e-09, 1.115584e-09, 1.116838e-09, 1.116064e-09, 
    1.112313e-09, 1.111698e-09, 1.109039e-09, 1.108305e-09, 1.106279e-09, 
    1.104602e-09, 1.106135e-09, 1.107744e-09, 1.112314e-09, 1.116433e-09, 
    1.120923e-09, 1.122022e-09, 1.127269e-09, 1.122998e-09, 1.130046e-09, 
    1.124054e-09, 1.134426e-09, 1.115789e-09, 1.123877e-09, 1.109223e-09, 
    1.110802e-09, 1.113657e-09, 1.120207e-09, 1.116671e-09, 1.120806e-09, 
    1.111674e-09, 1.106936e-09, 1.10571e-09, 1.103423e-09, 1.105762e-09, 
    1.105572e-09, 1.10781e-09, 1.107091e-09, 1.112466e-09, 1.109579e-09, 
    1.11778e-09, 1.120773e-09, 1.129225e-09, 1.134407e-09, 1.139681e-09, 
    1.142009e-09, 1.142718e-09, 1.143014e-09 ;

 SOIL2C_TO_SOIL3C =
  7.757511e-11, 7.79165e-11, 7.785013e-11, 7.812549e-11, 7.797274e-11, 
    7.815305e-11, 7.764431e-11, 7.793006e-11, 7.774764e-11, 7.760583e-11, 
    7.865988e-11, 7.813777e-11, 7.920217e-11, 7.88692e-11, 7.970562e-11, 
    7.915036e-11, 7.981758e-11, 7.968959e-11, 8.007477e-11, 7.996442e-11, 
    8.045712e-11, 8.01257e-11, 8.071251e-11, 8.037797e-11, 8.04303e-11, 
    8.011477e-11, 7.824284e-11, 7.859489e-11, 7.822198e-11, 7.827219e-11, 
    7.824966e-11, 7.79759e-11, 7.783795e-11, 7.7549e-11, 7.760146e-11, 
    7.781368e-11, 7.829476e-11, 7.813145e-11, 7.854301e-11, 7.853371e-11, 
    7.899191e-11, 7.878532e-11, 7.955542e-11, 7.933654e-11, 7.996903e-11, 
    7.980997e-11, 7.996156e-11, 7.991559e-11, 7.996216e-11, 7.972888e-11, 
    7.982882e-11, 7.962355e-11, 7.882401e-11, 7.9059e-11, 7.835817e-11, 
    7.793677e-11, 7.765685e-11, 7.745822e-11, 7.74863e-11, 7.753984e-11, 
    7.781492e-11, 7.807355e-11, 7.827064e-11, 7.840248e-11, 7.853238e-11, 
    7.892561e-11, 7.913371e-11, 7.959969e-11, 7.951558e-11, 7.965805e-11, 
    7.979414e-11, 8.002264e-11, 7.998503e-11, 8.00857e-11, 7.965428e-11, 
    7.994101e-11, 7.946768e-11, 7.959714e-11, 7.856773e-11, 7.81755e-11, 
    7.800881e-11, 7.786289e-11, 7.75079e-11, 7.775305e-11, 7.765641e-11, 
    7.788632e-11, 7.803241e-11, 7.796015e-11, 7.840608e-11, 7.823272e-11, 
    7.914604e-11, 7.875265e-11, 7.977827e-11, 7.953285e-11, 7.98371e-11, 
    7.968184e-11, 7.994786e-11, 7.970845e-11, 8.012317e-11, 8.021347e-11, 
    8.015177e-11, 8.038881e-11, 7.969517e-11, 7.996157e-11, 7.795813e-11, 
    7.796992e-11, 7.802482e-11, 7.778349e-11, 7.776873e-11, 7.754757e-11, 
    7.774435e-11, 7.782815e-11, 7.804087e-11, 7.81667e-11, 7.828631e-11, 
    7.85493e-11, 7.884302e-11, 7.925371e-11, 7.954876e-11, 7.974653e-11, 
    7.962525e-11, 7.973232e-11, 7.961264e-11, 7.955653e-11, 8.017964e-11, 
    7.982976e-11, 8.035472e-11, 8.032567e-11, 8.00881e-11, 8.032894e-11, 
    7.797819e-11, 7.791037e-11, 7.767494e-11, 7.785918e-11, 7.752348e-11, 
    7.77114e-11, 7.781945e-11, 7.823635e-11, 7.832793e-11, 7.841287e-11, 
    7.858061e-11, 7.879589e-11, 7.917354e-11, 7.950211e-11, 7.980206e-11, 
    7.978009e-11, 7.978782e-11, 7.985483e-11, 7.968885e-11, 7.988208e-11, 
    7.991451e-11, 7.982971e-11, 8.032178e-11, 8.01812e-11, 8.032505e-11, 
    8.023352e-11, 7.793242e-11, 7.804652e-11, 7.798486e-11, 7.810081e-11, 
    7.801913e-11, 7.838234e-11, 7.849124e-11, 7.900079e-11, 7.879166e-11, 
    7.912448e-11, 7.882547e-11, 7.887845e-11, 7.913534e-11, 7.884162e-11, 
    7.948401e-11, 7.90485e-11, 7.985743e-11, 7.942255e-11, 7.988469e-11, 
    7.980076e-11, 7.993971e-11, 8.006416e-11, 8.022071e-11, 8.050959e-11, 
    8.044269e-11, 8.068426e-11, 7.821663e-11, 7.836463e-11, 7.83516e-11, 
    7.850647e-11, 7.862102e-11, 7.886928e-11, 7.926746e-11, 7.911773e-11, 
    7.93926e-11, 7.944779e-11, 7.903018e-11, 7.928659e-11, 7.846368e-11, 
    7.859664e-11, 7.851747e-11, 7.822831e-11, 7.915224e-11, 7.867808e-11, 
    7.955363e-11, 7.929677e-11, 8.004641e-11, 7.967361e-11, 8.040587e-11, 
    8.071892e-11, 8.101352e-11, 8.135782e-11, 7.84454e-11, 7.834483e-11, 
    7.852489e-11, 7.877402e-11, 7.900515e-11, 7.931244e-11, 7.934387e-11, 
    7.940144e-11, 7.955055e-11, 7.967593e-11, 7.941965e-11, 7.970735e-11, 
    7.862749e-11, 7.919339e-11, 7.830682e-11, 7.85738e-11, 7.875933e-11, 
    7.867794e-11, 7.910061e-11, 7.920023e-11, 7.960505e-11, 7.939578e-11, 
    8.064166e-11, 8.009045e-11, 8.161997e-11, 8.119254e-11, 7.83097e-11, 
    7.844505e-11, 7.891612e-11, 7.869198e-11, 7.933295e-11, 7.949073e-11, 
    7.961897e-11, 7.978293e-11, 7.980062e-11, 7.989777e-11, 7.973858e-11, 
    7.989148e-11, 7.931309e-11, 7.957156e-11, 7.886226e-11, 7.903491e-11, 
    7.895548e-11, 7.886837e-11, 7.913723e-11, 7.942369e-11, 7.94298e-11, 
    7.952165e-11, 7.97805e-11, 7.933555e-11, 8.071283e-11, 7.986227e-11, 
    7.859264e-11, 7.885335e-11, 7.889058e-11, 7.878959e-11, 7.947491e-11, 
    7.922659e-11, 7.98954e-11, 7.971464e-11, 8.00108e-11, 7.986364e-11, 
    7.984199e-11, 7.965296e-11, 7.953529e-11, 7.923798e-11, 7.899607e-11, 
    7.880424e-11, 7.884884e-11, 7.905957e-11, 7.944121e-11, 7.980223e-11, 
    7.972315e-11, 7.99883e-11, 7.928647e-11, 7.958077e-11, 7.946703e-11, 
    7.97636e-11, 7.911375e-11, 7.966717e-11, 7.897229e-11, 7.903322e-11, 
    7.922166e-11, 7.960074e-11, 7.968459e-11, 7.977413e-11, 7.971888e-11, 
    7.94509e-11, 7.940699e-11, 7.921708e-11, 7.916465e-11, 7.901995e-11, 
    7.890015e-11, 7.900961e-11, 7.912456e-11, 7.9451e-11, 7.974519e-11, 
    8.006593e-11, 8.014442e-11, 8.05192e-11, 8.021412e-11, 8.071756e-11, 
    8.028957e-11, 8.103044e-11, 7.969922e-11, 8.027696e-11, 7.923023e-11, 
    7.9343e-11, 7.954697e-11, 8.001477e-11, 7.97622e-11, 8.005756e-11, 
    7.940527e-11, 7.906684e-11, 7.897927e-11, 7.881591e-11, 7.898301e-11, 
    7.896941e-11, 7.912931e-11, 7.907793e-11, 7.946184e-11, 7.925562e-11, 
    7.984145e-11, 8.005523e-11, 8.065895e-11, 8.102906e-11, 8.140578e-11, 
    8.15721e-11, 8.162273e-11, 8.164389e-11 ;

 SOIL2C_vr =
  20.00646, 20.00647, 20.00647, 20.00648, 20.00648, 20.00648, 20.00646, 
    20.00647, 20.00647, 20.00646, 20.00651, 20.00648, 20.00654, 20.00652, 
    20.00656, 20.00653, 20.00657, 20.00656, 20.00658, 20.00657, 20.0066, 
    20.00658, 20.00661, 20.00659, 20.0066, 20.00658, 20.00649, 20.00651, 
    20.00649, 20.00649, 20.00649, 20.00648, 20.00647, 20.00645, 20.00646, 
    20.00647, 20.00649, 20.00648, 20.0065, 20.0065, 20.00653, 20.00652, 
    20.00655, 20.00654, 20.00657, 20.00657, 20.00657, 20.00657, 20.00657, 
    20.00656, 20.00657, 20.00656, 20.00652, 20.00653, 20.00649, 20.00647, 
    20.00646, 20.00645, 20.00645, 20.00645, 20.00647, 20.00648, 20.00649, 
    20.0065, 20.0065, 20.00652, 20.00653, 20.00656, 20.00655, 20.00656, 
    20.00657, 20.00658, 20.00657, 20.00658, 20.00656, 20.00657, 20.00655, 
    20.00656, 20.00651, 20.00649, 20.00648, 20.00647, 20.00645, 20.00647, 
    20.00646, 20.00647, 20.00648, 20.00648, 20.0065, 20.00649, 20.00653, 
    20.00652, 20.00657, 20.00655, 20.00657, 20.00656, 20.00657, 20.00656, 
    20.00658, 20.00659, 20.00658, 20.0066, 20.00656, 20.00657, 20.00648, 
    20.00648, 20.00648, 20.00647, 20.00647, 20.00645, 20.00646, 20.00647, 
    20.00648, 20.00648, 20.00649, 20.0065, 20.00652, 20.00654, 20.00655, 
    20.00656, 20.00656, 20.00656, 20.00656, 20.00655, 20.00658, 20.00657, 
    20.00659, 20.00659, 20.00658, 20.00659, 20.00648, 20.00647, 20.00646, 
    20.00647, 20.00645, 20.00646, 20.00647, 20.00649, 20.00649, 20.0065, 
    20.00651, 20.00652, 20.00653, 20.00655, 20.00657, 20.00657, 20.00657, 
    20.00657, 20.00656, 20.00657, 20.00657, 20.00657, 20.00659, 20.00658, 
    20.00659, 20.00659, 20.00647, 20.00648, 20.00648, 20.00648, 20.00648, 
    20.0065, 20.0065, 20.00653, 20.00652, 20.00653, 20.00652, 20.00652, 
    20.00653, 20.00652, 20.00655, 20.00653, 20.00657, 20.00655, 20.00657, 
    20.00657, 20.00657, 20.00658, 20.00659, 20.0066, 20.0066, 20.00661, 
    20.00649, 20.0065, 20.00649, 20.0065, 20.00651, 20.00652, 20.00654, 
    20.00653, 20.00655, 20.00655, 20.00653, 20.00654, 20.0065, 20.00651, 
    20.0065, 20.00649, 20.00653, 20.00651, 20.00655, 20.00654, 20.00658, 
    20.00656, 20.0066, 20.00661, 20.00663, 20.00664, 20.0065, 20.00649, 
    20.0065, 20.00652, 20.00653, 20.00654, 20.00654, 20.00655, 20.00655, 
    20.00656, 20.00655, 20.00656, 20.00651, 20.00654, 20.00649, 20.00651, 
    20.00652, 20.00651, 20.00653, 20.00654, 20.00656, 20.00655, 20.00661, 
    20.00658, 20.00665, 20.00663, 20.00649, 20.0065, 20.00652, 20.00651, 
    20.00654, 20.00655, 20.00656, 20.00657, 20.00657, 20.00657, 20.00656, 
    20.00657, 20.00654, 20.00656, 20.00652, 20.00653, 20.00653, 20.00652, 
    20.00653, 20.00655, 20.00655, 20.00655, 20.00657, 20.00654, 20.00661, 
    20.00657, 20.00651, 20.00652, 20.00652, 20.00652, 20.00655, 20.00654, 
    20.00657, 20.00656, 20.00658, 20.00657, 20.00657, 20.00656, 20.00655, 
    20.00654, 20.00653, 20.00652, 20.00652, 20.00653, 20.00655, 20.00657, 
    20.00656, 20.00657, 20.00654, 20.00656, 20.00655, 20.00657, 20.00653, 
    20.00656, 20.00653, 20.00653, 20.00654, 20.00656, 20.00656, 20.00657, 
    20.00656, 20.00655, 20.00655, 20.00654, 20.00653, 20.00653, 20.00652, 
    20.00653, 20.00653, 20.00655, 20.00656, 20.00658, 20.00658, 20.0066, 
    20.00659, 20.00661, 20.00659, 20.00663, 20.00656, 20.00659, 20.00654, 
    20.00654, 20.00655, 20.00658, 20.00657, 20.00658, 20.00655, 20.00653, 
    20.00653, 20.00652, 20.00653, 20.00653, 20.00653, 20.00653, 20.00655, 
    20.00654, 20.00657, 20.00658, 20.00661, 20.00663, 20.00665, 20.00665, 
    20.00665, 20.00666,
  20.00607, 20.00609, 20.00609, 20.00611, 20.0061, 20.00611, 20.00607, 
    20.00609, 20.00608, 20.00607, 20.00614, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00617, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00625, 20.00626, 20.00624, 20.00611, 20.00614, 
    20.00611, 20.00611, 20.00611, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00608, 20.00612, 20.00611, 20.00613, 20.00613, 20.00616, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00622, 20.00623, 
    20.00621, 20.00622, 20.0062, 20.00615, 20.00617, 20.00612, 20.00609, 
    20.00607, 20.00606, 20.00606, 20.00607, 20.00608, 20.0061, 20.00611, 
    20.00612, 20.00613, 20.00616, 20.00617, 20.0062, 20.0062, 20.00621, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.0062, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00607, 20.00609, 20.0061, 20.00609, 20.00612, 20.00611, 20.00617, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00624, 20.00624, 20.00626, 20.00621, 20.00623, 20.00609, 
    20.0061, 20.0061, 20.00608, 20.00608, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00613, 20.00615, 20.00618, 20.0062, 
    20.00621, 20.0062, 20.00621, 20.0062, 20.0062, 20.00624, 20.00622, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00607, 
    20.00609, 20.00607, 20.00608, 20.00608, 20.00611, 20.00612, 20.00612, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00622, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00624, 20.00609, 20.0061, 20.0061, 20.0061, 20.0061, 
    20.00612, 20.00613, 20.00616, 20.00615, 20.00617, 20.00615, 20.00616, 
    20.00617, 20.00615, 20.0062, 20.00617, 20.00622, 20.00619, 20.00622, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00626, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00618, 
    20.00617, 20.00619, 20.00619, 20.00617, 20.00618, 20.00613, 20.00614, 
    20.00613, 20.00611, 20.00617, 20.00614, 20.0062, 20.00618, 20.00623, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00613, 20.00615, 20.00616, 20.00618, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.00619, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00614, 20.00617, 20.00618, 20.0062, 20.00619, 20.00627, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00614, 
    20.00619, 20.0062, 20.0062, 20.00622, 20.00622, 20.00622, 20.00621, 
    20.00622, 20.00618, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00617, 20.00619, 20.00619, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00615, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00622, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00616, 20.00615, 20.00615, 20.00617, 20.00619, 20.00622, 
    20.00621, 20.00623, 20.00618, 20.0062, 20.0062, 20.00621, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.0062, 20.00621, 20.00621, 
    20.00621, 20.00619, 20.00619, 20.00618, 20.00617, 20.00616, 20.00616, 
    20.00616, 20.00617, 20.00619, 20.00621, 20.00624, 20.00624, 20.00626, 
    20.00624, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00623, 20.00621, 20.00623, 20.00619, 20.00617, 
    20.00616, 20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00623, 20.00627, 20.0063, 20.00632, 20.00633, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00552, 
    20.00554, 20.00553, 20.00552, 20.0056, 20.00556, 20.00563, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00572, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00564, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00566, 20.00561, 20.00562, 20.00558, 20.00554, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00555, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.00569, 20.00569, 20.0057, 20.00567, 20.00569, 20.00565, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00551, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00567, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00553, 20.00553, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00566, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00571, 20.0057, 20.00571, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00557, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00571, 20.0057, 
    20.00571, 20.00571, 20.00554, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00558, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00558, 20.00559, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.00569, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00557, 
    20.00559, 20.0056, 20.00562, 20.00564, 20.00564, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.00559, 20.00563, 20.00557, 20.00559, 
    20.0056, 20.0056, 20.00563, 20.00563, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.0058, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00564, 20.00566, 20.00566, 20.00568, 20.00568, 20.00568, 20.00567, 
    20.00568, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00564, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00561, 20.00561, 20.00565, 20.00564, 
    20.00568, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00562, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00565, 20.00567, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00567, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00561, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00576, 20.00567, 20.00571, 20.00564, 
    20.00564, 20.00566, 20.00569, 20.00567, 20.0057, 20.00565, 20.00562, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00565, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00576, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.0051, 20.0051, 20.00512, 20.00511, 20.00512, 20.00508, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.00519, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00525, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.0052, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00518, 20.00513, 20.00511, 
    20.00508, 20.00507, 20.00507, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00517, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00508, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.00509, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00521, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00514, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00525, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00513, 20.00515, 20.00515, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00515, 20.00519, 20.00513, 20.00515, 
    20.00516, 20.00516, 20.00519, 20.00519, 20.00522, 20.00521, 20.00529, 
    20.00526, 20.00536, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.0052, 20.00521, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.0052, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00518, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00523, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00523, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00525, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00523, 20.00525, 20.00521, 20.00518, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00536, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00446, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00438, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.00439, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00445, 20.00448, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00442, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00445, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00444, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258258, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.5258269, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258233, 0.5258234, 
    0.5258234, 0.5258229, 0.5258226, 0.5258222, 0.5258223, 0.5258226, 
    0.5258234, 0.5258232, 0.5258238, 0.5258238, 0.5258246, 0.5258242, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258262, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258243, 0.5258247, 
    0.5258235, 0.5258228, 0.5258223, 0.525822, 0.525822, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258236, 0.5258238, 0.5258245, 
    0.5258248, 0.5258256, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.5258229, 0.5258227, 0.5258221, 0.5258225, 
    0.5258223, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258248, 0.5258242, 0.5258259, 0.5258255, 0.525826, 0.5258258, 
    0.5258262, 0.5258258, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258262, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258225, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.525825, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.5258239, 0.5258243, 0.5258249, 0.5258255, 
    0.525826, 0.5258259, 0.525826, 0.525826, 0.5258258, 0.5258261, 0.5258262, 
    0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 0.5258228, 
    0.525823, 0.5258229, 0.5258231, 0.525823, 0.5258236, 0.5258238, 
    0.5258246, 0.5258242, 0.5258248, 0.5258243, 0.5258244, 0.5258248, 
    0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258253, 0.5258261, 
    0.525826, 0.5258262, 0.5258264, 0.5258267, 0.5258272, 0.5258271, 
    0.5258275, 0.5258233, 0.5258235, 0.5258235, 0.5258238, 0.525824, 
    0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 0.5258247, 
    0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258233, 0.5258249, 
    0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258257, 0.525827, 
    0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 0.5258238, 
    0.5258242, 0.5258246, 0.5258251, 0.5258252, 0.5258253, 0.5258256, 
    0.5258257, 0.5258253, 0.5258258, 0.525824, 0.525825, 0.5258235, 
    0.5258239, 0.5258242, 0.5258241, 0.5258248, 0.525825, 0.5258256, 
    0.5258253, 0.5258274, 0.5258265, 0.525829, 0.5258283, 0.5258235, 
    0.5258237, 0.5258245, 0.5258241, 0.5258252, 0.5258254, 0.5258257, 
    0.5258259, 0.525826, 0.5258262, 0.5258259, 0.5258262, 0.5258251, 
    0.5258256, 0.5258244, 0.5258247, 0.5258245, 0.5258244, 0.5258248, 
    0.5258253, 0.5258253, 0.5258255, 0.5258259, 0.5258252, 0.5258275, 
    0.5258261, 0.525824, 0.5258244, 0.5258244, 0.5258242, 0.5258254, 
    0.525825, 0.5258262, 0.5258259, 0.5258263, 0.5258261, 0.525826, 
    0.5258257, 0.5258255, 0.525825, 0.5258246, 0.5258243, 0.5258244, 
    0.5258247, 0.5258254, 0.525826, 0.5258259, 0.5258263, 0.5258251, 
    0.5258256, 0.5258254, 0.5258259, 0.5258248, 0.5258257, 0.5258246, 
    0.5258247, 0.525825, 0.5258256, 0.5258258, 0.5258259, 0.5258259, 
    0.5258254, 0.5258253, 0.525825, 0.5258249, 0.5258247, 0.5258244, 
    0.5258247, 0.5258248, 0.5258254, 0.5258259, 0.5258264, 0.5258266, 
    0.5258272, 0.5258267, 0.5258275, 0.5258268, 0.5258281, 0.5258258, 
    0.5258268, 0.525825, 0.5258252, 0.5258256, 0.5258263, 0.5258259, 
    0.5258264, 0.5258253, 0.5258247, 0.5258246, 0.5258243, 0.5258246, 
    0.5258245, 0.5258248, 0.5258248, 0.5258254, 0.5258251, 0.525826, 
    0.5258264, 0.5258274, 0.5258281, 0.5258287, 0.525829, 0.525829, 0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  2.569961e-21, 1.798972e-20, 2.569961e-21, 1.541976e-20, 5.139921e-21, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, 1.027984e-20, -1.28498e-20, 
    5.139921e-21, 1.28498e-20, 1.28498e-20, -7.709882e-21, 1.027984e-20, 
    -1.027984e-20, -1.798972e-20, -5.139921e-21, 1.003089e-36, 2.569961e-21, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, 5.139921e-21, -1.28498e-20, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    -1.28498e-20, 7.709882e-21, 2.312965e-20, 2.569961e-21, -1.027984e-20, 
    7.709882e-21, 2.055969e-20, 2.055969e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-21, -1.28498e-20, 5.015443e-37, -1.798972e-20, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, 1.798972e-20, -2.312965e-20, -1.027984e-20, 
    2.826957e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    1.798972e-20, 1.28498e-20, -1.541976e-20, -1.003089e-36, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -2.055969e-20, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, 2.569961e-21, -1.003089e-36, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -1.541976e-20, -2.055969e-20, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -2.312965e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, 1.541976e-20, -1.798972e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 7.709882e-21, 0, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 1.027984e-20, -1.003089e-36, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 1.28498e-20, 5.139921e-21, -1.003089e-36, 
    -1.798972e-20, -1.541976e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -2.055969e-20, -1.28498e-20, 7.709882e-21, 1.28498e-20, 
    2.055969e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, 1.541976e-20, -1.28498e-20, 
    1.027984e-20, -1.28498e-20, -1.541976e-20, 2.569961e-21, -7.709882e-21, 
    -1.027984e-20, -5.139921e-21, -2.055969e-20, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, 1.003089e-36, 
    2.569961e-21, 7.709882e-21, 2.055969e-20, 2.569961e-21, -7.709882e-21, 
    1.003089e-36, -2.569961e-21, -1.798972e-20, 1.027984e-20, -7.709882e-21, 
    5.139921e-21, -1.003089e-36, 2.569961e-21, 1.003089e-36, -1.003089e-36, 
    -5.139921e-21, -1.541976e-20, -2.569961e-21, -1.28498e-20, 1.541976e-20, 
    -1.027984e-20, 5.139921e-21, 1.28498e-20, -1.28498e-20, -5.139921e-21, 
    1.003089e-36, 1.027984e-20, -1.003089e-36, -1.541976e-20, -1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, 2.569961e-21, -2.569961e-21, 
    1.541976e-20, 5.139921e-21, 7.709882e-21, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 1.003089e-36, 
    1.798972e-20, -5.139921e-21, -7.709882e-21, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, 1.027984e-20, 5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -7.709882e-21, -1.027984e-20, -1.541976e-20, 
    2.312965e-20, 5.139921e-21, 1.027984e-20, 0, -1.28498e-20, -5.139921e-21, 
    -1.798972e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 1.541976e-20, 2.569961e-21, 
    1.003089e-36, -1.027984e-20, 5.139921e-21, 2.569961e-21, 2.312965e-20, 
    5.139921e-21, 7.709882e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.28498e-20, -7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, 0, 5.139921e-21, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.003089e-36, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    -1.798972e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 1.003089e-36, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 2.055969e-20, 0, 5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -1.027984e-20, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, 1.28498e-20, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -7.709882e-21, 1.28498e-20, 1.027984e-20, 
    5.139921e-21, -2.055969e-20, -5.139921e-21, 0, -2.569961e-21, 
    -1.027984e-20, -2.055969e-20, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, 7.709882e-21, 1.003089e-36, -7.709882e-21, -1.541976e-20, 
    -1.28498e-20, -2.569961e-20, -7.709882e-21, 7.709882e-21, 0, 2.826957e-20,
  -2.569961e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, -1.027984e-20, 
    5.139921e-21, -1.28498e-20, 1.003089e-36, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -7.709882e-21, -1.28498e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, -7.709882e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, 0, 7.709882e-21, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -1.28498e-20, -1.027984e-20, 0, 7.709882e-21, 1.28498e-20, -1.798972e-20, 
    5.139921e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, -1.28498e-20, -1.027984e-20, 1.541976e-20, 2.569961e-21, 
    1.28498e-20, 1.003089e-36, -1.027984e-20, 7.709882e-21, -1.027984e-20, 0, 
    -5.139921e-21, -5.139921e-21, -1.28498e-20, -1.027984e-20, -1.003089e-36, 
    0, -1.28498e-20, 7.709882e-21, 0, 0, -5.139921e-21, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    0, 1.28498e-20, -2.569961e-21, -1.027984e-20, 0, -5.139921e-21, 
    -1.003089e-36, -5.139921e-21, 0, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 1.541976e-20, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.312965e-20, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -7.709882e-21, 0, 0, -2.569961e-21, 
    1.003089e-36, -1.027984e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 0, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, -7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 1.003089e-36, -1.28498e-20, 0, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 1.027984e-20, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, 0, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 0, 1.027984e-20, -2.569961e-21, 2.569961e-21, -1.28498e-20, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, 5.139921e-21, 0, -7.709882e-21, -2.569961e-21, -5.139921e-21, 0, 
    5.139921e-21, -2.569961e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 0, 
    7.709882e-21, 5.139921e-21, -2.569961e-21, -1.003089e-36, -5.139921e-21, 
    1.541976e-20, -1.027984e-20, 7.709882e-21, 1.541976e-20, 0, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 0, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 0, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 1.541976e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    1.003089e-36, -2.569961e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -7.709882e-21, 1.541976e-20, 1.003089e-36, -1.027984e-20, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 
    0, -1.28498e-20, 1.28498e-20, 1.003089e-36, 0, -1.003089e-36, 
    -1.798972e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 1.003089e-36, 
    -2.569961e-21, -1.28498e-20, 5.139921e-21, -1.027984e-20, -7.709882e-21, 
    0, 1.541976e-20, 2.569961e-21, -1.28498e-20, 0, -7.709882e-21, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 0, -5.139921e-21, 
    7.709882e-21, 5.139921e-21, 0, 0, 1.28498e-20, -5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 1.541976e-20, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, -1.28498e-20, -5.139921e-21, -2.055969e-20, -1.798972e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 0, 1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.312965e-20, 
    -2.569961e-21, -7.709882e-21, 1.28498e-20, 5.139921e-21, -1.027984e-20, 
    7.709882e-21, 1.003089e-36, 1.027984e-20, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 1.541976e-20, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21,
  7.709882e-21, 2.569961e-21, 2.569961e-21, 1.541976e-20, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, 7.709882e-21, 1.003089e-36, 1.027984e-20, 
    -5.139921e-21, 7.709882e-21, -1.541976e-20, 2.569961e-21, -1.28498e-20, 
    -1.027984e-20, -1.28498e-20, 7.709882e-21, 7.709882e-21, 1.798972e-20, 
    2.569961e-21, 0, 7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, 1.027984e-20, 1.798972e-20, 
    -7.709882e-21, 1.027984e-20, 0, 2.569961e-21, 5.139921e-21, 1.003089e-36, 
    5.139921e-21, -2.569961e-21, 2.312965e-20, -1.027984e-20, 1.541976e-20, 
    -1.798972e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    2.312965e-20, 7.709882e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, -1.28498e-20, 0, 
    7.709882e-21, 0, -5.139921e-21, -1.027984e-20, 1.28498e-20, 
    -1.003089e-36, 1.027984e-20, -5.139921e-21, -1.28498e-20, -7.709882e-21, 
    1.003089e-36, -1.027984e-20, 1.798972e-20, -1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, -1.28498e-20, 
    1.003089e-36, 0, 2.569961e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    0, 2.569961e-21, 1.798972e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, 2.312965e-20, 
    -7.709882e-21, 1.541976e-20, -1.541976e-20, -1.28498e-20, 1.798972e-20, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    1.28498e-20, -1.541976e-20, 5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 2.055969e-20, -2.055969e-20, 
    7.709882e-21, 2.569961e-21, 5.139921e-21, -1.003089e-36, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 0, 
    7.709882e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    1.027984e-20, -1.003089e-36, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, 0, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, -2.569961e-21, 1.28498e-20, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 0, -2.569961e-21, 0, -5.139921e-21, 
    -1.28498e-20, 1.027984e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, 0, 7.709882e-21, -1.027984e-20, 0, 
    -1.541976e-20, -7.709882e-21, -1.003089e-36, -5.139921e-21, -1.28498e-20, 
    1.541976e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    0, 5.139921e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -1.28498e-20, 1.28498e-20, -2.569961e-21, 0, 1.027984e-20, 7.709882e-21, 
    1.28498e-20, 1.027984e-20, -7.709882e-21, 0, 2.569961e-21, 1.003089e-36, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -1.28498e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, -7.709882e-21, 0, 5.139921e-21, 
    -1.541976e-20, 2.569961e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, 
    -7.709882e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -1.027984e-20, 1.541976e-20, -1.027984e-20, -2.569961e-21, 
    0, -5.139921e-21, -7.709882e-21, 0, -1.28498e-20, -1.541976e-20, 0, 
    -1.28498e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -5.139921e-21, 1.28498e-20, -1.28498e-20, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 0, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 1.798972e-20, -1.28498e-20, 
    -2.055969e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, 7.709882e-21, 1.541976e-20, -1.027984e-20, -7.709882e-21, 
    -1.28498e-20, 5.139921e-21, -1.003089e-36, 5.139921e-21, -1.798972e-20, 
    5.139921e-21, 5.139921e-21, -1.28498e-20, 5.139921e-21, -2.569961e-21, 
    7.709882e-21, -1.541976e-20, 7.709882e-21, 1.28498e-20, -1.28498e-20, 
    -7.709882e-21, -7.709882e-21, 1.027984e-20,
  1.541976e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 1.003089e-36, 1.28498e-20, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, 1.28498e-20, -1.798972e-20, 
    -5.139921e-21, -1.798972e-20, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, 1.28498e-20, 5.139921e-21, 1.28498e-20, -1.28498e-20, 
    7.709882e-21, 5.139921e-21, 0, -2.569961e-21, -1.027984e-20, 
    -1.003089e-36, 1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    0, -7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 7.709882e-21, 2.055969e-20, 1.541976e-20, 0, 5.139921e-21, 
    -1.003089e-36, 7.709882e-21, 2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -2.569961e-21, 1.798972e-20, -5.139921e-21, 7.709882e-21, -1.28498e-20, 
    2.569961e-21, 5.139921e-21, -1.541976e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, 0, 
    1.027984e-20, 0, -1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -2.055969e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, 7.709882e-21, -1.28498e-20, -1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.798972e-20, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, 0, -5.139921e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 7.709882e-21, 
    1.28498e-20, -7.709882e-21, -1.28498e-20, 2.569961e-21, 5.139921e-21, 
    -2.569961e-20, -5.139921e-21, -7.709882e-21, 1.027984e-20, 1.027984e-20, 
    1.003089e-36, 1.28498e-20, -2.569961e-21, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 7.709882e-21, 1.541976e-20, -7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 1.28498e-20, 1.027984e-20, 1.027984e-20, 
    -1.798972e-20, -1.003089e-36, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 7.709882e-21, 0, 
    5.139921e-21, 7.709882e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, 7.709882e-21, 1.798972e-20, 
    -1.28498e-20, 7.709882e-21, 2.569961e-21, -1.027984e-20, -1.541976e-20, 
    0, 1.027984e-20, 1.027984e-20, -7.709882e-21, 1.541976e-20, 2.569961e-21, 
    7.709882e-21, -1.541976e-20, -7.709882e-21, 0, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, 1.027984e-20, -2.569961e-21, 
    2.569961e-21, -1.28498e-20, 7.709882e-21, -1.003089e-36, 7.709882e-21, 
    2.055969e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 
    1.541976e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, -1.798972e-20, 
    1.003089e-36, 0, -7.709882e-21, -1.003089e-36, 1.28498e-20, 2.569961e-20, 
    1.027984e-20, 1.28498e-20, -5.139921e-21, 1.003089e-36, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, -1.28498e-20, 1.541976e-20, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, -1.541976e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, 2.569961e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -2.055969e-20, -1.798972e-20, -1.027984e-20, 0, 
    2.569961e-21, -2.312965e-20, 1.798972e-20, 1.003089e-36, 0, 7.709882e-21, 
    1.027984e-20, 1.027984e-20, 2.312965e-20, 5.139921e-21, 0, -1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 1.28498e-20, 7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, -1.027984e-20, 1.798972e-20, 
    5.139921e-21, 0, -2.569961e-21, 2.569961e-21, -5.139921e-21, 1.28498e-20, 
    5.139921e-21, 1.28498e-20, 1.28498e-20, 2.569961e-21, -1.798972e-20, 
    7.709882e-21, -1.798972e-20, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    7.709882e-21, -1.003089e-36, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, 1.28498e-20, 5.139921e-21, 
    1.28498e-20, 2.569961e-21, 0, -2.569961e-21, -2.569961e-21, 0, 
    -5.139921e-21, -1.003089e-36, 1.28498e-20, 5.139921e-21, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-20, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, -1.003089e-36, -1.003089e-36, 
    -2.569961e-21, 1.28498e-20, -1.798972e-20, -2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 0, -1.28498e-20, -1.027984e-20, -2.569961e-21, 
    2.312965e-20, 1.28498e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 1.28498e-20, 0, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 0, 7.709882e-21, 1.28498e-20, -2.569961e-21,
  1.798972e-20, -2.569961e-21, -1.28498e-20, 2.569961e-21, -7.709882e-21, 
    3.083953e-20, 1.798972e-20, 1.003089e-36, 7.709882e-21, -1.28498e-20, 
    -1.027984e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    -1.003089e-36, 2.055969e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -1.28498e-20, -2.569961e-21, -2.569961e-21, 1.28498e-20, -2.055969e-20, 
    -2.569961e-21, -2.569961e-20, 1.027984e-20, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, -1.003089e-36, -1.027984e-20, 1.28498e-20, -1.28498e-20, 
    1.003089e-36, 1.798972e-20, 1.28498e-20, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 1.798972e-20, 2.055969e-20, 1.798972e-20, -2.569961e-21, 
    1.003089e-36, 1.28498e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 2.569961e-21, -1.798972e-20, 
    1.003089e-36, 7.709882e-21, -5.139921e-21, 2.055969e-20, 2.569961e-21, 
    1.541976e-20, 5.139921e-21, -1.798972e-20, 7.709882e-21, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, -5.139921e-21, 1.027984e-20, 1.28498e-20, 
    1.28498e-20, 7.709882e-21, -5.139921e-21, 1.541976e-20, -2.055969e-20, 
    -1.798972e-20, -7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -2.055969e-20, 2.569961e-21, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, 0, 1.541976e-20, 2.055969e-20, 
    -2.312965e-20, 1.003089e-36, 1.28498e-20, -1.28498e-20, 7.709882e-21, 
    2.312965e-20, -1.28498e-20, -5.139921e-21, 1.541976e-20, -1.28498e-20, 
    1.027984e-20, -1.28498e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    1.027984e-20, -1.003089e-36, 2.312965e-20, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, -2.569961e-21, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, 1.28498e-20, 2.569961e-21, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, 5.139921e-21, 1.28498e-20, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 1.28498e-20, 
    1.003089e-36, 1.003089e-36, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    7.709882e-21, -1.541976e-20, 2.055969e-20, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, 1.798972e-20, -1.003089e-36, 5.139921e-21, 1.541976e-20, 
    1.027984e-20, 7.709882e-21, 1.28498e-20, -7.709882e-21, -2.569961e-20, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, 1.28498e-20, -1.798972e-20, 2.569961e-20, 0, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, 2.569961e-21, 1.28498e-20, 
    1.28498e-20, -2.055969e-20, 5.139921e-21, -1.798972e-20, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.003089e-36, -1.541976e-20, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 1.28498e-20, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 1.541976e-20, 1.541976e-20, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 1.003089e-36, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 0, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -1.541976e-20, 2.055969e-20, -1.28498e-20, 
    1.28498e-20, -1.541976e-20, 2.569961e-20, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, 1.798972e-20, -2.569961e-21, 1.28498e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, 2.055969e-20, -1.28498e-20, -7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 1.28498e-20, -1.28498e-20, 
    -5.139921e-21, 1.28498e-20, 0, 7.709882e-21, -1.28498e-20, -1.027984e-20, 
    1.798972e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 5.139921e-21, 
    2.826957e-20, 5.139921e-21, 7.709882e-21, -1.798972e-20, -5.015443e-37, 
    -1.027984e-20, -7.709882e-21, 1.541976e-20, -1.027984e-20, 2.569961e-21, 
    1.027984e-20, -7.709882e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, -1.541976e-20, 5.139921e-21, -1.003089e-36, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -1.003089e-36, -1.541976e-20, 
    -5.139921e-21, 1.28498e-20, 7.709882e-21, -2.569961e-20, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 0, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, 2.569961e-21, -1.003089e-36, 2.569961e-21, 
    -5.139921e-21, -1.027984e-20, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -2.312965e-20, 1.027984e-20, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, -1.28498e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, -1.28498e-20, 2.055969e-20, 
    -1.003089e-36, 7.709882e-21, -2.569961e-21, 2.055969e-20, -7.709882e-21, 
    -5.139921e-21, 1.003089e-36, -1.798972e-20, -1.027984e-20, 2.312965e-20, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    2.569961e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 1.28498e-20, -1.28498e-20, -1.28498e-20, 2.569961e-20, 
    7.709882e-21,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259424e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.25942e-29, 6.259417e-29, 6.259414e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259453e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259466e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259426e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.25944e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259458e-29, 6.259458e-29, 6.259458e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259441e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259413e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.259459e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.259419e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259421e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259461e-29, 6.259463e-29, 
    6.259462e-29, 6.259467e-29, 6.259453e-29, 6.259458e-29, 6.259421e-29, 
    6.259422e-29, 6.259422e-29, 6.259418e-29, 6.259417e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259427e-29, 
    6.259432e-29, 6.259438e-29, 6.259445e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259454e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.259429e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259455e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259455e-29, 6.259458e-29, 6.259461e-29, 6.259463e-29, 6.259469e-29, 
    6.259467e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259428e-29, 
    6.259431e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259443e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.25943e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259432e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.25943e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259455e-29, 6.259457e-29, 6.259455e-29, 
    6.259457e-29, 6.259446e-29, 6.259451e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259456e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.259449e-29, 
    6.259445e-29, 6.259457e-29, 6.259454e-29, 6.259459e-29, 6.259456e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.25944e-29, 
    6.259437e-29, 6.259438e-29, 6.259441e-29, 6.259449e-29, 6.259455e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259444e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259444e-29, 6.259444e-29, 6.259441e-29, 
    6.259438e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259453e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.25946e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.25946e-29, 6.259472e-29, 6.259479e-29, 6.259485e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.194043e-10, 2.203699e-10, 2.201822e-10, 2.20961e-10, 2.20529e-10, 
    2.210389e-10, 2.196001e-10, 2.204082e-10, 2.198923e-10, 2.194912e-10, 
    2.224724e-10, 2.209957e-10, 2.240061e-10, 2.230644e-10, 2.2543e-10, 
    2.238596e-10, 2.257467e-10, 2.253847e-10, 2.264741e-10, 2.26162e-10, 
    2.275555e-10, 2.266182e-10, 2.282778e-10, 2.273316e-10, 2.274796e-10, 
    2.265872e-10, 2.212929e-10, 2.222886e-10, 2.212339e-10, 2.213759e-10, 
    2.213122e-10, 2.205379e-10, 2.201477e-10, 2.193305e-10, 2.194789e-10, 
    2.200791e-10, 2.214397e-10, 2.209778e-10, 2.221418e-10, 2.221156e-10, 
    2.234115e-10, 2.228272e-10, 2.250052e-10, 2.243862e-10, 2.26175e-10, 
    2.257252e-10, 2.261539e-10, 2.260239e-10, 2.261556e-10, 2.254958e-10, 
    2.257785e-10, 2.251979e-10, 2.229366e-10, 2.236012e-10, 2.216191e-10, 
    2.204272e-10, 2.196355e-10, 2.190738e-10, 2.191532e-10, 2.193046e-10, 
    2.200826e-10, 2.208141e-10, 2.213715e-10, 2.217444e-10, 2.221118e-10, 
    2.232239e-10, 2.238125e-10, 2.251304e-10, 2.248926e-10, 2.252955e-10, 
    2.256804e-10, 2.263267e-10, 2.262203e-10, 2.26505e-10, 2.252848e-10, 
    2.260958e-10, 2.247571e-10, 2.251232e-10, 2.222118e-10, 2.211024e-10, 
    2.20631e-10, 2.202183e-10, 2.192142e-10, 2.199076e-10, 2.196343e-10, 
    2.202845e-10, 2.206977e-10, 2.204934e-10, 2.217546e-10, 2.212643e-10, 
    2.238474e-10, 2.227348e-10, 2.256355e-10, 2.249414e-10, 2.258019e-10, 
    2.253628e-10, 2.261152e-10, 2.25438e-10, 2.26611e-10, 2.268664e-10, 
    2.266919e-10, 2.273623e-10, 2.254005e-10, 2.261539e-10, 2.204876e-10, 
    2.20521e-10, 2.206762e-10, 2.199937e-10, 2.19952e-10, 2.193265e-10, 
    2.19883e-10, 2.2012e-10, 2.207217e-10, 2.210775e-10, 2.214158e-10, 
    2.221596e-10, 2.229903e-10, 2.241519e-10, 2.249864e-10, 2.255457e-10, 
    2.252027e-10, 2.255056e-10, 2.25167e-10, 2.250084e-10, 2.267707e-10, 
    2.257811e-10, 2.272659e-10, 2.271837e-10, 2.265118e-10, 2.27193e-10, 
    2.205444e-10, 2.203526e-10, 2.196867e-10, 2.202078e-10, 2.192583e-10, 
    2.197898e-10, 2.200954e-10, 2.212745e-10, 2.215336e-10, 2.217738e-10, 
    2.222482e-10, 2.228571e-10, 2.239252e-10, 2.248545e-10, 2.257028e-10, 
    2.256406e-10, 2.256625e-10, 2.25852e-10, 2.253826e-10, 2.259291e-10, 
    2.260208e-10, 2.25781e-10, 2.271727e-10, 2.267751e-10, 2.27182e-10, 
    2.269231e-10, 2.204149e-10, 2.207376e-10, 2.205632e-10, 2.208912e-10, 
    2.206602e-10, 2.216874e-10, 2.219954e-10, 2.234366e-10, 2.228451e-10, 
    2.237864e-10, 2.229407e-10, 2.230906e-10, 2.238171e-10, 2.229864e-10, 
    2.248033e-10, 2.235715e-10, 2.258594e-10, 2.246295e-10, 2.259365e-10, 
    2.256991e-10, 2.260921e-10, 2.264441e-10, 2.268869e-10, 2.277039e-10, 
    2.275147e-10, 2.281979e-10, 2.212187e-10, 2.216373e-10, 2.216005e-10, 
    2.220385e-10, 2.223625e-10, 2.230646e-10, 2.241908e-10, 2.237673e-10, 
    2.245447e-10, 2.247008e-10, 2.235197e-10, 2.242449e-10, 2.219175e-10, 
    2.222935e-10, 2.220696e-10, 2.212518e-10, 2.238649e-10, 2.225239e-10, 
    2.250002e-10, 2.242737e-10, 2.263939e-10, 2.253395e-10, 2.274105e-10, 
    2.282959e-10, 2.291291e-10, 2.301029e-10, 2.218658e-10, 2.215814e-10, 
    2.220906e-10, 2.227952e-10, 2.234489e-10, 2.24318e-10, 2.244069e-10, 
    2.245697e-10, 2.249915e-10, 2.25346e-10, 2.246212e-10, 2.254349e-10, 
    2.223808e-10, 2.239813e-10, 2.214738e-10, 2.222289e-10, 2.227537e-10, 
    2.225235e-10, 2.237189e-10, 2.240007e-10, 2.251456e-10, 2.245537e-10, 
    2.280774e-10, 2.265184e-10, 2.308443e-10, 2.296355e-10, 2.21482e-10, 
    2.218648e-10, 2.231971e-10, 2.225632e-10, 2.24376e-10, 2.248222e-10, 
    2.25185e-10, 2.256487e-10, 2.256987e-10, 2.259735e-10, 2.255233e-10, 
    2.259557e-10, 2.243199e-10, 2.250509e-10, 2.230448e-10, 2.235331e-10, 
    2.233084e-10, 2.230621e-10, 2.238225e-10, 2.246327e-10, 2.246499e-10, 
    2.249097e-10, 2.256418e-10, 2.243834e-10, 2.282787e-10, 2.258731e-10, 
    2.222822e-10, 2.230196e-10, 2.231249e-10, 2.228392e-10, 2.247775e-10, 
    2.240752e-10, 2.259668e-10, 2.254556e-10, 2.262932e-10, 2.25877e-10, 
    2.258157e-10, 2.252811e-10, 2.249483e-10, 2.241074e-10, 2.234232e-10, 
    2.228807e-10, 2.230068e-10, 2.236028e-10, 2.246822e-10, 2.257033e-10, 
    2.254796e-10, 2.262295e-10, 2.242446e-10, 2.250769e-10, 2.247552e-10, 
    2.25594e-10, 2.237561e-10, 2.253213e-10, 2.23356e-10, 2.235283e-10, 
    2.240613e-10, 2.251334e-10, 2.253705e-10, 2.256238e-10, 2.254675e-10, 
    2.247096e-10, 2.245854e-10, 2.240483e-10, 2.239e-10, 2.234908e-10, 
    2.231519e-10, 2.234615e-10, 2.237866e-10, 2.247099e-10, 2.255419e-10, 
    2.264491e-10, 2.266711e-10, 2.277311e-10, 2.268682e-10, 2.282921e-10, 
    2.270816e-10, 2.29177e-10, 2.254119e-10, 2.27046e-10, 2.240855e-10, 
    2.244044e-10, 2.249813e-10, 2.263044e-10, 2.255901e-10, 2.264254e-10, 
    2.245805e-10, 2.236234e-10, 2.233757e-10, 2.229137e-10, 2.233863e-10, 
    2.233478e-10, 2.238001e-10, 2.236547e-10, 2.247406e-10, 2.241573e-10, 
    2.258142e-10, 2.264188e-10, 2.281263e-10, 2.291731e-10, 2.302386e-10, 
    2.30709e-10, 2.308522e-10, 2.30912e-10 ;

 SOIL2N_TO_SOIL3N =
  1.567174e-11, 1.574071e-11, 1.57273e-11, 1.578293e-11, 1.575207e-11, 
    1.57885e-11, 1.568572e-11, 1.574345e-11, 1.570659e-11, 1.567795e-11, 
    1.589089e-11, 1.578541e-11, 1.600044e-11, 1.593317e-11, 1.610214e-11, 
    1.598997e-11, 1.612476e-11, 1.609891e-11, 1.617672e-11, 1.615443e-11, 
    1.625396e-11, 1.618701e-11, 1.630556e-11, 1.623797e-11, 1.624855e-11, 
    1.61848e-11, 1.580663e-11, 1.587775e-11, 1.580242e-11, 1.581256e-11, 
    1.580801e-11, 1.575271e-11, 1.572484e-11, 1.566647e-11, 1.567706e-11, 
    1.571993e-11, 1.581712e-11, 1.578413e-11, 1.586727e-11, 1.58654e-11, 
    1.595796e-11, 1.591623e-11, 1.60718e-11, 1.602759e-11, 1.615536e-11, 
    1.612323e-11, 1.615385e-11, 1.614456e-11, 1.615397e-11, 1.610684e-11, 
    1.612704e-11, 1.608557e-11, 1.592404e-11, 1.597151e-11, 1.582993e-11, 
    1.57448e-11, 1.568825e-11, 1.564813e-11, 1.56538e-11, 1.566461e-11, 
    1.572019e-11, 1.577243e-11, 1.581225e-11, 1.583888e-11, 1.586513e-11, 
    1.594457e-11, 1.598661e-11, 1.608074e-11, 1.606375e-11, 1.609254e-11, 
    1.612003e-11, 1.616619e-11, 1.615859e-11, 1.617893e-11, 1.609178e-11, 
    1.61497e-11, 1.605408e-11, 1.608023e-11, 1.587227e-11, 1.579303e-11, 
    1.575936e-11, 1.572988e-11, 1.565816e-11, 1.570769e-11, 1.568816e-11, 
    1.573461e-11, 1.576412e-11, 1.574952e-11, 1.583961e-11, 1.580459e-11, 
    1.59891e-11, 1.590963e-11, 1.611682e-11, 1.606724e-11, 1.612871e-11, 
    1.609734e-11, 1.615108e-11, 1.610272e-11, 1.61865e-11, 1.620474e-11, 
    1.619227e-11, 1.624017e-11, 1.610003e-11, 1.615385e-11, 1.574912e-11, 
    1.57515e-11, 1.576259e-11, 1.571384e-11, 1.571085e-11, 1.566617e-11, 
    1.570593e-11, 1.572286e-11, 1.576583e-11, 1.579125e-11, 1.581542e-11, 
    1.586855e-11, 1.592788e-11, 1.601085e-11, 1.607046e-11, 1.611041e-11, 
    1.608591e-11, 1.610754e-11, 1.608336e-11, 1.607203e-11, 1.619791e-11, 
    1.612722e-11, 1.623328e-11, 1.622741e-11, 1.617941e-11, 1.622807e-11, 
    1.575317e-11, 1.573947e-11, 1.569191e-11, 1.572913e-11, 1.566131e-11, 
    1.569927e-11, 1.57211e-11, 1.580532e-11, 1.582382e-11, 1.584098e-11, 
    1.587487e-11, 1.591836e-11, 1.599466e-11, 1.606103e-11, 1.612163e-11, 
    1.611719e-11, 1.611875e-11, 1.613229e-11, 1.609876e-11, 1.613779e-11, 
    1.614435e-11, 1.612722e-11, 1.622662e-11, 1.619822e-11, 1.622728e-11, 
    1.620879e-11, 1.574392e-11, 1.576697e-11, 1.575452e-11, 1.577794e-11, 
    1.576144e-11, 1.583482e-11, 1.585682e-11, 1.595975e-11, 1.591751e-11, 
    1.598474e-11, 1.592434e-11, 1.593504e-11, 1.598694e-11, 1.59276e-11, 
    1.605738e-11, 1.596939e-11, 1.613282e-11, 1.604496e-11, 1.613832e-11, 
    1.612137e-11, 1.614944e-11, 1.617458e-11, 1.62062e-11, 1.626456e-11, 
    1.625105e-11, 1.629985e-11, 1.580134e-11, 1.583124e-11, 1.58286e-11, 
    1.585989e-11, 1.588303e-11, 1.593319e-11, 1.601363e-11, 1.598338e-11, 
    1.603891e-11, 1.605006e-11, 1.596569e-11, 1.601749e-11, 1.585125e-11, 
    1.587811e-11, 1.586212e-11, 1.58037e-11, 1.599035e-11, 1.589456e-11, 
    1.607144e-11, 1.601955e-11, 1.617099e-11, 1.609568e-11, 1.624361e-11, 
    1.630685e-11, 1.636637e-11, 1.643592e-11, 1.584756e-11, 1.582724e-11, 
    1.586361e-11, 1.591394e-11, 1.596064e-11, 1.602271e-11, 1.602907e-11, 
    1.60407e-11, 1.607082e-11, 1.609615e-11, 1.604437e-11, 1.61025e-11, 
    1.588434e-11, 1.599867e-11, 1.581956e-11, 1.58735e-11, 1.591098e-11, 
    1.589453e-11, 1.597992e-11, 1.600005e-11, 1.608183e-11, 1.603955e-11, 
    1.629124e-11, 1.617989e-11, 1.648888e-11, 1.640253e-11, 1.582014e-11, 
    1.584748e-11, 1.594265e-11, 1.589737e-11, 1.602686e-11, 1.605873e-11, 
    1.608464e-11, 1.611776e-11, 1.612134e-11, 1.614096e-11, 1.610881e-11, 
    1.613969e-11, 1.602285e-11, 1.607506e-11, 1.593177e-11, 1.596665e-11, 
    1.59506e-11, 1.5933e-11, 1.598732e-11, 1.604519e-11, 1.604642e-11, 
    1.606498e-11, 1.611727e-11, 1.602738e-11, 1.630562e-11, 1.613379e-11, 
    1.58773e-11, 1.592997e-11, 1.593749e-11, 1.591709e-11, 1.605554e-11, 
    1.600537e-11, 1.614048e-11, 1.610397e-11, 1.61638e-11, 1.613407e-11, 
    1.612969e-11, 1.609151e-11, 1.606774e-11, 1.600767e-11, 1.59588e-11, 
    1.592005e-11, 1.592906e-11, 1.597163e-11, 1.604873e-11, 1.612166e-11, 
    1.610569e-11, 1.615925e-11, 1.601747e-11, 1.607692e-11, 1.605394e-11, 
    1.611386e-11, 1.598257e-11, 1.609438e-11, 1.5954e-11, 1.596631e-11, 
    1.600438e-11, 1.608096e-11, 1.60979e-11, 1.611599e-11, 1.610482e-11, 
    1.605069e-11, 1.604182e-11, 1.600345e-11, 1.599286e-11, 1.596363e-11, 
    1.593943e-11, 1.596154e-11, 1.598476e-11, 1.605071e-11, 1.611014e-11, 
    1.617493e-11, 1.619079e-11, 1.62665e-11, 1.620487e-11, 1.630658e-11, 
    1.622011e-11, 1.636979e-11, 1.610085e-11, 1.621757e-11, 1.600611e-11, 
    1.602889e-11, 1.607009e-11, 1.61646e-11, 1.611358e-11, 1.617325e-11, 
    1.604147e-11, 1.59731e-11, 1.595541e-11, 1.59224e-11, 1.595616e-11, 
    1.595342e-11, 1.598572e-11, 1.597534e-11, 1.60529e-11, 1.601124e-11, 
    1.612959e-11, 1.617277e-11, 1.629474e-11, 1.636951e-11, 1.644561e-11, 
    1.647921e-11, 1.648944e-11, 1.649371e-11 ;

 SOIL2N_vr =
  1.818769, 1.81877, 1.81877, 1.818771, 1.818771, 1.818771, 1.818769, 
    1.81877, 1.81877, 1.818769, 1.818774, 1.818771, 1.818776, 1.818775, 
    1.818778, 1.818776, 1.818779, 1.818778, 1.81878, 1.818779, 1.818782, 
    1.81878, 1.818783, 1.818781, 1.818782, 1.81878, 1.818772, 1.818773, 
    1.818772, 1.818772, 1.818772, 1.818771, 1.81877, 1.818769, 1.818769, 
    1.81877, 1.818772, 1.818771, 1.818773, 1.818773, 1.818775, 1.818774, 
    1.818778, 1.818777, 1.818779, 1.818779, 1.818779, 1.818779, 1.818779, 
    1.818778, 1.818779, 1.818778, 1.818774, 1.818775, 1.818772, 1.81877, 
    1.818769, 1.818768, 1.818768, 1.818769, 1.81877, 1.818771, 1.818772, 
    1.818772, 1.818773, 1.818775, 1.818776, 1.818778, 1.818777, 1.818778, 
    1.818779, 1.81878, 1.81878, 1.81878, 1.818778, 1.818779, 1.818777, 
    1.818778, 1.818773, 1.818771, 1.818771, 1.81877, 1.818769, 1.81877, 
    1.818769, 1.81877, 1.818771, 1.818771, 1.818773, 1.818772, 1.818776, 
    1.818774, 1.818779, 1.818778, 1.818779, 1.818778, 1.818779, 1.818778, 
    1.81878, 1.818781, 1.81878, 1.818781, 1.818778, 1.818779, 1.818771, 
    1.818771, 1.818771, 1.81877, 1.81877, 1.818769, 1.81877, 1.81877, 
    1.818771, 1.818771, 1.818772, 1.818773, 1.818774, 1.818776, 1.818778, 
    1.818779, 1.818778, 1.818778, 1.818778, 1.818778, 1.81878, 1.818779, 
    1.818781, 1.818781, 1.81878, 1.818781, 1.818771, 1.81877, 1.818769, 
    1.81877, 1.818769, 1.818769, 1.81877, 1.818772, 1.818772, 1.818773, 
    1.818773, 1.818774, 1.818776, 1.818777, 1.818779, 1.818779, 1.818779, 
    1.818779, 1.818778, 1.818779, 1.818779, 1.818779, 1.818781, 1.81878, 
    1.818781, 1.818781, 1.81877, 1.818771, 1.818771, 1.818771, 1.818771, 
    1.818772, 1.818773, 1.818775, 1.818774, 1.818776, 1.818774, 1.818775, 
    1.818776, 1.818774, 1.818777, 1.818775, 1.818779, 1.818777, 1.818779, 
    1.818779, 1.818779, 1.81878, 1.818781, 1.818782, 1.818782, 1.818783, 
    1.818772, 1.818772, 1.818772, 1.818773, 1.818774, 1.818775, 1.818776, 
    1.818776, 1.818777, 1.818777, 1.818775, 1.818776, 1.818773, 1.818773, 
    1.818773, 1.818772, 1.818776, 1.818774, 1.818778, 1.818776, 1.81878, 
    1.818778, 1.818781, 1.818783, 1.818784, 1.818786, 1.818773, 1.818772, 
    1.818773, 1.818774, 1.818775, 1.818777, 1.818777, 1.818777, 1.818778, 
    1.818778, 1.818777, 1.818778, 1.818774, 1.818776, 1.818772, 1.818773, 
    1.818774, 1.818774, 1.818776, 1.818776, 1.818778, 1.818777, 1.818782, 
    1.81878, 1.818787, 1.818785, 1.818772, 1.818773, 1.818775, 1.818774, 
    1.818777, 1.818777, 1.818778, 1.818779, 1.818779, 1.818779, 1.818779, 
    1.818779, 1.818777, 1.818778, 1.818775, 1.818775, 1.818775, 1.818775, 
    1.818776, 1.818777, 1.818777, 1.818778, 1.818779, 1.818777, 1.818783, 
    1.818779, 1.818773, 1.818774, 1.818775, 1.818774, 1.818777, 1.818776, 
    1.818779, 1.818778, 1.81878, 1.818779, 1.818779, 1.818778, 1.818778, 
    1.818776, 1.818775, 1.818774, 1.818774, 1.818775, 1.818777, 1.818779, 
    1.818778, 1.81878, 1.818776, 1.818778, 1.818777, 1.818779, 1.818776, 
    1.818778, 1.818775, 1.818775, 1.818776, 1.818778, 1.818778, 1.818779, 
    1.818778, 1.818777, 1.818777, 1.818776, 1.818776, 1.818775, 1.818775, 
    1.818775, 1.818776, 1.818777, 1.818779, 1.81878, 1.81878, 1.818782, 
    1.818781, 1.818783, 1.818781, 1.818784, 1.818778, 1.818781, 1.818776, 
    1.818777, 1.818778, 1.81878, 1.818779, 1.81878, 1.818777, 1.818775, 
    1.818775, 1.818774, 1.818775, 1.818775, 1.818776, 1.818776, 1.818777, 
    1.818776, 1.818779, 1.81878, 1.818783, 1.818784, 1.818786, 1.818787, 
    1.818787, 1.818787,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818743, 1.818741, 
    1.818746, 1.818743, 1.818747, 1.818746, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818752, 1.81875, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818733, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.818739, 1.818739, 1.818742, 1.818741, 
    1.818745, 1.818744, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818738, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818733, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.818739, 1.818742, 1.818743, 1.818746, 1.818745, 1.818746, 
    1.818747, 1.818748, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818737, 1.818736, 1.818735, 1.818733, 1.818735, 
    1.818734, 1.818735, 1.818736, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 
    1.818749, 1.818749, 1.818749, 1.818751, 1.818746, 1.818748, 1.818736, 
    1.818736, 1.818736, 1.818735, 1.818735, 1.818733, 1.818735, 1.818735, 
    1.818736, 1.818737, 1.818738, 1.818739, 1.818741, 1.818744, 1.818745, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818745, 1.818749, 1.818747, 
    1.81875, 1.81875, 1.818749, 1.81875, 1.818736, 1.818736, 1.818734, 
    1.818735, 1.818733, 1.818734, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818747, 1.818746, 1.818747, 1.818748, 1.818747, 1.81875, 1.818749, 
    1.81875, 1.81875, 1.818736, 1.818736, 1.818736, 1.818737, 1.818736, 
    1.818738, 1.818739, 1.818742, 1.818741, 1.818743, 1.818741, 1.818741, 
    1.818743, 1.818741, 1.818745, 1.818742, 1.818747, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818751, 1.818751, 1.818752, 
    1.818737, 1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818742, 1.818744, 1.818739, 1.81874, 
    1.818739, 1.818738, 1.818743, 1.81874, 1.818745, 1.818744, 1.818748, 
    1.818746, 1.818751, 1.818753, 1.818754, 1.818756, 1.818739, 1.818738, 
    1.818739, 1.818741, 1.818742, 1.818744, 1.818744, 1.818745, 1.818745, 
    1.818746, 1.818745, 1.818746, 1.81874, 1.818743, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818743, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818755, 1.818738, 1.818739, 1.818742, 1.81874, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818741, 1.818742, 1.818742, 1.818741, 
    1.818743, 1.818745, 1.818745, 1.818745, 1.818747, 1.818744, 1.818752, 
    1.818747, 1.81874, 1.818741, 1.818741, 1.818741, 1.818745, 1.818743, 
    1.818748, 1.818746, 1.818748, 1.818747, 1.818747, 1.818746, 1.818745, 
    1.818744, 1.818742, 1.818741, 1.818741, 1.818743, 1.818745, 1.818747, 
    1.818746, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818742, 1.818743, 1.818746, 1.818746, 1.818747, 
    1.818746, 1.818745, 1.818745, 1.818743, 1.818743, 1.818742, 1.818742, 
    1.818742, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818751, 
    1.818749, 1.818752, 1.81875, 1.818754, 1.818746, 1.81875, 1.818744, 
    1.818744, 1.818745, 1.818748, 1.818747, 1.818748, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818747, 1.818748, 1.818752, 1.818754, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818685, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818683, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818697, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818683, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818687, 1.818686, 1.818685, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818686, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818686, 1.818685, 1.818685, 1.818683, 1.818685, 1.818685, 
    1.818687, 1.818687, 1.818688, 1.81869, 1.818692, 1.818694, 1.818696, 
    1.818698, 1.818697, 1.818697, 1.818697, 1.818696, 1.8187, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818701, 1.818686, 1.818686, 1.818684, 
    1.818685, 1.818683, 1.818684, 1.818685, 1.818688, 1.818688, 1.818689, 
    1.81869, 1.818691, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818698, 1.818699, 1.818698, 1.818701, 1.8187, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818686, 
    1.818689, 1.818689, 1.818693, 1.818691, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818695, 1.818698, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818702, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.81869, 1.818692, 1.818694, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.818699, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818695, 1.818696, 
    1.818697, 1.818695, 1.818697, 1.81869, 1.818694, 1.818688, 1.81869, 
    1.818691, 1.818691, 1.818693, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.818709, 1.818707, 1.818688, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818697, 
    1.818699, 1.818695, 1.818696, 1.818692, 1.818693, 1.818692, 1.818692, 
    1.818694, 1.818695, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818691, 1.818696, 1.818694, 
    1.818699, 1.818697, 1.818699, 1.818698, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818691, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818697, 1.818699, 1.818695, 1.818696, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818697, 1.818696, 1.818695, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818702, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818695, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818694, 1.818698, 1.818699, 1.818703, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818643, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818657, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818643, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818646, 1.818645, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.81866, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818643, 1.818645, 1.818645, 
    1.818647, 1.818647, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818657, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818645, 1.818643, 1.818645, 1.818645, 1.818648, 1.818648, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818646, 
    1.818649, 1.81865, 1.818653, 1.818651, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.81866, 1.818662, 1.818662, 1.818663, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818654, 
    1.818653, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.818659, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.818669, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818658, 1.818657, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818655, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818651, 1.818656, 1.818654, 
    1.818658, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818651, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818656, 1.818656, 1.818658, 1.818653, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818662, 
    1.81866, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818659, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818586, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.81859, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818587, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.818589, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.81859, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.327396e-09, 1.333238e-09, 1.332102e-09, 1.336814e-09, 1.3342e-09, 
    1.337286e-09, 1.32858e-09, 1.33347e-09, 1.330349e-09, 1.327922e-09, 
    1.345958e-09, 1.337024e-09, 1.355237e-09, 1.34954e-09, 1.363852e-09, 
    1.354351e-09, 1.365767e-09, 1.363577e-09, 1.370168e-09, 1.36828e-09, 
    1.376711e-09, 1.37104e-09, 1.381081e-09, 1.375356e-09, 1.376252e-09, 
    1.370853e-09, 1.338822e-09, 1.344846e-09, 1.338465e-09, 1.339324e-09, 
    1.338939e-09, 1.334254e-09, 1.331894e-09, 1.32695e-09, 1.327847e-09, 
    1.331478e-09, 1.33971e-09, 1.336916e-09, 1.343958e-09, 1.343799e-09, 
    1.351639e-09, 1.348104e-09, 1.361282e-09, 1.357536e-09, 1.368359e-09, 
    1.365637e-09, 1.368231e-09, 1.367445e-09, 1.368241e-09, 1.36425e-09, 
    1.36596e-09, 1.362447e-09, 1.348766e-09, 1.352787e-09, 1.340795e-09, 
    1.333585e-09, 1.328795e-09, 1.325396e-09, 1.325877e-09, 1.326793e-09, 
    1.3315e-09, 1.335925e-09, 1.339298e-09, 1.341554e-09, 1.343776e-09, 
    1.350505e-09, 1.354066e-09, 1.362039e-09, 1.3606e-09, 1.363038e-09, 
    1.365366e-09, 1.369276e-09, 1.368633e-09, 1.370355e-09, 1.362973e-09, 
    1.367879e-09, 1.35978e-09, 1.361996e-09, 1.344381e-09, 1.33767e-09, 
    1.334818e-09, 1.332321e-09, 1.326246e-09, 1.330441e-09, 1.328787e-09, 
    1.332721e-09, 1.335221e-09, 1.333985e-09, 1.341615e-09, 1.338649e-09, 
    1.354277e-09, 1.347545e-09, 1.365095e-09, 1.360895e-09, 1.366101e-09, 
    1.363445e-09, 1.367997e-09, 1.3639e-09, 1.370996e-09, 1.372542e-09, 
    1.371486e-09, 1.375542e-09, 1.363673e-09, 1.368231e-09, 1.33395e-09, 
    1.334152e-09, 1.335091e-09, 1.330962e-09, 1.330709e-09, 1.326925e-09, 
    1.330292e-09, 1.331726e-09, 1.335366e-09, 1.337519e-09, 1.339566e-09, 
    1.344066e-09, 1.349092e-09, 1.356119e-09, 1.361168e-09, 1.364552e-09, 
    1.362477e-09, 1.364309e-09, 1.362261e-09, 1.361301e-09, 1.371963e-09, 
    1.365976e-09, 1.374959e-09, 1.374461e-09, 1.370396e-09, 1.374517e-09, 
    1.334293e-09, 1.333133e-09, 1.329104e-09, 1.332257e-09, 1.326513e-09, 
    1.329728e-09, 1.331577e-09, 1.338711e-09, 1.340278e-09, 1.341731e-09, 
    1.344602e-09, 1.348285e-09, 1.354747e-09, 1.360369e-09, 1.365502e-09, 
    1.365126e-09, 1.365258e-09, 1.366405e-09, 1.363565e-09, 1.366871e-09, 
    1.367426e-09, 1.365975e-09, 1.374395e-09, 1.371989e-09, 1.374451e-09, 
    1.372885e-09, 1.33351e-09, 1.335463e-09, 1.334408e-09, 1.336392e-09, 
    1.334994e-09, 1.341209e-09, 1.343072e-09, 1.351791e-09, 1.348213e-09, 
    1.353908e-09, 1.348791e-09, 1.349698e-09, 1.354094e-09, 1.349068e-09, 
    1.36006e-09, 1.352608e-09, 1.366449e-09, 1.359008e-09, 1.366916e-09, 
    1.36548e-09, 1.367857e-09, 1.369987e-09, 1.372665e-09, 1.377608e-09, 
    1.376464e-09, 1.380597e-09, 1.338373e-09, 1.340906e-09, 1.340683e-09, 
    1.343333e-09, 1.345293e-09, 1.349541e-09, 1.356354e-09, 1.353792e-09, 
    1.358496e-09, 1.35944e-09, 1.352294e-09, 1.356682e-09, 1.342601e-09, 
    1.344876e-09, 1.343521e-09, 1.338573e-09, 1.354383e-09, 1.346269e-09, 
    1.361251e-09, 1.356856e-09, 1.369683e-09, 1.363304e-09, 1.375834e-09, 
    1.38119e-09, 1.386231e-09, 1.392123e-09, 1.342288e-09, 1.340567e-09, 
    1.343648e-09, 1.347911e-09, 1.351866e-09, 1.357124e-09, 1.357662e-09, 
    1.358647e-09, 1.361198e-09, 1.363344e-09, 1.358959e-09, 1.363881e-09, 
    1.345404e-09, 1.355087e-09, 1.339917e-09, 1.344485e-09, 1.34766e-09, 
    1.346267e-09, 1.353499e-09, 1.355204e-09, 1.362131e-09, 1.35855e-09, 
    1.379868e-09, 1.370437e-09, 1.396608e-09, 1.389295e-09, 1.339966e-09, 
    1.342282e-09, 1.350342e-09, 1.346507e-09, 1.357475e-09, 1.360175e-09, 
    1.362369e-09, 1.365175e-09, 1.365477e-09, 1.36714e-09, 1.364416e-09, 
    1.367032e-09, 1.357135e-09, 1.361558e-09, 1.349421e-09, 1.352375e-09, 
    1.351016e-09, 1.349525e-09, 1.354126e-09, 1.359028e-09, 1.359132e-09, 
    1.360704e-09, 1.365133e-09, 1.357519e-09, 1.381086e-09, 1.366532e-09, 
    1.344807e-09, 1.349269e-09, 1.349906e-09, 1.348177e-09, 1.359904e-09, 
    1.355655e-09, 1.367099e-09, 1.364006e-09, 1.369074e-09, 1.366556e-09, 
    1.366185e-09, 1.362951e-09, 1.360937e-09, 1.35585e-09, 1.351711e-09, 
    1.348428e-09, 1.349191e-09, 1.352797e-09, 1.359327e-09, 1.365505e-09, 
    1.364152e-09, 1.368689e-09, 1.35668e-09, 1.361715e-09, 1.359769e-09, 
    1.364844e-09, 1.353724e-09, 1.363194e-09, 1.351304e-09, 1.352346e-09, 
    1.355571e-09, 1.362057e-09, 1.363492e-09, 1.365024e-09, 1.364079e-09, 
    1.359493e-09, 1.358742e-09, 1.355492e-09, 1.354595e-09, 1.352119e-09, 
    1.350069e-09, 1.351942e-09, 1.353909e-09, 1.359495e-09, 1.364529e-09, 
    1.370017e-09, 1.37136e-09, 1.377773e-09, 1.372553e-09, 1.381167e-09, 
    1.373844e-09, 1.386521e-09, 1.363742e-09, 1.373628e-09, 1.355717e-09, 
    1.357647e-09, 1.361137e-09, 1.369141e-09, 1.36482e-09, 1.369874e-09, 
    1.358712e-09, 1.352922e-09, 1.351423e-09, 1.348628e-09, 1.351487e-09, 
    1.351254e-09, 1.35399e-09, 1.353111e-09, 1.35968e-09, 1.356152e-09, 
    1.366176e-09, 1.369834e-09, 1.380164e-09, 1.386497e-09, 1.392943e-09, 
    1.395789e-09, 1.396656e-09, 1.397018e-09 ;

 SOIL2_HR_S3 =
  9.481402e-11, 9.523128e-11, 9.515016e-11, 9.548672e-11, 9.530002e-11, 
    9.55204e-11, 9.489861e-11, 9.524785e-11, 9.50249e-11, 9.485157e-11, 
    9.613986e-11, 9.550172e-11, 9.680265e-11, 9.639569e-11, 9.741798e-11, 
    9.673932e-11, 9.755481e-11, 9.739839e-11, 9.786916e-11, 9.773429e-11, 
    9.833648e-11, 9.793141e-11, 9.864862e-11, 9.823974e-11, 9.830371e-11, 
    9.791806e-11, 9.563014e-11, 9.606042e-11, 9.560465e-11, 9.5666e-11, 
    9.563847e-11, 9.530388e-11, 9.513527e-11, 9.478212e-11, 9.484623e-11, 
    9.51056e-11, 9.569359e-11, 9.549399e-11, 9.599702e-11, 9.598566e-11, 
    9.654567e-11, 9.629317e-11, 9.72344e-11, 9.696689e-11, 9.773993e-11, 
    9.754551e-11, 9.77308e-11, 9.767461e-11, 9.773152e-11, 9.744641e-11, 
    9.756856e-11, 9.731767e-11, 9.634046e-11, 9.662766e-11, 9.577109e-11, 
    9.525605e-11, 9.491393e-11, 9.467116e-11, 9.470548e-11, 9.477091e-11, 
    9.510712e-11, 9.542322e-11, 9.566412e-11, 9.582525e-11, 9.598402e-11, 
    9.646463e-11, 9.671898e-11, 9.72885e-11, 9.718571e-11, 9.735984e-11, 
    9.752617e-11, 9.780545e-11, 9.775948e-11, 9.788253e-11, 9.735523e-11, 
    9.770568e-11, 9.712717e-11, 9.72854e-11, 9.602722e-11, 9.554784e-11, 
    9.534411e-11, 9.516576e-11, 9.473187e-11, 9.50315e-11, 9.491339e-11, 
    9.519439e-11, 9.537295e-11, 9.528463e-11, 9.582966e-11, 9.561777e-11, 
    9.673406e-11, 9.625323e-11, 9.750677e-11, 9.720681e-11, 9.757867e-11, 
    9.738892e-11, 9.771405e-11, 9.742143e-11, 9.792832e-11, 9.80387e-11, 
    9.796327e-11, 9.8253e-11, 9.740522e-11, 9.77308e-11, 9.528216e-11, 
    9.529656e-11, 9.536366e-11, 9.506871e-11, 9.505067e-11, 9.478036e-11, 
    9.502087e-11, 9.51233e-11, 9.538329e-11, 9.553708e-11, 9.568327e-11, 
    9.60047e-11, 9.636368e-11, 9.686564e-11, 9.722625e-11, 9.746799e-11, 
    9.731976e-11, 9.745062e-11, 9.730433e-11, 9.723576e-11, 9.799734e-11, 
    9.756971e-11, 9.821133e-11, 9.817582e-11, 9.788546e-11, 9.817982e-11, 
    9.530667e-11, 9.522379e-11, 9.493603e-11, 9.516123e-11, 9.475092e-11, 
    9.49806e-11, 9.511266e-11, 9.56222e-11, 9.573414e-11, 9.583796e-11, 
    9.604298e-11, 9.63061e-11, 9.676766e-11, 9.716925e-11, 9.753585e-11, 
    9.750899e-11, 9.751844e-11, 9.760034e-11, 9.739748e-11, 9.763365e-11, 
    9.767329e-11, 9.756965e-11, 9.817107e-11, 9.799925e-11, 9.817507e-11, 
    9.806319e-11, 9.525073e-11, 9.53902e-11, 9.531483e-11, 9.545655e-11, 
    9.535672e-11, 9.580064e-11, 9.593374e-11, 9.655651e-11, 9.630092e-11, 
    9.670769e-11, 9.634223e-11, 9.640699e-11, 9.672098e-11, 9.636198e-11, 
    9.714712e-11, 9.661483e-11, 9.760353e-11, 9.707201e-11, 9.763684e-11, 
    9.753427e-11, 9.770409e-11, 9.785619e-11, 9.804754e-11, 9.84006e-11, 
    9.831885e-11, 9.86141e-11, 9.55981e-11, 9.5779e-11, 9.576306e-11, 
    9.595236e-11, 9.609236e-11, 9.639579e-11, 9.688245e-11, 9.669944e-11, 
    9.703541e-11, 9.710285e-11, 9.659244e-11, 9.690584e-11, 9.590005e-11, 
    9.606256e-11, 9.59658e-11, 9.561237e-11, 9.674162e-11, 9.61621e-11, 
    9.723222e-11, 9.691827e-11, 9.78345e-11, 9.737885e-11, 9.827384e-11, 
    9.865646e-11, 9.901652e-11, 9.943734e-11, 9.587771e-11, 9.57548e-11, 
    9.597487e-11, 9.627936e-11, 9.656185e-11, 9.693742e-11, 9.697584e-11, 
    9.704621e-11, 9.722845e-11, 9.738169e-11, 9.706846e-11, 9.74201e-11, 
    9.610026e-11, 9.679192e-11, 9.570834e-11, 9.603464e-11, 9.626141e-11, 
    9.616193e-11, 9.667852e-11, 9.680028e-11, 9.729506e-11, 9.703929e-11, 
    9.856203e-11, 9.788833e-11, 9.975774e-11, 9.923532e-11, 9.571186e-11, 
    9.587728e-11, 9.645303e-11, 9.617909e-11, 9.696249e-11, 9.715533e-11, 
    9.731208e-11, 9.751247e-11, 9.75341e-11, 9.765283e-11, 9.745827e-11, 
    9.764514e-11, 9.693822e-11, 9.725413e-11, 9.638721e-11, 9.659822e-11, 
    9.650115e-11, 9.639467e-11, 9.672329e-11, 9.70734e-11, 9.708086e-11, 
    9.719313e-11, 9.750951e-11, 9.696566e-11, 9.864901e-11, 9.760944e-11, 
    9.605767e-11, 9.637632e-11, 9.642182e-11, 9.629839e-11, 9.713599e-11, 
    9.68325e-11, 9.764993e-11, 9.742901e-11, 9.779098e-11, 9.761111e-11, 
    9.758465e-11, 9.735363e-11, 9.72098e-11, 9.684642e-11, 9.655075e-11, 
    9.631629e-11, 9.637081e-11, 9.662836e-11, 9.709481e-11, 9.753606e-11, 
    9.74394e-11, 9.776348e-11, 9.690569e-11, 9.726538e-11, 9.712637e-11, 
    9.748884e-11, 9.669458e-11, 9.737098e-11, 9.652169e-11, 9.659615e-11, 
    9.682648e-11, 9.728979e-11, 9.739227e-11, 9.750172e-11, 9.743418e-11, 
    9.710665e-11, 9.705298e-11, 9.682088e-11, 9.67568e-11, 9.657994e-11, 
    9.643352e-11, 9.65673e-11, 9.670779e-11, 9.710678e-11, 9.746634e-11, 
    9.785836e-11, 9.795428e-11, 9.841235e-11, 9.803949e-11, 9.86548e-11, 
    9.813169e-11, 9.90372e-11, 9.741016e-11, 9.811629e-11, 9.683696e-11, 
    9.697478e-11, 9.722407e-11, 9.779582e-11, 9.748714e-11, 9.784814e-11, 
    9.705088e-11, 9.663725e-11, 9.653022e-11, 9.633055e-11, 9.653479e-11, 
    9.651818e-11, 9.671361e-11, 9.665081e-11, 9.712003e-11, 9.686798e-11, 
    9.758399e-11, 9.784528e-11, 9.858316e-11, 9.903552e-11, 9.949595e-11, 
    9.969923e-11, 9.976111e-11, 9.978698e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.617577e-11, 2.629094e-11, 2.626855e-11, 2.636144e-11, 2.630991e-11, 
    2.637074e-11, 2.619912e-11, 2.629551e-11, 2.623398e-11, 2.618613e-11, 
    2.654172e-11, 2.636559e-11, 2.672466e-11, 2.661233e-11, 2.68945e-11, 
    2.670718e-11, 2.693227e-11, 2.688909e-11, 2.701903e-11, 2.69818e-11, 
    2.714801e-11, 2.703621e-11, 2.723417e-11, 2.712131e-11, 2.713897e-11, 
    2.703252e-11, 2.640103e-11, 2.651979e-11, 2.639399e-11, 2.641093e-11, 
    2.640333e-11, 2.631098e-11, 2.626444e-11, 2.616696e-11, 2.618466e-11, 
    2.625625e-11, 2.641854e-11, 2.636345e-11, 2.650229e-11, 2.649916e-11, 
    2.665373e-11, 2.658404e-11, 2.684383e-11, 2.676999e-11, 2.698336e-11, 
    2.69297e-11, 2.698084e-11, 2.696533e-11, 2.698104e-11, 2.690234e-11, 
    2.693606e-11, 2.686681e-11, 2.659709e-11, 2.667636e-11, 2.643994e-11, 
    2.629778e-11, 2.620335e-11, 2.613634e-11, 2.614581e-11, 2.616387e-11, 
    2.625667e-11, 2.634392e-11, 2.641041e-11, 2.645488e-11, 2.649871e-11, 
    2.663136e-11, 2.670156e-11, 2.685876e-11, 2.683039e-11, 2.687845e-11, 
    2.692436e-11, 2.700144e-11, 2.698875e-11, 2.702272e-11, 2.687718e-11, 
    2.697391e-11, 2.681423e-11, 2.68579e-11, 2.651063e-11, 2.637831e-11, 
    2.632208e-11, 2.627285e-11, 2.61531e-11, 2.62358e-11, 2.62032e-11, 
    2.628076e-11, 2.633004e-11, 2.630567e-11, 2.64561e-11, 2.639761e-11, 
    2.670573e-11, 2.657301e-11, 2.691901e-11, 2.683621e-11, 2.693885e-11, 
    2.688648e-11, 2.697622e-11, 2.689545e-11, 2.703536e-11, 2.706582e-11, 
    2.7045e-11, 2.712497e-11, 2.689097e-11, 2.698084e-11, 2.630498e-11, 
    2.630896e-11, 2.632748e-11, 2.624607e-11, 2.624109e-11, 2.616648e-11, 
    2.623286e-11, 2.626114e-11, 2.63329e-11, 2.637534e-11, 2.64157e-11, 
    2.650441e-11, 2.66035e-11, 2.674205e-11, 2.684158e-11, 2.69083e-11, 
    2.686739e-11, 2.690351e-11, 2.686313e-11, 2.68442e-11, 2.705441e-11, 
    2.693638e-11, 2.711347e-11, 2.710367e-11, 2.702353e-11, 2.710477e-11, 
    2.631175e-11, 2.628887e-11, 2.620945e-11, 2.62716e-11, 2.615835e-11, 
    2.622175e-11, 2.62582e-11, 2.639884e-11, 2.642974e-11, 2.645839e-11, 
    2.651498e-11, 2.65876e-11, 2.6715e-11, 2.682585e-11, 2.692703e-11, 
    2.691962e-11, 2.692223e-11, 2.694483e-11, 2.688884e-11, 2.695402e-11, 
    2.696497e-11, 2.693636e-11, 2.710236e-11, 2.705493e-11, 2.710346e-11, 
    2.707258e-11, 2.629631e-11, 2.63348e-11, 2.6314e-11, 2.635312e-11, 
    2.632556e-11, 2.644809e-11, 2.648483e-11, 2.665672e-11, 2.658617e-11, 
    2.669845e-11, 2.659758e-11, 2.661545e-11, 2.670212e-11, 2.660303e-11, 
    2.681974e-11, 2.667282e-11, 2.694571e-11, 2.679901e-11, 2.695491e-11, 
    2.692659e-11, 2.697347e-11, 2.701545e-11, 2.706826e-11, 2.716571e-11, 
    2.714315e-11, 2.722464e-11, 2.639219e-11, 2.644212e-11, 2.643772e-11, 
    2.648997e-11, 2.652861e-11, 2.661236e-11, 2.674668e-11, 2.669617e-11, 
    2.67889e-11, 2.680752e-11, 2.666664e-11, 2.675314e-11, 2.647553e-11, 
    2.652038e-11, 2.649368e-11, 2.639613e-11, 2.670781e-11, 2.654786e-11, 
    2.684322e-11, 2.675657e-11, 2.700946e-11, 2.68837e-11, 2.713072e-11, 
    2.723633e-11, 2.733571e-11, 2.745186e-11, 2.646936e-11, 2.643544e-11, 
    2.649618e-11, 2.658022e-11, 2.665819e-11, 2.676186e-11, 2.677246e-11, 
    2.679188e-11, 2.684218e-11, 2.688448e-11, 2.679803e-11, 2.689508e-11, 
    2.653079e-11, 2.67217e-11, 2.642261e-11, 2.651268e-11, 2.657527e-11, 
    2.654781e-11, 2.66904e-11, 2.6724e-11, 2.686057e-11, 2.678997e-11, 
    2.721027e-11, 2.702432e-11, 2.754029e-11, 2.73961e-11, 2.642359e-11, 
    2.646925e-11, 2.662816e-11, 2.655255e-11, 2.676878e-11, 2.6822e-11, 
    2.686527e-11, 2.692058e-11, 2.692655e-11, 2.695932e-11, 2.690562e-11, 
    2.69572e-11, 2.676208e-11, 2.684927e-11, 2.660999e-11, 2.666823e-11, 
    2.664144e-11, 2.661205e-11, 2.670275e-11, 2.679939e-11, 2.680145e-11, 
    2.683244e-11, 2.691976e-11, 2.676965e-11, 2.723427e-11, 2.694734e-11, 
    2.651904e-11, 2.660699e-11, 2.661955e-11, 2.658548e-11, 2.681667e-11, 
    2.67329e-11, 2.695852e-11, 2.689754e-11, 2.699745e-11, 2.694781e-11, 
    2.69405e-11, 2.687674e-11, 2.683704e-11, 2.673674e-11, 2.665513e-11, 
    2.659042e-11, 2.660546e-11, 2.667655e-11, 2.68053e-11, 2.692709e-11, 
    2.690041e-11, 2.698986e-11, 2.67531e-11, 2.685238e-11, 2.681401e-11, 
    2.691406e-11, 2.669483e-11, 2.688152e-11, 2.664711e-11, 2.666766e-11, 
    2.673124e-11, 2.685911e-11, 2.68874e-11, 2.691761e-11, 2.689897e-11, 
    2.680857e-11, 2.679375e-11, 2.672969e-11, 2.6712e-11, 2.666319e-11, 
    2.662277e-11, 2.66597e-11, 2.669848e-11, 2.68086e-11, 2.690785e-11, 
    2.701605e-11, 2.704252e-11, 2.716895e-11, 2.706604e-11, 2.723587e-11, 
    2.709149e-11, 2.734142e-11, 2.689234e-11, 2.708724e-11, 2.673413e-11, 
    2.677217e-11, 2.684098e-11, 2.699879e-11, 2.691359e-11, 2.701322e-11, 
    2.679317e-11, 2.667901e-11, 2.664946e-11, 2.659435e-11, 2.665073e-11, 
    2.664614e-11, 2.670008e-11, 2.668275e-11, 2.681226e-11, 2.674269e-11, 
    2.694032e-11, 2.701244e-11, 2.72161e-11, 2.734095e-11, 2.746804e-11, 
    2.752415e-11, 2.754122e-11, 2.754836e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -1.003089e-36, 1.28498e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, 1.798972e-20, -5.139921e-21, 0, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -1.28498e-20, 7.709882e-21, 5.139921e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -1.28498e-20, 1.28498e-20, 
    2.312965e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-20, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -1.541976e-20, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 0, 7.709882e-21, -1.798972e-20, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -1.28498e-20, -1.027984e-20, 1.003089e-36, 2.569961e-21, 0, 1.541976e-20, 
    -1.027984e-20, 1.541976e-20, 1.28498e-20, -1.027984e-20, -2.055969e-20, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, 0, 1.28498e-20, -5.139921e-21, 1.798972e-20, 
    -1.027984e-20, 7.709882e-21, 7.709882e-21, -2.569961e-21, -1.003089e-36, 
    1.003089e-36, 5.139921e-21, 1.003089e-36, 1.28498e-20, -7.709882e-21, 
    -1.541976e-20, -7.709882e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, 1.541976e-20, 0, 0, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, 1.28498e-20, -1.28498e-20, 1.798972e-20, -2.569961e-21, 
    1.027984e-20, -1.027984e-20, -7.709882e-21, 2.312965e-20, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, -5.139921e-21, 
    1.28498e-20, -1.28498e-20, -1.541976e-20, -2.569961e-21, 1.027984e-20, 
    -1.28498e-20, 5.139921e-21, 1.003089e-36, 7.709882e-21, 0, -1.798972e-20, 
    1.28498e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, 1.003089e-36, 
    1.28498e-20, 2.569961e-21, 5.139921e-21, -1.28498e-20, 7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -7.709882e-21, 2.312965e-20, 2.055969e-20, 
    -1.003089e-36, 7.709882e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, 
    2.569961e-21, -2.055969e-20, -2.569961e-21, 1.28498e-20, -1.027984e-20, 
    -5.139921e-21, 0, -5.139921e-21, 1.027984e-20, -2.055969e-20, 
    7.709882e-21, -1.28498e-20, 1.28498e-20, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, 5.139921e-21, 7.709882e-21, 7.709882e-21, 0, 2.312965e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, 0, 7.709882e-21, 
    2.569961e-21, -1.003089e-36, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    1.798972e-20, 0, -1.027984e-20, 0, -1.003089e-36, 0, 2.569961e-21, 
    -2.312965e-20, 2.055969e-20, -1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -1.003089e-36, 0, -1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, -5.139921e-21, 2.055969e-20, 
    0, 7.709882e-21, -7.709882e-21, 1.541976e-20, 2.055969e-20, 7.709882e-21, 
    -7.709882e-21, 1.003089e-36, -1.003089e-36, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-20, -7.709882e-21, -2.569961e-21, 1.541976e-20, 
    -7.709882e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, -1.541976e-20, 1.003089e-36, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -1.027984e-20, 1.28498e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.312965e-20, 1.28498e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 1.541976e-20, 7.709882e-21, -1.28498e-20, 5.139921e-21, 
    -1.28498e-20, 7.709882e-21, 7.709882e-21, -1.003089e-36, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, -1.003089e-36, -7.709882e-21, -1.28498e-20, -2.569961e-21, 
    -1.003089e-36, -1.003089e-36, -1.003089e-36, 1.28498e-20, 2.569961e-21, 
    2.569961e-21, 1.003089e-36, -1.28498e-20, -5.139921e-21, -1.798972e-20, 
    1.003089e-36, 1.798972e-20, -1.541976e-20, 1.28498e-20, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -2.055969e-20, 
    1.027984e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -2.569961e-21, -7.709882e-21, 1.003089e-36, -7.709882e-21, 1.003089e-36, 
    5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    1.027984e-20, -5.139921e-21, -1.28498e-20, -1.541976e-20, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    0, 2.569961e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, 2.569961e-21, -1.28498e-20, 1.027984e-20, 
    -1.541976e-20, -1.027984e-20, -5.139921e-21, 1.28498e-20, -1.003089e-36,
  -2.569961e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    1.027984e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -1.541976e-20, 1.28498e-20, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 0, -2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, 1.003089e-36, 0, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, -1.541976e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.003089e-36, 7.709882e-21, -2.569961e-21, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, 0, -2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 2.569961e-21, 1.541976e-20, -1.541976e-20, 
    -2.569961e-21, 7.709882e-21, -1.027984e-20, -7.709882e-21, -5.139921e-21, 
    0, -2.569961e-21, -1.003089e-36, 7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, -2.055969e-20, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.003089e-36, -7.709882e-21, 0, 
    1.027984e-20, 1.027984e-20, 0, -1.027984e-20, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -1.027984e-20, 2.055969e-20, -7.709882e-21, 0, 1.798972e-20, 0, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 1.003089e-36, 
    1.28498e-20, 5.139921e-21, 1.541976e-20, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 0, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    2.569961e-21, 1.003089e-36, -2.569961e-21, 0, 5.139921e-21, 0, 
    -1.003089e-36, 0, 0, 2.569961e-21, -2.569961e-21, 0, 0, -7.709882e-21, 
    -5.139921e-21, -1.798972e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 1.027984e-20, 5.139921e-21, 0, -2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    0, 7.709882e-21, -1.027984e-20, 2.569961e-21, 0, 1.003089e-36, 
    1.027984e-20, 7.709882e-21, -1.003089e-36, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.541976e-20, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 0, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, 1.541976e-20, 7.709882e-21, 
    1.28498e-20, 1.798972e-20, 1.003089e-36, -7.709882e-21, 0, -1.28498e-20, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 0, -1.28498e-20, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 0, 
    -5.139921e-21, -1.027984e-20, -1.003089e-36, 1.027984e-20, -1.28498e-20, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, -1.28498e-20, -1.28498e-20, 
    1.28498e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    1.28498e-20, -1.027984e-20, -1.541976e-20, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, 5.139921e-21, -5.139921e-21, 
    1.003089e-36, 2.569961e-21, 7.709882e-21, 0, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 0, 
    1.027984e-20, -1.003089e-36, -1.28498e-20, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, 0, 0, -7.709882e-21, 0, 5.139921e-21, -7.709882e-21, 0, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    0, 0, 5.139921e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    7.709882e-21, 0, -2.569961e-21, -5.139921e-21, -1.541976e-20, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 0, 1.027984e-20, 7.709882e-21, 
    -1.003089e-36, 7.709882e-21, 1.541976e-20, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, 0, 1.027984e-20, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, 1.003089e-36, 2.569961e-21, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 0,
  5.139921e-21, -1.798972e-20, 2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -1.28498e-20, -7.709882e-21, 0, -2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -1.027984e-20, 7.709882e-21, 0, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -1.541976e-20, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, -1.28498e-20, -1.027984e-20, 
    -1.541976e-20, 1.003089e-36, -2.569961e-21, -1.541976e-20, -1.541976e-20, 
    1.003089e-36, -2.569961e-21, 5.139921e-21, -7.709882e-21, 1.003089e-36, 
    0, 7.709882e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 0, 
    -1.798972e-20, 5.139921e-21, 1.798972e-20, 7.709882e-21, -2.569961e-21, 
    -1.28498e-20, -7.709882e-21, 1.28498e-20, -5.139921e-21, 0, 1.003089e-36, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 1.28498e-20, 1.28498e-20, 
    1.28498e-20, 7.709882e-21, -1.541976e-20, 7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, 
    5.139921e-21, -1.28498e-20, 1.027984e-20, 1.027984e-20, -1.003089e-36, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, -1.003089e-36, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -2.055969e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, -5.139921e-21, 
    1.027984e-20, 7.709882e-21, 0, 1.027984e-20, 1.28498e-20, -1.541976e-20, 
    -1.003089e-36, -5.139921e-21, 7.709882e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, 0, 0, 7.709882e-21, 1.003089e-36, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 1.798972e-20, -1.003089e-36, 
    -1.541976e-20, -7.709882e-21, -1.541976e-20, 1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    1.541976e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 0, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 0, 2.569961e-21, 
    -1.003089e-36, -5.139921e-21, 1.003089e-36, 1.003089e-36, -5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -1.003089e-36, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -2.312965e-20, -2.569961e-21, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 1.541976e-20, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 0, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 0, 1.027984e-20, 5.139921e-21, 1.541976e-20, 0, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, 1.28498e-20, 
    2.569961e-21, 7.709882e-21, 0, 1.003089e-36, 0, -2.569961e-21, 
    -1.28498e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, 0, 
    5.139921e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, -1.541976e-20, 
    1.28498e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, 1.28498e-20, 
    1.28498e-20, -5.139921e-21, 1.003089e-36, -1.027984e-20, 7.709882e-21, 
    7.709882e-21, -1.541976e-20, 1.541976e-20, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -1.027984e-20, 0, -7.709882e-21, -1.28498e-20, 
    -7.709882e-21, 5.139921e-21, 2.055969e-20, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, 7.709882e-21, -1.027984e-20, 0, -1.027984e-20, 
    7.709882e-21, 1.003089e-36, -1.541976e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21,
  -7.709882e-21, -1.798972e-20, -1.027984e-20, 1.027984e-20, -7.709882e-21, 
    1.027984e-20, -2.055969e-20, 7.709882e-21, -7.709882e-21, 1.027984e-20, 
    1.28498e-20, 1.003089e-36, 2.569961e-21, -1.28498e-20, 2.569961e-21, 
    1.003089e-36, 1.027984e-20, -7.709882e-21, -7.709882e-21, 1.28498e-20, 
    1.28498e-20, 1.027984e-20, -7.709882e-21, 0, 0, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 0, 
    -1.027984e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 1.541976e-20, 
    -5.139921e-21, 7.709882e-21, 7.709882e-21, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, 1.28498e-20, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, -1.003089e-36, 
    5.139921e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.003089e-36, -1.003089e-36, 2.569961e-21, -2.569961e-21, -1.003089e-36, 
    -5.139921e-21, -1.003089e-36, -7.709882e-21, 0, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 0, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    1.003089e-36, 0, 7.709882e-21, -1.027984e-20, -7.709882e-21, 0, 
    1.027984e-20, -1.28498e-20, -1.28498e-20, 1.027984e-20, 0, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, -1.003089e-36, -1.798972e-20, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 0, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -1.28498e-20, -7.709882e-21, 1.541976e-20, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 0, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, 0, -7.709882e-21, 1.027984e-20, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -2.569961e-21, -1.003089e-36, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 1.541976e-20, -1.003089e-36, -2.569961e-21, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -2.569961e-21, -2.569961e-21, 1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 1.003089e-36, 
    -1.798972e-20, -2.569961e-21, -1.027984e-20, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    2.055969e-20, -1.027984e-20, 2.569961e-21, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -1.541976e-20, -1.28498e-20, -7.709882e-21, 1.027984e-20, 
    -1.003089e-36, -1.027984e-20, 2.569961e-21, 1.28498e-20, 1.003089e-36, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, 1.28498e-20, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.28498e-20, 1.541976e-20, 5.139921e-21, 2.569961e-21, 1.541976e-20, 
    1.027984e-20, 7.709882e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    1.003089e-36, 1.003089e-36, -2.312965e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, 1.28498e-20, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -1.28498e-20, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    1.027984e-20, 1.28498e-20, 5.139921e-21, -5.139921e-21, -1.003089e-36, 
    7.709882e-21, 1.027984e-20, -1.027984e-20, -2.569961e-21, 1.541976e-20, 
    5.139921e-21, 7.709882e-21, -1.28498e-20, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, 1.541976e-20, 1.798972e-20, 2.569961e-21, 1.28498e-20, 
    1.541976e-20, -1.027984e-20, -2.569961e-21, 1.027984e-20, 7.709882e-21, 
    7.709882e-21, -1.541976e-20, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 1.003089e-36, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, -7.709882e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, 1.798972e-20, -1.541976e-20, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 7.709882e-21, 1.541976e-20, -2.569961e-21, 1.28498e-20, 
    1.003089e-36, 1.28498e-20, 0, 1.28498e-20, 2.569961e-21, -2.055969e-20, 
    -1.798972e-20, 1.027984e-20, -2.569961e-21, 1.28498e-20,
  -1.28498e-20, 1.28498e-20, -1.541976e-20, -5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, 
    1.28498e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -2.312965e-20, 1.027984e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 1.541976e-20, -7.709882e-21, 1.28498e-20, 1.541976e-20, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, 1.003089e-36, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    1.798972e-20, 2.569961e-21, 1.28498e-20, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, -7.709882e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, -1.541976e-20, -7.709882e-21, -1.027984e-20, 1.027984e-20, 
    0, 2.569961e-20, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, 1.28498e-20, -7.709882e-21, -7.709882e-21, 1.541976e-20, 
    5.139921e-21, 2.826957e-20, 1.027984e-20, 1.798972e-20, 5.139921e-21, 
    -1.003089e-36, -5.139921e-21, 1.798972e-20, 2.569961e-21, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, -1.798972e-20, 
    1.541976e-20, 1.28498e-20, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    2.826957e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -1.541976e-20, -5.139921e-21, -1.003089e-36, -1.28498e-20, 1.798972e-20, 
    -5.139921e-21, 1.28498e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, 
    1.027984e-20, -2.055969e-20, 0, -7.709882e-21, 2.312965e-20, 
    1.541976e-20, -2.569961e-21, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 1.28498e-20, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 1.28498e-20, 2.055969e-20, 
    -2.569961e-21, -7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.055969e-20, 7.709882e-21, 
    -2.055969e-20, -2.569961e-21, 7.709882e-21, 1.541976e-20, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, -1.003089e-36, 2.312965e-20, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, -7.709882e-21, -1.28498e-20, 
    2.569961e-21, 1.003089e-36, -1.541976e-20, 1.541976e-20, 1.003089e-36, 
    -2.569961e-21, -1.798972e-20, -1.003089e-36, 1.541976e-20, 1.027984e-20, 
    7.709882e-21, -1.28498e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, -1.003089e-36, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, -2.569961e-21, 
    1.28498e-20, 1.541976e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, -2.569961e-21, -3.083953e-20, 1.541976e-20, -1.28498e-20, 
    5.139921e-21, -1.28498e-20, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, -1.28498e-20, -1.798972e-20, 7.709882e-21, 2.055969e-20, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, 1.28498e-20, -5.139921e-21, 
    -1.798972e-20, -7.709882e-21, -1.28498e-20, -7.709882e-21, -2.055969e-20, 
    -5.139921e-21, -1.28498e-20, 1.003089e-36, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -1.798972e-20, -1.798972e-20, 
    7.709882e-21, -7.709882e-21, -1.003089e-36, -2.569961e-21, 1.798972e-20, 
    -1.027984e-20, 1.003089e-36, -1.541976e-20, -1.28498e-20, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -7.709882e-21, 1.798972e-20, 
    -2.569961e-21, 3.083953e-20, 1.541976e-20, 1.027984e-20, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, 0, -1.28498e-20, 
    -1.003089e-36, -5.139921e-21, -2.569961e-21, 0, -5.139921e-21, 
    2.312965e-20, 1.798972e-20, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    1.027984e-20, 1.003089e-36, 5.139921e-21, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -1.798972e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, -1.798972e-20, 
    -5.139921e-21, 1.28498e-20, -1.027984e-20, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, -3.340949e-20, -1.003089e-36, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, -1.541976e-20, 
    0, 2.569961e-21, -5.139921e-21, 7.709882e-21, -1.541976e-20, 
    -5.139921e-21, 2.312965e-20, -1.003089e-36, 2.569961e-20, -2.569961e-21, 
    -5.139921e-21, -1.003089e-36, -1.003089e-36, 1.003089e-36, -1.798972e-20, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-20, -2.569961e-21, -1.541976e-20, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.288034e-12, 5.311301e-12, 5.306778e-12, 5.325544e-12, 5.315134e-12, 
    5.327422e-12, 5.292751e-12, 5.312225e-12, 5.299793e-12, 5.290129e-12, 
    5.361963e-12, 5.326381e-12, 5.398921e-12, 5.376229e-12, 5.433232e-12, 
    5.39539e-12, 5.440862e-12, 5.432139e-12, 5.45839e-12, 5.450869e-12, 
    5.484447e-12, 5.461861e-12, 5.501852e-12, 5.479053e-12, 5.48262e-12, 
    5.461116e-12, 5.333541e-12, 5.357534e-12, 5.33212e-12, 5.335541e-12, 
    5.334006e-12, 5.315349e-12, 5.305948e-12, 5.286255e-12, 5.28983e-12, 
    5.304293e-12, 5.33708e-12, 5.32595e-12, 5.353998e-12, 5.353365e-12, 
    5.384592e-12, 5.370512e-12, 5.422995e-12, 5.408079e-12, 5.451183e-12, 
    5.440343e-12, 5.450674e-12, 5.447542e-12, 5.450715e-12, 5.434817e-12, 
    5.441628e-12, 5.427638e-12, 5.373149e-12, 5.389164e-12, 5.341401e-12, 
    5.312682e-12, 5.293605e-12, 5.280068e-12, 5.281982e-12, 5.28563e-12, 
    5.304378e-12, 5.322004e-12, 5.335436e-12, 5.344421e-12, 5.353274e-12, 
    5.380073e-12, 5.394255e-12, 5.426012e-12, 5.420281e-12, 5.42999e-12, 
    5.439264e-12, 5.454837e-12, 5.452274e-12, 5.459135e-12, 5.429733e-12, 
    5.449274e-12, 5.417016e-12, 5.425839e-12, 5.355683e-12, 5.328953e-12, 
    5.317592e-12, 5.307647e-12, 5.283454e-12, 5.300161e-12, 5.293575e-12, 
    5.309244e-12, 5.3192e-12, 5.314276e-12, 5.344667e-12, 5.332852e-12, 
    5.395096e-12, 5.368286e-12, 5.438183e-12, 5.421457e-12, 5.442192e-12, 
    5.431611e-12, 5.449741e-12, 5.433424e-12, 5.461688e-12, 5.467843e-12, 
    5.463637e-12, 5.479792e-12, 5.43252e-12, 5.450675e-12, 5.314138e-12, 
    5.314941e-12, 5.318683e-12, 5.302236e-12, 5.30123e-12, 5.286157e-12, 
    5.299569e-12, 5.30528e-12, 5.319777e-12, 5.328353e-12, 5.336504e-12, 
    5.354427e-12, 5.374444e-12, 5.402434e-12, 5.422541e-12, 5.43602e-12, 
    5.427755e-12, 5.435052e-12, 5.426895e-12, 5.423071e-12, 5.465537e-12, 
    5.441692e-12, 5.477468e-12, 5.475489e-12, 5.459298e-12, 5.475712e-12, 
    5.315505e-12, 5.310883e-12, 5.294838e-12, 5.307395e-12, 5.284516e-12, 
    5.297323e-12, 5.304687e-12, 5.333099e-12, 5.339341e-12, 5.34513e-12, 
    5.356562e-12, 5.371233e-12, 5.39697e-12, 5.419362e-12, 5.439804e-12, 
    5.438306e-12, 5.438834e-12, 5.443401e-12, 5.432089e-12, 5.445258e-12, 
    5.447468e-12, 5.441689e-12, 5.475224e-12, 5.465643e-12, 5.475446e-12, 
    5.469209e-12, 5.312386e-12, 5.320162e-12, 5.31596e-12, 5.323862e-12, 
    5.318295e-12, 5.343049e-12, 5.350471e-12, 5.385197e-12, 5.370944e-12, 
    5.393626e-12, 5.373248e-12, 5.376859e-12, 5.394367e-12, 5.374349e-12, 
    5.418129e-12, 5.388448e-12, 5.443578e-12, 5.413941e-12, 5.445435e-12, 
    5.439716e-12, 5.449185e-12, 5.457666e-12, 5.468335e-12, 5.488023e-12, 
    5.483464e-12, 5.499927e-12, 5.331755e-12, 5.341842e-12, 5.340953e-12, 
    5.351509e-12, 5.359315e-12, 5.376234e-12, 5.40337e-12, 5.393166e-12, 
    5.4119e-12, 5.415661e-12, 5.387199e-12, 5.404675e-12, 5.348592e-12, 
    5.357654e-12, 5.352258e-12, 5.332551e-12, 5.395518e-12, 5.363204e-12, 
    5.422874e-12, 5.405368e-12, 5.456457e-12, 5.43105e-12, 5.480954e-12, 
    5.502289e-12, 5.522366e-12, 5.545831e-12, 5.347346e-12, 5.340492e-12, 
    5.352764e-12, 5.369742e-12, 5.385494e-12, 5.406436e-12, 5.408579e-12, 
    5.412502e-12, 5.422664e-12, 5.431208e-12, 5.413743e-12, 5.43335e-12, 
    5.359756e-12, 5.398323e-12, 5.337902e-12, 5.356097e-12, 5.368741e-12, 
    5.363194e-12, 5.392e-12, 5.398789e-12, 5.426378e-12, 5.412116e-12, 
    5.497023e-12, 5.459458e-12, 5.563695e-12, 5.534566e-12, 5.338098e-12, 
    5.347322e-12, 5.379426e-12, 5.364151e-12, 5.407834e-12, 5.418586e-12, 
    5.427327e-12, 5.4385e-12, 5.439706e-12, 5.446327e-12, 5.435478e-12, 
    5.445898e-12, 5.406481e-12, 5.424095e-12, 5.375756e-12, 5.387522e-12, 
    5.382109e-12, 5.376172e-12, 5.394496e-12, 5.414018e-12, 5.414434e-12, 
    5.420694e-12, 5.438335e-12, 5.408011e-12, 5.501873e-12, 5.443907e-12, 
    5.357381e-12, 5.375149e-12, 5.377686e-12, 5.370803e-12, 5.417508e-12, 
    5.400586e-12, 5.446165e-12, 5.433847e-12, 5.45403e-12, 5.444001e-12, 
    5.442525e-12, 5.429643e-12, 5.421624e-12, 5.401362e-12, 5.384875e-12, 
    5.371802e-12, 5.374842e-12, 5.389203e-12, 5.415212e-12, 5.439816e-12, 
    5.434426e-12, 5.452497e-12, 5.404666e-12, 5.424723e-12, 5.416972e-12, 
    5.437183e-12, 5.392895e-12, 5.430611e-12, 5.383255e-12, 5.387407e-12, 
    5.40025e-12, 5.426084e-12, 5.431798e-12, 5.437901e-12, 5.434135e-12, 
    5.415872e-12, 5.412879e-12, 5.399937e-12, 5.396364e-12, 5.386502e-12, 
    5.378338e-12, 5.385798e-12, 5.393632e-12, 5.41588e-12, 5.435929e-12, 
    5.457787e-12, 5.463136e-12, 5.488678e-12, 5.467887e-12, 5.502196e-12, 
    5.473028e-12, 5.523519e-12, 5.432796e-12, 5.472169e-12, 5.400834e-12, 
    5.408519e-12, 5.422419e-12, 5.4543e-12, 5.437088e-12, 5.457217e-12, 
    5.412762e-12, 5.389699e-12, 5.38373e-12, 5.372596e-12, 5.383985e-12, 
    5.383059e-12, 5.393956e-12, 5.390454e-12, 5.416618e-12, 5.402564e-12, 
    5.442488e-12, 5.457058e-12, 5.498202e-12, 5.523425e-12, 5.549099e-12, 
    5.560434e-12, 5.563884e-12, 5.565326e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.199261e-11, 3.213337e-11, 3.210601e-11, 3.221954e-11, 3.215656e-11, 
    3.223091e-11, 3.202114e-11, 3.213896e-11, 3.206375e-11, 3.200528e-11, 
    3.243988e-11, 3.22246e-11, 3.266347e-11, 3.252618e-11, 3.287105e-11, 
    3.264211e-11, 3.291721e-11, 3.286444e-11, 3.302326e-11, 3.297776e-11, 
    3.318091e-11, 3.304426e-11, 3.32862e-11, 3.314827e-11, 3.316985e-11, 
    3.303975e-11, 3.226792e-11, 3.241308e-11, 3.225933e-11, 3.228003e-11, 
    3.227074e-11, 3.215786e-11, 3.210098e-11, 3.198184e-11, 3.200347e-11, 
    3.209098e-11, 3.228933e-11, 3.2222e-11, 3.239169e-11, 3.238786e-11, 
    3.257678e-11, 3.24916e-11, 3.280912e-11, 3.271888e-11, 3.297966e-11, 
    3.291408e-11, 3.297658e-11, 3.295763e-11, 3.297683e-11, 3.288064e-11, 
    3.292185e-11, 3.283721e-11, 3.250755e-11, 3.260444e-11, 3.231548e-11, 
    3.214173e-11, 3.202631e-11, 3.194441e-11, 3.195599e-11, 3.197807e-11, 
    3.209149e-11, 3.219812e-11, 3.227939e-11, 3.233375e-11, 3.238731e-11, 
    3.254944e-11, 3.263525e-11, 3.282737e-11, 3.27927e-11, 3.285144e-11, 
    3.290755e-11, 3.300176e-11, 3.298626e-11, 3.302776e-11, 3.284989e-11, 
    3.296811e-11, 3.277295e-11, 3.282632e-11, 3.240188e-11, 3.224016e-11, 
    3.217144e-11, 3.211127e-11, 3.19649e-11, 3.206598e-11, 3.202613e-11, 
    3.212092e-11, 3.218116e-11, 3.215137e-11, 3.233524e-11, 3.226375e-11, 
    3.264033e-11, 3.247813e-11, 3.290101e-11, 3.279981e-11, 3.292526e-11, 
    3.286125e-11, 3.297093e-11, 3.287222e-11, 3.304321e-11, 3.308045e-11, 
    3.3055e-11, 3.315274e-11, 3.286674e-11, 3.297658e-11, 3.215054e-11, 
    3.215539e-11, 3.217803e-11, 3.207853e-11, 3.207244e-11, 3.198125e-11, 
    3.206239e-11, 3.209694e-11, 3.218465e-11, 3.223653e-11, 3.228585e-11, 
    3.239429e-11, 3.251539e-11, 3.268472e-11, 3.280637e-11, 3.288792e-11, 
    3.283792e-11, 3.288206e-11, 3.283271e-11, 3.280958e-11, 3.30665e-11, 
    3.292224e-11, 3.313869e-11, 3.312671e-11, 3.302875e-11, 3.312806e-11, 
    3.215881e-11, 3.213084e-11, 3.203377e-11, 3.210974e-11, 3.197132e-11, 
    3.20488e-11, 3.209336e-11, 3.226525e-11, 3.230301e-11, 3.233804e-11, 
    3.24072e-11, 3.249596e-11, 3.265167e-11, 3.278714e-11, 3.291082e-11, 
    3.290175e-11, 3.290494e-11, 3.293257e-11, 3.286414e-11, 3.294381e-11, 
    3.295718e-11, 3.292222e-11, 3.31251e-11, 3.306714e-11, 3.312645e-11, 
    3.308871e-11, 3.213993e-11, 3.218698e-11, 3.216156e-11, 3.220936e-11, 
    3.217569e-11, 3.232544e-11, 3.237035e-11, 3.258044e-11, 3.249421e-11, 
    3.263144e-11, 3.250815e-11, 3.253e-11, 3.263592e-11, 3.251481e-11, 
    3.277968e-11, 3.260011e-11, 3.293365e-11, 3.275434e-11, 3.294488e-11, 
    3.291028e-11, 3.296757e-11, 3.301888e-11, 3.308343e-11, 3.320254e-11, 
    3.317496e-11, 3.327456e-11, 3.225712e-11, 3.231814e-11, 3.231277e-11, 
    3.237663e-11, 3.242386e-11, 3.252622e-11, 3.269039e-11, 3.262865e-11, 
    3.274199e-11, 3.276475e-11, 3.259256e-11, 3.269828e-11, 3.235898e-11, 
    3.24138e-11, 3.238116e-11, 3.226193e-11, 3.264288e-11, 3.244738e-11, 
    3.280838e-11, 3.270248e-11, 3.301157e-11, 3.285785e-11, 3.315977e-11, 
    3.328885e-11, 3.341031e-11, 3.355228e-11, 3.235144e-11, 3.230998e-11, 
    3.238422e-11, 3.248694e-11, 3.258224e-11, 3.270894e-11, 3.27219e-11, 
    3.274564e-11, 3.280711e-11, 3.285881e-11, 3.275314e-11, 3.287177e-11, 
    3.242652e-11, 3.265985e-11, 3.229431e-11, 3.240438e-11, 3.248088e-11, 
    3.244732e-11, 3.26216e-11, 3.266267e-11, 3.282959e-11, 3.27433e-11, 
    3.325699e-11, 3.302972e-11, 3.366036e-11, 3.348413e-11, 3.229549e-11, 
    3.23513e-11, 3.254553e-11, 3.245312e-11, 3.271739e-11, 3.278245e-11, 
    3.283532e-11, 3.290293e-11, 3.291022e-11, 3.295028e-11, 3.288464e-11, 
    3.294768e-11, 3.270921e-11, 3.281578e-11, 3.252332e-11, 3.259451e-11, 
    3.256176e-11, 3.252584e-11, 3.26367e-11, 3.275481e-11, 3.275733e-11, 
    3.27952e-11, 3.290193e-11, 3.271847e-11, 3.328634e-11, 3.293564e-11, 
    3.241215e-11, 3.251965e-11, 3.2535e-11, 3.249336e-11, 3.277592e-11, 
    3.267354e-11, 3.29493e-11, 3.287477e-11, 3.299688e-11, 3.293621e-11, 
    3.292728e-11, 3.284934e-11, 3.280082e-11, 3.267824e-11, 3.25785e-11, 
    3.24994e-11, 3.251779e-11, 3.260468e-11, 3.276203e-11, 3.291089e-11, 
    3.287828e-11, 3.298761e-11, 3.269823e-11, 3.281957e-11, 3.277268e-11, 
    3.289496e-11, 3.262702e-11, 3.28552e-11, 3.256869e-11, 3.259381e-11, 
    3.267151e-11, 3.282781e-11, 3.286238e-11, 3.28993e-11, 3.287652e-11, 
    3.276603e-11, 3.274792e-11, 3.266962e-11, 3.264801e-11, 3.258834e-11, 
    3.253895e-11, 3.258408e-11, 3.263147e-11, 3.276607e-11, 3.288737e-11, 
    3.301961e-11, 3.305197e-11, 3.32065e-11, 3.308072e-11, 3.328829e-11, 
    3.311182e-11, 3.341729e-11, 3.286841e-11, 3.310662e-11, 3.267504e-11, 
    3.272154e-11, 3.280564e-11, 3.299852e-11, 3.289438e-11, 3.301616e-11, 
    3.274721e-11, 3.260768e-11, 3.257157e-11, 3.250421e-11, 3.257311e-11, 
    3.25675e-11, 3.263343e-11, 3.261225e-11, 3.277054e-11, 3.268551e-11, 
    3.292705e-11, 3.30152e-11, 3.326412e-11, 3.341672e-11, 3.357205e-11, 
    3.364063e-11, 3.36615e-11, 3.367022e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.356944e-08, 6.384899e-08, 6.379465e-08, 6.402013e-08, 6.389505e-08, 
    6.404269e-08, 6.362611e-08, 6.38601e-08, 6.371073e-08, 6.359461e-08, 
    6.445772e-08, 6.403019e-08, 6.490177e-08, 6.462912e-08, 6.531402e-08, 
    6.485934e-08, 6.540569e-08, 6.53009e-08, 6.56163e-08, 6.552594e-08, 
    6.592938e-08, 6.565801e-08, 6.61385e-08, 6.586457e-08, 6.590742e-08, 
    6.564905e-08, 6.411622e-08, 6.44045e-08, 6.409914e-08, 6.414025e-08, 
    6.41218e-08, 6.389764e-08, 6.378468e-08, 6.354806e-08, 6.359102e-08, 
    6.376479e-08, 6.415873e-08, 6.4025e-08, 6.436202e-08, 6.435441e-08, 
    6.47296e-08, 6.456043e-08, 6.519103e-08, 6.50118e-08, 6.552971e-08, 
    6.539947e-08, 6.552359e-08, 6.548596e-08, 6.552408e-08, 6.533306e-08, 
    6.541491e-08, 6.524682e-08, 6.459211e-08, 6.478453e-08, 6.421065e-08, 
    6.386559e-08, 6.363638e-08, 6.347373e-08, 6.349672e-08, 6.354056e-08, 
    6.376582e-08, 6.397759e-08, 6.413898e-08, 6.424694e-08, 6.435332e-08, 
    6.467531e-08, 6.484571e-08, 6.522728e-08, 6.515841e-08, 6.527507e-08, 
    6.538651e-08, 6.557362e-08, 6.554281e-08, 6.562525e-08, 6.527198e-08, 
    6.550677e-08, 6.511919e-08, 6.522519e-08, 6.438226e-08, 6.406108e-08, 
    6.392459e-08, 6.38051e-08, 6.351441e-08, 6.371515e-08, 6.363602e-08, 
    6.382428e-08, 6.394391e-08, 6.388474e-08, 6.42499e-08, 6.410793e-08, 
    6.485581e-08, 6.453368e-08, 6.537351e-08, 6.517254e-08, 6.542168e-08, 
    6.529455e-08, 6.551238e-08, 6.531634e-08, 6.565593e-08, 6.572988e-08, 
    6.567934e-08, 6.587345e-08, 6.530546e-08, 6.55236e-08, 6.388309e-08, 
    6.389273e-08, 6.393769e-08, 6.374008e-08, 6.372799e-08, 6.354689e-08, 
    6.370803e-08, 6.377665e-08, 6.395084e-08, 6.405388e-08, 6.415182e-08, 
    6.436717e-08, 6.460768e-08, 6.494398e-08, 6.518557e-08, 6.534752e-08, 
    6.524822e-08, 6.533589e-08, 6.523788e-08, 6.519194e-08, 6.570217e-08, 
    6.541567e-08, 6.584553e-08, 6.582174e-08, 6.562721e-08, 6.582443e-08, 
    6.389951e-08, 6.384398e-08, 6.365119e-08, 6.380206e-08, 6.352717e-08, 
    6.368104e-08, 6.376953e-08, 6.411091e-08, 6.41859e-08, 6.425545e-08, 
    6.439281e-08, 6.456909e-08, 6.487833e-08, 6.514738e-08, 6.539299e-08, 
    6.537499e-08, 6.538133e-08, 6.54362e-08, 6.530028e-08, 6.545852e-08, 
    6.548507e-08, 6.541563e-08, 6.581856e-08, 6.570345e-08, 6.582124e-08, 
    6.574629e-08, 6.386203e-08, 6.395546e-08, 6.390498e-08, 6.399992e-08, 
    6.393303e-08, 6.423046e-08, 6.431962e-08, 6.473687e-08, 6.456563e-08, 
    6.483815e-08, 6.45933e-08, 6.463669e-08, 6.484705e-08, 6.460653e-08, 
    6.513255e-08, 6.477594e-08, 6.543834e-08, 6.508223e-08, 6.546065e-08, 
    6.539193e-08, 6.55057e-08, 6.560761e-08, 6.57358e-08, 6.597234e-08, 
    6.591757e-08, 6.611538e-08, 6.409476e-08, 6.421595e-08, 6.420527e-08, 
    6.43321e-08, 6.44259e-08, 6.462918e-08, 6.495523e-08, 6.483262e-08, 
    6.505771e-08, 6.51029e-08, 6.476093e-08, 6.49709e-08, 6.429705e-08, 
    6.440593e-08, 6.43411e-08, 6.410432e-08, 6.486088e-08, 6.447262e-08, 
    6.518957e-08, 6.497923e-08, 6.559308e-08, 6.528781e-08, 6.588741e-08, 
    6.614376e-08, 6.638498e-08, 6.666692e-08, 6.428208e-08, 6.419974e-08, 
    6.434718e-08, 6.455118e-08, 6.474044e-08, 6.499207e-08, 6.501781e-08, 
    6.506495e-08, 6.518705e-08, 6.52897e-08, 6.507986e-08, 6.531544e-08, 
    6.443119e-08, 6.489459e-08, 6.416861e-08, 6.438723e-08, 6.453915e-08, 
    6.44725e-08, 6.481861e-08, 6.490018e-08, 6.523167e-08, 6.506031e-08, 
    6.60805e-08, 6.562914e-08, 6.688157e-08, 6.653157e-08, 6.417097e-08, 
    6.42818e-08, 6.466754e-08, 6.448401e-08, 6.500886e-08, 6.513805e-08, 
    6.524307e-08, 6.537733e-08, 6.539182e-08, 6.547136e-08, 6.534101e-08, 
    6.546621e-08, 6.49926e-08, 6.520425e-08, 6.462344e-08, 6.476481e-08, 
    6.469977e-08, 6.462844e-08, 6.48486e-08, 6.508316e-08, 6.508817e-08, 
    6.516338e-08, 6.537534e-08, 6.501099e-08, 6.613876e-08, 6.544229e-08, 
    6.440266e-08, 6.461615e-08, 6.464663e-08, 6.456393e-08, 6.51251e-08, 
    6.492177e-08, 6.546942e-08, 6.532141e-08, 6.556392e-08, 6.544342e-08, 
    6.542568e-08, 6.52709e-08, 6.517455e-08, 6.493109e-08, 6.473301e-08, 
    6.457592e-08, 6.461245e-08, 6.4785e-08, 6.509751e-08, 6.539313e-08, 
    6.532837e-08, 6.554549e-08, 6.497081e-08, 6.521179e-08, 6.511865e-08, 
    6.53615e-08, 6.482936e-08, 6.528253e-08, 6.471353e-08, 6.476342e-08, 
    6.491774e-08, 6.522814e-08, 6.52968e-08, 6.537012e-08, 6.532488e-08, 
    6.510544e-08, 6.506949e-08, 6.491398e-08, 6.487105e-08, 6.475256e-08, 
    6.465446e-08, 6.474409e-08, 6.483822e-08, 6.510553e-08, 6.534642e-08, 
    6.560906e-08, 6.567333e-08, 6.598021e-08, 6.57304e-08, 6.614265e-08, 
    6.579219e-08, 6.639884e-08, 6.530878e-08, 6.578186e-08, 6.492476e-08, 
    6.501709e-08, 6.518411e-08, 6.556716e-08, 6.536035e-08, 6.560221e-08, 
    6.506808e-08, 6.479096e-08, 6.471925e-08, 6.458548e-08, 6.472231e-08, 
    6.471118e-08, 6.484211e-08, 6.480003e-08, 6.511441e-08, 6.494554e-08, 
    6.542524e-08, 6.56003e-08, 6.609465e-08, 6.639771e-08, 6.670619e-08, 
    6.684238e-08, 6.688383e-08, 6.690116e-08 ;

 SOILC_LOSS =
  6.356944e-08, 6.384899e-08, 6.379465e-08, 6.402013e-08, 6.389505e-08, 
    6.404269e-08, 6.362611e-08, 6.38601e-08, 6.371073e-08, 6.359461e-08, 
    6.445772e-08, 6.403019e-08, 6.490177e-08, 6.462912e-08, 6.531402e-08, 
    6.485934e-08, 6.540569e-08, 6.53009e-08, 6.56163e-08, 6.552594e-08, 
    6.592938e-08, 6.565801e-08, 6.61385e-08, 6.586457e-08, 6.590742e-08, 
    6.564905e-08, 6.411622e-08, 6.44045e-08, 6.409914e-08, 6.414025e-08, 
    6.41218e-08, 6.389764e-08, 6.378468e-08, 6.354806e-08, 6.359102e-08, 
    6.376479e-08, 6.415873e-08, 6.4025e-08, 6.436202e-08, 6.435441e-08, 
    6.47296e-08, 6.456043e-08, 6.519103e-08, 6.50118e-08, 6.552971e-08, 
    6.539947e-08, 6.552359e-08, 6.548596e-08, 6.552408e-08, 6.533306e-08, 
    6.541491e-08, 6.524682e-08, 6.459211e-08, 6.478453e-08, 6.421065e-08, 
    6.386559e-08, 6.363638e-08, 6.347373e-08, 6.349672e-08, 6.354056e-08, 
    6.376582e-08, 6.397759e-08, 6.413898e-08, 6.424694e-08, 6.435332e-08, 
    6.467531e-08, 6.484571e-08, 6.522728e-08, 6.515841e-08, 6.527507e-08, 
    6.538651e-08, 6.557362e-08, 6.554281e-08, 6.562525e-08, 6.527198e-08, 
    6.550677e-08, 6.511919e-08, 6.522519e-08, 6.438226e-08, 6.406108e-08, 
    6.392459e-08, 6.38051e-08, 6.351441e-08, 6.371515e-08, 6.363602e-08, 
    6.382428e-08, 6.394391e-08, 6.388474e-08, 6.42499e-08, 6.410793e-08, 
    6.485581e-08, 6.453368e-08, 6.537351e-08, 6.517254e-08, 6.542168e-08, 
    6.529455e-08, 6.551238e-08, 6.531634e-08, 6.565593e-08, 6.572988e-08, 
    6.567934e-08, 6.587345e-08, 6.530546e-08, 6.55236e-08, 6.388309e-08, 
    6.389273e-08, 6.393769e-08, 6.374008e-08, 6.372799e-08, 6.354689e-08, 
    6.370803e-08, 6.377665e-08, 6.395084e-08, 6.405388e-08, 6.415182e-08, 
    6.436717e-08, 6.460768e-08, 6.494398e-08, 6.518557e-08, 6.534752e-08, 
    6.524822e-08, 6.533589e-08, 6.523788e-08, 6.519194e-08, 6.570217e-08, 
    6.541567e-08, 6.584553e-08, 6.582174e-08, 6.562721e-08, 6.582443e-08, 
    6.389951e-08, 6.384398e-08, 6.365119e-08, 6.380206e-08, 6.352717e-08, 
    6.368104e-08, 6.376953e-08, 6.411091e-08, 6.41859e-08, 6.425545e-08, 
    6.439281e-08, 6.456909e-08, 6.487833e-08, 6.514738e-08, 6.539299e-08, 
    6.537499e-08, 6.538133e-08, 6.54362e-08, 6.530028e-08, 6.545852e-08, 
    6.548507e-08, 6.541563e-08, 6.581856e-08, 6.570345e-08, 6.582124e-08, 
    6.574629e-08, 6.386203e-08, 6.395546e-08, 6.390498e-08, 6.399992e-08, 
    6.393303e-08, 6.423046e-08, 6.431962e-08, 6.473687e-08, 6.456563e-08, 
    6.483815e-08, 6.45933e-08, 6.463669e-08, 6.484705e-08, 6.460653e-08, 
    6.513255e-08, 6.477594e-08, 6.543834e-08, 6.508223e-08, 6.546065e-08, 
    6.539193e-08, 6.55057e-08, 6.560761e-08, 6.57358e-08, 6.597234e-08, 
    6.591757e-08, 6.611538e-08, 6.409476e-08, 6.421595e-08, 6.420527e-08, 
    6.43321e-08, 6.44259e-08, 6.462918e-08, 6.495523e-08, 6.483262e-08, 
    6.505771e-08, 6.51029e-08, 6.476093e-08, 6.49709e-08, 6.429705e-08, 
    6.440593e-08, 6.43411e-08, 6.410432e-08, 6.486088e-08, 6.447262e-08, 
    6.518957e-08, 6.497923e-08, 6.559308e-08, 6.528781e-08, 6.588741e-08, 
    6.614376e-08, 6.638498e-08, 6.666692e-08, 6.428208e-08, 6.419974e-08, 
    6.434718e-08, 6.455118e-08, 6.474044e-08, 6.499207e-08, 6.501781e-08, 
    6.506495e-08, 6.518705e-08, 6.52897e-08, 6.507986e-08, 6.531544e-08, 
    6.443119e-08, 6.489459e-08, 6.416861e-08, 6.438723e-08, 6.453915e-08, 
    6.44725e-08, 6.481861e-08, 6.490018e-08, 6.523167e-08, 6.506031e-08, 
    6.60805e-08, 6.562914e-08, 6.688157e-08, 6.653157e-08, 6.417097e-08, 
    6.42818e-08, 6.466754e-08, 6.448401e-08, 6.500886e-08, 6.513805e-08, 
    6.524307e-08, 6.537733e-08, 6.539182e-08, 6.547136e-08, 6.534101e-08, 
    6.546621e-08, 6.49926e-08, 6.520425e-08, 6.462344e-08, 6.476481e-08, 
    6.469977e-08, 6.462844e-08, 6.48486e-08, 6.508316e-08, 6.508817e-08, 
    6.516338e-08, 6.537534e-08, 6.501099e-08, 6.613876e-08, 6.544229e-08, 
    6.440266e-08, 6.461615e-08, 6.464663e-08, 6.456393e-08, 6.51251e-08, 
    6.492177e-08, 6.546942e-08, 6.532141e-08, 6.556392e-08, 6.544342e-08, 
    6.542568e-08, 6.52709e-08, 6.517455e-08, 6.493109e-08, 6.473301e-08, 
    6.457592e-08, 6.461245e-08, 6.4785e-08, 6.509751e-08, 6.539313e-08, 
    6.532837e-08, 6.554549e-08, 6.497081e-08, 6.521179e-08, 6.511865e-08, 
    6.53615e-08, 6.482936e-08, 6.528253e-08, 6.471353e-08, 6.476342e-08, 
    6.491774e-08, 6.522814e-08, 6.52968e-08, 6.537012e-08, 6.532488e-08, 
    6.510544e-08, 6.506949e-08, 6.491398e-08, 6.487105e-08, 6.475256e-08, 
    6.465446e-08, 6.474409e-08, 6.483822e-08, 6.510553e-08, 6.534642e-08, 
    6.560906e-08, 6.567333e-08, 6.598021e-08, 6.57304e-08, 6.614265e-08, 
    6.579219e-08, 6.639884e-08, 6.530878e-08, 6.578186e-08, 6.492476e-08, 
    6.501709e-08, 6.518411e-08, 6.556716e-08, 6.536035e-08, 6.560221e-08, 
    6.506808e-08, 6.479096e-08, 6.471925e-08, 6.458548e-08, 6.472231e-08, 
    6.471118e-08, 6.484211e-08, 6.480003e-08, 6.511441e-08, 6.494554e-08, 
    6.542524e-08, 6.56003e-08, 6.609465e-08, 6.639771e-08, 6.670619e-08, 
    6.684238e-08, 6.688383e-08, 6.690116e-08 ;

 SOILICE =
  57.49552, 57.6865, 57.64934, 57.80369, 57.71803, 57.81916, 57.5342, 
    57.6941, 57.59198, 57.5127, 58.10423, 57.81059, 58.41063, 58.22237, 
    58.69618, 58.38129, 58.75983, 58.68709, 58.9063, 58.84343, 59.12453, 
    58.93533, 59.27069, 59.07931, 59.10921, 58.9291, 57.86959, 58.0676, 
    57.85787, 57.88607, 57.87341, 57.71979, 57.6425, 57.48095, 57.51025, 
    57.62892, 57.89875, 57.80704, 58.03843, 58.0332, 58.29169, 58.17502, 
    58.61089, 58.48677, 58.84605, 58.75552, 58.84179, 58.81562, 58.84213, 
    58.70941, 58.76625, 58.64957, 58.19686, 58.32962, 57.9344, 57.69784, 
    57.5412, 57.43027, 57.44594, 57.47582, 57.62962, 57.77455, 57.88521, 
    57.95933, 58.03244, 58.2542, 58.37188, 58.63601, 58.58829, 58.66916, 
    58.74652, 58.87658, 58.85516, 58.91252, 58.66703, 58.83009, 58.56112, 
    58.63458, 58.0523, 57.83177, 57.73823, 57.65648, 57.45799, 57.595, 
    57.54095, 57.66961, 57.75148, 57.71097, 57.96136, 57.8639, 58.37886, 
    58.15658, 58.7375, 58.59808, 58.77095, 58.68269, 58.83399, 58.69781, 
    58.93388, 58.98539, 58.95018, 59.08551, 58.69026, 58.84179, 57.70984, 
    57.71644, 57.74722, 57.61203, 57.60377, 57.48015, 57.59014, 57.63703, 
    57.75623, 57.82683, 57.89401, 58.04197, 58.20758, 58.43982, 58.60711, 
    58.71945, 58.65055, 58.71138, 58.64338, 58.61153, 58.96608, 58.76677, 
    59.06603, 59.04944, 58.91388, 59.05131, 57.72108, 57.68308, 57.55132, 
    57.65441, 57.4667, 57.5717, 57.63215, 57.86593, 57.91741, 57.96517, 
    58.05961, 58.18099, 58.39443, 58.58064, 58.75103, 58.73853, 58.74293, 
    58.78104, 58.68667, 58.79655, 58.815, 58.76675, 59.04722, 58.96698, 
    59.04909, 58.99683, 57.69543, 57.75939, 57.72482, 57.78984, 57.74403, 
    57.94799, 58.00926, 58.2967, 58.1786, 58.36666, 58.19768, 58.22759, 
    58.37279, 58.2068, 58.57035, 58.32367, 58.78252, 58.53549, 58.79803, 
    58.75029, 58.82935, 58.90024, 58.98952, 59.15454, 59.1163, 59.25453, 
    57.85487, 57.93803, 57.93071, 58.01785, 58.08237, 58.22242, 58.44762, 
    58.36285, 58.51854, 58.54983, 58.31333, 58.45845, 57.99376, 58.06862, 
    58.02404, 57.86142, 58.38237, 58.11452, 58.60987, 58.46423, 58.89013, 
    58.678, 59.09525, 59.27436, 59.44335, 59.64131, 57.98347, 57.92691, 
    58.02822, 58.16863, 58.29918, 58.47311, 58.49092, 58.52355, 58.60814, 
    58.67933, 58.53386, 58.69719, 58.08598, 58.40567, 57.90554, 58.05575, 
    58.16035, 58.11445, 58.35317, 58.40955, 58.63906, 58.52034, 59.23011, 
    58.91521, 59.7924, 59.5462, 57.90716, 57.98328, 58.24886, 58.12237, 
    58.48473, 58.57418, 58.64698, 58.74014, 58.75021, 58.80547, 58.71494, 
    58.8019, 58.47348, 58.62006, 58.21846, 58.316, 58.27111, 58.2219, 
    58.37389, 58.53615, 58.53963, 58.59172, 58.73871, 58.48621, 59.27083, 
    58.78523, 58.06638, 58.21341, 58.23445, 58.17744, 58.5652, 58.42448, 
    58.80413, 58.70133, 58.86984, 58.78606, 58.77374, 58.66629, 58.59947, 
    58.43092, 58.29404, 58.1857, 58.21088, 58.32994, 58.54609, 58.75112, 
    58.70615, 58.85703, 58.4584, 58.62527, 58.56073, 58.72915, 58.3606, 
    58.6743, 58.28061, 58.31505, 58.42168, 58.6366, 58.68425, 58.73514, 
    58.70373, 58.55158, 58.52669, 58.41909, 58.3894, 58.30755, 58.23986, 
    58.3017, 58.36671, 58.55165, 58.71868, 58.90125, 58.946, 59.16002, 
    58.98574, 59.27354, 59.02877, 59.45303, 58.69254, 59.0216, 58.42654, 
    58.49043, 58.60608, 58.87208, 58.72836, 58.89647, 58.52571, 58.33405, 
    58.28456, 58.19228, 58.28667, 58.27899, 58.36941, 58.34034, 58.5578, 
    58.44092, 58.77342, 58.89515, 59.24002, 59.45226, 59.66895, 59.7648, 
    59.79401, 59.80622,
  78.78071, 79.08004, 79.02182, 79.26369, 79.1295, 79.28794, 78.84139, 
    79.09187, 78.93194, 78.80772, 79.73457, 79.27451, 80.2154, 79.92023, 
    80.66348, 80.16932, 80.76344, 80.64936, 80.9935, 80.8948, 81.33589, 
    81.03909, 81.56555, 81.26502, 81.31191, 81.02928, 79.36708, 79.67712, 
    79.3487, 79.39286, 79.37308, 79.13222, 79.01095, 78.75798, 78.80389, 
    78.98977, 79.41272, 79.26905, 79.63186, 79.62366, 80.02898, 79.84602, 
    80.52978, 80.33504, 80.89892, 80.75679, 80.89221, 80.85115, 80.89275, 
    80.68439, 80.7736, 80.5905, 79.88023, 80.08842, 79.46866, 79.0976, 
    78.85233, 78.67854, 78.70309, 78.74988, 78.99086, 79.21812, 79.39162, 
    79.50782, 79.62247, 79.96989, 80.15462, 80.56911, 80.49434, 80.62116, 
    80.74268, 80.94681, 80.91321, 81.00321, 80.61792, 80.87377, 80.45173, 
    80.56697, 79.65311, 79.30782, 79.16094, 79.03298, 78.72196, 78.93661, 
    78.85192, 79.05363, 79.18195, 79.11849, 79.511, 79.35819, 80.16557, 
    79.81702, 80.72849, 80.50969, 80.78102, 80.64251, 80.87992, 80.66623, 
    81.03677, 81.11757, 81.06234, 81.27486, 80.65438, 80.89216, 79.11668, 
    79.12703, 79.17529, 78.96329, 78.95037, 78.75669, 78.92906, 79.00251, 
    79.18943, 79.30006, 79.40539, 79.63735, 79.89697, 80.26128, 80.52386, 
    80.7002, 80.59207, 80.68753, 80.5808, 80.53085, 81.08725, 80.7744, 
    81.24427, 81.21823, 81.00533, 81.22116, 79.1343, 79.07478, 78.86819, 
    79.02982, 78.73563, 78.90012, 78.9948, 79.36126, 79.4421, 79.51694, 
    79.66505, 79.85538, 80.19009, 80.48226, 80.74977, 80.73016, 80.73705, 
    80.79684, 80.64873, 80.82118, 80.85011, 80.77443, 81.21474, 81.08876, 
    81.21767, 81.13564, 79.09413, 79.19437, 79.14018, 79.24207, 79.17023, 
    79.48988, 79.58592, 80.0367, 79.85159, 80.1465, 79.88156, 79.92842, 
    80.1559, 79.8959, 80.46603, 80.07895, 80.79916, 80.4112, 80.82352, 
    80.74861, 80.87272, 80.98394, 81.12415, 81.38316, 81.32315, 81.54024, 
    79.34403, 79.47433, 79.46296, 79.59957, 79.7007, 79.92038, 80.27357, 
    80.14064, 80.38491, 80.43397, 80.06299, 80.29052, 79.56172, 79.67901, 
    79.60924, 79.35425, 80.17111, 79.751, 80.52818, 80.29965, 80.96806, 
    80.63499, 81.29011, 81.57116, 81.83686, 82.14764, 79.54564, 79.45701, 
    79.61586, 79.83587, 80.04073, 80.31355, 80.34157, 80.39273, 80.52551, 
    80.63722, 80.40881, 80.66526, 79.70602, 80.2077, 79.42342, 79.6588, 
    79.82294, 79.75101, 80.12549, 80.21391, 80.57393, 80.38773, 81.50163, 
    81.00731, 82.38524, 81.99828, 79.42603, 79.54539, 79.96175, 79.76344, 
    80.33185, 80.47217, 80.58647, 80.7326, 80.74847, 80.83517, 80.69312, 
    80.8296, 80.31414, 80.54418, 79.9142, 80.06712, 79.99678, 79.91959, 
    80.15798, 80.41238, 80.41798, 80.49966, 80.72984, 80.33417, 81.56529, 
    80.80294, 79.67569, 79.90606, 79.93922, 79.84985, 80.45808, 80.23728, 
    80.83308, 80.67176, 80.93627, 80.80473, 80.78538, 80.61675, 80.51186, 
    80.24736, 80.03267, 79.86282, 79.90231, 80.08897, 80.42799, 80.74983, 
    80.67922, 80.91615, 80.29053, 80.55231, 80.451, 80.71541, 80.13708, 
    80.62884, 80.01168, 80.06568, 80.2329, 80.56997, 80.64495, 80.72475, 
    80.67554, 80.43665, 80.39764, 80.22887, 80.18224, 80.05393, 79.94775, 
    80.04472, 80.14662, 80.43681, 80.69891, 80.9855, 81.05582, 81.39149, 
    81.11794, 81.56952, 81.18511, 81.85162, 80.65766, 81.17416, 80.24057, 
    80.3408, 80.52212, 80.93956, 80.71416, 80.9779, 80.39612, 80.09533, 
    80.01785, 79.87312, 80.02116, 80.00912, 80.15096, 80.10537, 80.44646, 
    80.26312, 80.78485, 80.97586, 81.5174, 81.85068, 82.19129, 82.34193, 
    82.38783, 82.40701,
  118.1164, 118.6721, 118.5639, 119.0132, 118.7639, 119.0583, 118.2289, 
    118.6942, 118.397, 118.1664, 119.8886, 119.0333, 120.7651, 120.233, 
    121.5715, 120.6823, 121.7514, 121.5458, 122.1655, 121.9877, 122.7827, 
    122.2476, 123.1964, 122.6548, 122.7394, 122.2299, 119.2051, 119.7819, 
    119.171, 119.2531, 119.2163, 118.769, 118.544, 118.074, 118.1593, 
    118.5045, 119.29, 119.023, 119.6969, 119.6817, 120.4296, 120.095, 
    121.3305, 120.98, 121.9951, 121.7392, 121.9831, 121.9091, 121.984, 
    121.6089, 121.7695, 121.4398, 120.1586, 120.5366, 119.3939, 118.7051, 
    118.2493, 117.9266, 117.9722, 118.0591, 118.5066, 118.9284, 119.2506, 
    119.4665, 119.6795, 120.3238, 120.6557, 121.4015, 121.2667, 121.4952, 
    121.7138, 122.0814, 122.0209, 122.1831, 121.4892, 121.95, 121.1899, 
    121.3975, 119.7373, 119.095, 118.8226, 118.5847, 118.0073, 118.4058, 
    118.2486, 118.6229, 118.8612, 118.7433, 119.4724, 119.1886, 120.6754, 
    120.0412, 121.6883, 121.2944, 121.7828, 121.5334, 121.961, 121.5761, 
    122.2435, 122.3891, 122.2896, 122.6724, 121.5548, 121.9831, 118.74, 
    118.7592, 118.8488, 118.4554, 118.4313, 118.0717, 118.3917, 118.5281, 
    118.8751, 119.0806, 119.2763, 119.7072, 120.1899, 120.8475, 121.3199, 
    121.6373, 121.4426, 121.6145, 121.4223, 121.3324, 122.3345, 121.771, 
    122.6172, 122.5703, 122.1869, 122.5756, 118.7728, 118.6622, 118.2787, 
    118.5787, 118.0326, 118.338, 118.5139, 119.1945, 119.3444, 119.4835, 
    119.7586, 120.1124, 120.7194, 121.2451, 121.7265, 121.6912, 121.7036, 
    121.8113, 121.5446, 121.8552, 121.9073, 121.771, 122.564, 122.3371, 
    122.5693, 122.4215, 118.6981, 118.8843, 118.7836, 118.9729, 118.8395, 
    119.4334, 119.6119, 120.4437, 120.1054, 120.641, 120.161, 120.2482, 
    120.6583, 120.1876, 121.216, 120.5197, 121.8155, 121.1175, 121.8594, 
    121.7244, 121.9479, 122.1483, 122.4008, 122.8677, 122.7595, 123.1507, 
    119.1622, 119.4044, 119.3831, 119.637, 119.8249, 120.2331, 120.8695, 
    120.6303, 121.0697, 121.1581, 120.4906, 120.9, 119.5668, 119.7849, 
    119.655, 119.1813, 120.6853, 119.9186, 121.3277, 120.9163, 122.1197, 
    121.5201, 122.6999, 123.2067, 123.6853, 124.2462, 119.5368, 119.3721, 
    119.6672, 120.0763, 120.4507, 120.9414, 120.9917, 121.0838, 121.3228, 
    121.5239, 121.1129, 121.5744, 119.8354, 120.7511, 119.3098, 119.7474, 
    120.0522, 119.9184, 120.603, 120.7621, 121.4101, 121.0748, 123.0815, 
    122.1906, 124.6745, 123.9767, 119.3145, 119.5363, 120.3088, 119.9415, 
    120.9742, 121.2268, 121.4325, 121.6957, 121.7242, 121.8804, 121.6245, 
    121.8703, 120.9424, 121.3564, 120.2216, 120.4982, 120.3716, 120.2316, 
    120.6615, 121.1194, 121.1292, 121.2764, 121.6916, 120.9784, 123.1967, 
    121.8231, 119.7784, 120.2069, 120.2681, 120.102, 121.2015, 120.8042, 
    121.8766, 121.5861, 122.0624, 121.8255, 121.7907, 121.4871, 121.2983, 
    120.8223, 120.4362, 120.1261, 120.1995, 120.5375, 121.1475, 121.7268, 
    121.5997, 122.0261, 120.8999, 121.3712, 121.1888, 121.6647, 120.6239, 
    121.5096, 120.3984, 120.4955, 120.7963, 121.4031, 121.5378, 121.6816, 
    121.5929, 121.163, 121.0927, 120.789, 120.7052, 120.4743, 120.2834, 
    120.4578, 120.6412, 121.1632, 121.6351, 122.1512, 122.2777, 122.8831, 
    122.3901, 123.2044, 122.5117, 123.7126, 121.5612, 122.4915, 120.81, 
    120.9903, 121.3169, 122.0687, 121.6625, 122.1376, 121.09, 120.549, 
    120.4095, 120.1453, 120.4154, 120.3938, 120.6488, 120.5668, 121.1806, 
    120.8506, 121.7898, 122.1339, 123.1096, 123.7105, 124.3245, 124.5963, 
    124.6791, 124.7137,
  186.9665, 187.9677, 187.7727, 188.5827, 188.133, 188.6639, 187.1691, 
    188.0076, 187.472, 187.0564, 190.1565, 188.6189, 191.7155, 190.757, 
    193.172, 191.5661, 193.4971, 193.1255, 194.2455, 193.9241, 195.3624, 
    194.394, 196.1113, 195.1308, 195.2839, 194.3621, 188.9286, 189.9695, 
    188.8671, 189.0152, 188.9487, 188.1423, 187.737, 186.8901, 187.0436, 
    187.6657, 189.0819, 188.6002, 189.8158, 189.7883, 191.1098, 190.5162, 
    192.7365, 192.1034, 193.9375, 193.475, 193.9158, 193.782, 193.9175, 
    193.2395, 193.5298, 192.934, 190.6272, 191.3029, 189.2691, 188.0273, 
    187.2058, 186.6246, 186.7067, 186.8633, 187.6694, 188.4296, 189.0106, 
    189.4, 189.7843, 190.9191, 191.5181, 192.8648, 192.6212, 193.034, 
    193.429, 194.0936, 193.9841, 194.2774, 193.0231, 193.856, 192.4825, 
    192.8574, 189.8891, 188.73, 188.2392, 187.8102, 186.7698, 187.4878, 
    187.2045, 187.879, 188.3085, 188.096, 189.4107, 188.8988, 191.5537, 
    190.4224, 193.3829, 192.6712, 193.5538, 193.103, 193.8759, 193.1802, 
    194.3866, 194.6501, 194.47, 195.1625, 193.1417, 193.9158, 188.0901, 
    188.1247, 188.2862, 187.5771, 187.5338, 186.8859, 187.4623, 187.7082, 
    188.3335, 188.7041, 189.0569, 189.8344, 190.6818, 191.8642, 192.7172, 
    193.2907, 192.9389, 193.2495, 192.9023, 192.7398, 194.5514, 193.5325, 
    195.0628, 194.9779, 194.2844, 194.9874, 188.149, 187.9497, 187.2588, 
    187.7993, 186.8154, 187.3657, 187.6827, 188.9095, 189.1798, 189.4308, 
    189.9272, 190.5465, 191.6329, 192.5822, 193.452, 193.3882, 193.4106, 
    193.6053, 193.1233, 193.6846, 193.7789, 193.5323, 194.9665, 194.5559, 
    194.976, 194.7086, 188.0145, 188.3501, 188.1687, 188.5099, 188.2695, 
    189.3406, 189.6626, 191.1353, 190.5344, 191.4915, 190.6314, 190.7836, 
    191.5229, 190.6778, 192.5298, 191.2727, 193.6129, 192.352, 193.6922, 
    193.4482, 193.8522, 194.2146, 194.6712, 195.5161, 195.3202, 196.0283, 
    188.8513, 189.2882, 189.2497, 189.7076, 190.0451, 190.7572, 191.9039, 
    191.472, 192.2654, 192.425, 191.2199, 191.9591, 189.581, 189.9747, 
    189.7402, 188.8857, 191.5715, 190.2086, 192.7314, 191.9885, 194.1629, 
    193.0791, 195.2124, 196.1301, 196.9967, 198.0135, 189.5269, 189.2297, 
    189.7622, 190.4837, 191.1479, 192.0337, 192.1245, 192.2909, 192.7224, 
    193.0858, 192.3436, 193.177, 190.0637, 191.6902, 189.1175, 189.907, 
    190.4416, 190.2082, 191.4227, 191.7099, 192.8804, 192.2746, 195.9033, 
    194.2913, 198.7904, 197.5249, 189.1259, 189.5259, 190.8918, 190.2485, 
    192.093, 192.5492, 192.9207, 193.3964, 193.4478, 193.7302, 193.2677, 
    193.7119, 192.0356, 192.7833, 190.7371, 191.2335, 191.005, 190.7546, 
    191.5283, 192.3553, 192.3729, 192.6387, 193.3895, 192.1005, 196.1123, 
    193.6271, 189.9628, 190.7115, 190.8184, 190.5284, 192.5034, 191.7859, 
    193.7233, 193.1982, 194.0592, 193.631, 193.568, 193.0193, 192.6782, 
    191.8188, 191.1218, 190.5704, 190.6985, 191.3045, 192.406, 193.4525, 
    193.2229, 193.9936, 191.9588, 192.81, 192.4807, 193.3403, 191.4606, 
    193.0605, 191.0533, 191.2287, 191.7717, 192.8679, 193.111, 193.3709, 
    193.2104, 192.434, 192.307, 191.7585, 191.6073, 191.1905, 190.8459, 
    191.1607, 191.4917, 192.4343, 193.2868, 194.2198, 194.4486, 195.5443, 
    194.652, 196.1262, 194.8725, 197.0467, 193.1535, 194.8356, 191.7964, 
    192.122, 192.7121, 194.0707, 193.3362, 194.1954, 192.302, 191.3255, 
    191.0734, 190.6039, 191.0842, 191.0451, 191.5054, 191.3574, 192.4656, 
    191.8697, 193.5665, 194.1886, 195.954, 197.0426, 198.1554, 198.6483, 
    198.7986, 198.8614,
  314.7132, 316.4507, 316.1122, 317.5189, 316.7377, 317.6599, 315.0646, 
    316.5199, 315.5901, 314.8691, 320.2661, 317.5817, 323.077, 321.3481, 
    325.708, 322.8074, 326.2959, 325.6238, 327.6396, 327.0685, 329.5957, 
    327.8995, 330.9085, 329.1897, 329.458, 327.8437, 318.1201, 319.9308, 
    318.0131, 318.2706, 318.155, 316.7539, 316.0502, 314.5807, 314.8469, 
    315.9264, 318.3865, 317.5493, 319.663, 319.6151, 321.9841, 320.9139, 
    324.9208, 323.7771, 327.0927, 326.2558, 327.0534, 326.8113, 327.0565, 
    325.83, 326.3549, 325.2776, 321.1141, 322.3324, 318.7121, 316.5543, 
    315.1284, 314.1204, 314.2627, 314.5342, 315.9327, 317.2529, 318.2626, 
    318.9398, 319.6083, 321.6405, 322.7208, 325.1526, 324.7123, 325.4585, 
    326.1727, 327.3739, 327.177, 327.6954, 325.4387, 326.9452, 324.4618, 
    325.1393, 319.7908, 317.7749, 316.9222, 316.1772, 314.3722, 315.6177, 
    315.1261, 316.2966, 317.0426, 316.6734, 318.9583, 318.0681, 322.7849, 
    320.745, 326.0893, 324.8026, 326.3984, 325.5831, 326.9813, 325.7227, 
    327.8866, 328.3479, 328.0326, 329.2452, 325.6531, 327.0534, 316.6631, 
    316.7233, 317.0038, 315.7727, 315.6975, 314.5734, 315.5734, 316.0002, 
    317.0858, 317.7298, 318.3431, 319.6955, 321.2125, 323.3453, 324.8859, 
    325.9226, 325.2865, 325.848, 325.2204, 324.9266, 328.175, 326.3599, 
    329.0705, 328.9218, 327.7076, 328.9385, 316.7655, 316.4193, 315.2203, 
    316.1583, 314.4512, 315.4057, 315.9558, 318.0868, 318.5567, 318.9932, 
    319.8569, 320.9686, 322.9279, 324.6419, 326.2142, 326.0988, 326.1394, 
    326.4916, 325.6199, 326.635, 326.8057, 326.3596, 328.9018, 328.1829, 
    328.9186, 328.4503, 316.5318, 317.1147, 316.7996, 317.3925, 316.9747, 
    318.8364, 319.3965, 322.0303, 320.9467, 322.6727, 321.1216, 321.3959, 
    322.7294, 321.2052, 324.5473, 322.278, 326.5053, 324.2263, 326.6487, 
    326.2074, 326.9383, 327.5855, 328.3848, 329.8648, 329.5215, 330.763, 
    317.9856, 318.7453, 318.6782, 319.4749, 320.0653, 321.3484, 323.4169, 
    322.6375, 324.0696, 324.3579, 322.1827, 323.5167, 319.2546, 319.9396, 
    319.5315, 318.0456, 322.8171, 320.3598, 324.9114, 323.5696, 327.4951, 
    325.5401, 329.3327, 330.9417, 332.4626, 334.2497, 319.1605, 318.6435, 
    319.5697, 320.8556, 322.0528, 323.6514, 323.8153, 324.1158, 324.8953, 
    325.5521, 324.211, 325.717, 320.0989, 323.0312, 318.4484, 319.8219, 
    320.7796, 320.359, 322.5485, 323.0667, 325.1807, 324.0862, 330.5439, 
    327.7197, 335.6165, 333.3906, 318.4631, 319.1587, 321.5911, 320.4315, 
    323.7583, 324.5823, 325.2536, 326.1138, 326.2067, 326.7176, 325.8809, 
    326.6844, 323.6548, 325.0053, 321.3121, 322.2073, 321.7951, 321.3437, 
    322.739, 324.2321, 324.2639, 324.7441, 326.1015, 323.7718, 330.9105, 
    326.5312, 319.9189, 321.2661, 321.4588, 320.936, 324.4996, 323.204, 
    326.7051, 325.7552, 327.3129, 326.538, 326.4241, 325.4318, 324.8154, 
    323.2633, 322.0057, 321.0117, 321.2426, 322.3354, 324.3236, 326.2152, 
    325.8, 327.1942, 323.516, 325.0536, 324.4585, 326.0122, 322.6169, 
    325.5066, 321.8823, 322.1985, 323.1783, 325.1582, 325.5975, 326.0676, 
    325.7774, 324.3742, 324.1447, 323.1544, 322.8816, 322.1296, 321.5083, 
    322.0759, 322.6731, 324.3747, 325.9156, 327.5946, 327.995, 329.9144, 
    328.3513, 330.9349, 328.7375, 332.5506, 325.6746, 328.6727, 323.2229, 
    323.8107, 324.8767, 327.3339, 326.0049, 327.552, 324.1357, 322.3732, 
    321.9185, 321.0721, 321.9379, 321.8674, 322.6978, 322.4307, 324.4313, 
    323.3552, 326.4213, 327.5401, 330.6327, 332.5432, 334.4991, 335.3664, 
    335.6309, 335.7415,
  523.2208, 526.4933, 525.8551, 528.509, 527.0347, 528.7754, 523.8821, 
    526.6238, 524.8715, 523.5142, 533.7062, 528.6277, 539.0436, 535.7582, 
    544.0582, 538.5309, 545.1812, 543.8974, 547.7717, 546.6583, 551.6522, 
    548.2866, 554.2629, 550.8459, 551.3788, 548.176, 529.6447, 533.0709, 
    529.4426, 529.9293, 529.7108, 527.0652, 525.7383, 522.9714, 523.4724, 
    525.5051, 530.1483, 528.5663, 532.5636, 532.473, 536.966, 534.9344, 
    542.5559, 540.3761, 546.7047, 545.1046, 546.6295, 546.1664, 546.6355, 
    544.2911, 545.294, 543.2366, 535.3143, 537.6278, 530.7639, 526.6887, 
    524.0021, 522.1059, 522.3735, 522.884, 525.517, 528.0069, 529.9141, 
    531.1946, 532.4599, 536.3134, 538.3661, 542.9982, 542.1583, 543.5818, 
    544.9457, 547.2454, 546.866, 547.8823, 543.544, 546.4225, 541.6807, 
    542.9726, 532.8057, 528.9925, 527.3828, 525.9777, 522.5793, 524.9234, 
    523.9979, 526.2028, 527.6099, 526.9133, 531.2296, 529.5465, 538.4881, 
    534.6141, 544.7864, 542.3306, 545.377, 543.8198, 546.4915, 544.0862, 
    548.261, 549.1755, 548.5504, 550.9561, 543.9533, 546.6296, 526.8939, 
    527.0074, 527.5366, 525.2154, 525.0737, 522.9578, 524.84, 525.644, 
    527.6915, 528.9073, 530.0662, 532.6251, 535.501, 539.5542, 542.4893, 
    544.468, 543.2535, 544.3255, 543.1274, 542.5669, 548.8327, 545.3035, 
    550.6093, 550.314, 547.9066, 550.3472, 527.0872, 526.4342, 524.1751, 
    525.942, 522.728, 524.5242, 525.5605, 529.5819, 530.4702, 531.2958, 
    532.9307, 535.0382, 538.76, 542.0241, 545.0251, 544.8045, 544.8821, 
    545.5553, 543.89, 545.8293, 546.1557, 545.3029, 550.2745, 548.8483, 
    550.3077, 549.3785, 526.6463, 527.746, 527.1515, 528.2703, 527.4819, 
    530.999, 532.0591, 537.0537, 534.9966, 538.2747, 535.3284, 535.8491, 
    538.3826, 535.4871, 541.8438, 537.5245, 545.5815, 541.2319, 545.8555, 
    545.0121, 546.4093, 547.6646, 549.2487, 552.1871, 551.5048, 553.9733, 
    529.3906, 530.8268, 530.6999, 532.2073, 533.3256, 535.7589, 539.6904, 
    538.2078, 540.9333, 541.4827, 537.3432, 539.8803, 531.7903, 533.0875, 
    532.3146, 529.5038, 538.5493, 533.8839, 542.538, 539.9812, 547.4854, 
    543.7376, 551.1298, 554.3289, 557.2599, 560.7106, 531.6123, 530.6342, 
    532.3868, 534.8238, 537.0965, 540.1368, 540.4489, 541.0213, 542.5072, 
    543.7606, 541.2027, 544.0753, 533.3893, 538.9565, 530.2652, 532.8645, 
    534.6797, 533.8823, 538.0386, 539.024, 543.0518, 540.9649, 553.5374, 
    547.9305, 563.3561, 559.0507, 530.2931, 531.6088, 536.2197, 534.0197, 
    540.3404, 541.9104, 543.1907, 544.8332, 545.0107, 545.9872, 544.3882, 
    545.9238, 540.1432, 542.717, 535.6899, 537.39, 536.607, 535.7499, 
    538.4006, 541.2429, 541.3035, 542.2189, 544.8098, 540.3661, 554.267, 
    545.6309, 533.0482, 535.6027, 535.9684, 534.9763, 541.7528, 539.2853, 
    545.9633, 544.1483, 547.126, 545.6438, 545.4262, 543.5308, 542.3549, 
    539.3982, 537.007, 535.12, 535.558, 537.6334, 541.4173, 545.027, 
    544.2338, 546.8989, 539.879, 542.8091, 541.6744, 544.6392, 538.1685, 
    543.6737, 536.7725, 537.3732, 539.2365, 543.0088, 543.8472, 544.7449, 
    544.1907, 541.5137, 541.0765, 539.191, 538.672, 537.2423, 536.0624, 
    537.1404, 538.2755, 541.5146, 544.4547, 547.6825, 548.476, 552.2856, 
    549.1824, 554.3157, 549.9484, 557.4296, 543.9943, 549.8199, 539.3213, 
    540.4402, 542.4717, 547.1663, 544.6252, 547.5982, 541.0593, 537.7054, 
    536.8413, 535.2346, 536.8781, 536.7442, 538.3223, 537.8145, 541.6226, 
    539.5729, 545.4208, 547.5746, 553.7141, 557.4154, 561.1931, 562.8717, 
    563.3839, 563.5983,
  947.124, 953.9968, 952.6537, 958.2476, 955.1371, 958.8105, 948.5101, 
    954.2717, 950.5864, 947.7388, 969.1208, 958.4984, 980.1606, 973.3537, 
    990.6221, 979.096, 992.9768, 990.2852, 998.4262, 996.0811, 1006.634, 
    999.5121, 1012.188, 1004.924, 1006.054, 999.2789, 960.6486, 967.8129, 
    960.221, 961.2509, 960.7884, 955.2015, 952.4081, 946.6017, 947.6512, 
    951.9177, 961.7147, 958.3687, 966.7698, 966.5834, 975.8518, 971.6527, 
    987.4788, 982.932, 996.1787, 992.816, 996.0204, 995.0466, 996.0331, 
    991.1099, 993.2137, 988.9019, 972.4367, 977.2228, 963.019, 954.4083, 
    948.7616, 944.7905, 945.3502, 946.4188, 951.9427, 957.1875, 961.2188, 
    963.9323, 966.5566, 974.5015, 978.754, 988.4033, 986.6482, 989.6245, 
    992.4826, 997.3172, 996.5183, 998.6593, 989.5452, 995.5851, 985.6512, 
    988.3498, 967.2675, 959.2693, 955.8708, 952.9117, 945.7809, 950.6954, 
    948.7528, 953.3853, 956.3499, 954.8815, 964.0067, 960.4409, 979.0072, 
    970.9919, 992.1484, 987.0079, 993.3879, 990.1226, 995.7302, 990.6807, 
    999.4581, 1001.389, 1000.069, 1005.158, 990.4023, 996.0206, 954.8406, 
    955.0798, 956.1953, 951.3088, 951.0112, 946.5731, 950.5201, 952.2098, 
    956.522, 959.0893, 961.5409, 966.8961, 972.8223, 981.2219, 987.3397, 
    991.4807, 988.9374, 991.1822, 988.6735, 987.5017, 1000.665, 993.2335, 
    1004.423, 1003.798, 998.7104, 1003.868, 955.2477, 953.8723, 949.1246, 
    952.8365, 946.092, 949.8573, 952.0343, 960.5157, 962.3965, 964.147, 
    967.5247, 971.8668, 979.5717, 986.368, 992.6492, 992.1864, 992.3494, 
    993.7623, 990.2696, 994.3379, 995.024, 993.2323, 1003.714, 1000.698, 
    1003.784, 1001.818, 954.319, 956.6371, 955.3833, 957.7435, 956.0798, 
    963.5175, 965.7331, 976.0334, 971.7811, 978.5643, 972.466, 973.5416, 
    978.7881, 972.7936, 985.9915, 977.0087, 993.8173, 984.715, 994.393, 
    992.6219, 995.5572, 998.2003, 1001.544, 1007.77, 1006.322, 1011.571, 
    960.1111, 963.1523, 962.8834, 966.0375, 968.337, 973.3551, 981.5052, 
    978.4255, 984.0927, 985.238, 976.6331, 981.9001, 965.1812, 967.8472, 
    966.2579, 960.3507, 979.1342, 969.4866, 987.4415, 982.11, 997.8227, 
    989.9506, 1005.526, 1012.329, 1018.81, 1026.488, 964.8157, 962.7442, 
    966.4064, 971.4244, 976.1221, 982.4338, 983.0836, 984.2761, 987.377, 
    989.9986, 984.6542, 990.6578, 968.4683, 979.9798, 961.9623, 967.3884, 
    971.1271, 969.4833, 978.0745, 980.1201, 988.5153, 984.1585, 1010.642, 
    998.761, 1032.287, 1022.788, 962.0213, 964.8085, 974.3076, 969.7665, 
    982.8576, 986.1307, 988.806, 992.2466, 992.6191, 994.6697, 991.3137, 
    994.5366, 982.4473, 987.8155, 973.2126, 976.73, 975.1088, 973.3365, 
    978.8256, 984.738, 984.8643, 986.7748, 992.1975, 982.9113, 1012.197, 
    993.9211, 967.7662, 973.0325, 973.7881, 971.739, 985.8016, 980.6629, 
    994.6195, 990.8108, 997.0656, 993.9482, 993.4912, 989.5176, 987.0589, 
    980.8976, 975.9368, 972.0356, 972.9401, 977.2344, 985.1017, 992.6532, 
    990.9899, 996.5876, 981.8974, 988.008, 985.6381, 991.8398, 978.3441, 
    989.8168, 975.4514, 976.6952, 980.5614, 988.4255, 990.1802, 992.0616, 
    990.8997, 985.3028, 984.3911, 980.4669, 979.3889, 976.4241, 973.9824, 
    976.213, 978.5659, 985.3048, 991.4528, 998.2382, 999.9117, 1007.98, 
    1001.404, 1012.301, 1003.024, 1019.186, 990.4882, 1002.752, 980.7377, 
    983.0655, 987.3029, 997.1504, 991.8104, 998.0605, 984.3553, 977.3836, 
    975.5938, 972.2721, 975.6699, 975.3928, 978.6631, 977.6099, 985.53, 
    981.2609, 993.4799, 998.0106, 1011.018, 1019.154, 1027.565, 1031.236, 
    1032.348, 1032.813,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.785, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.367, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.287, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.25, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.494, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.374, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.823, 1995.068, 1990.795, 2007.355, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.698, 1840.854, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.441, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.948, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.383, 1967.079, 1965.616, 1966.13, 
    1970.605, 1959.577, 1972.432, 1974.615, 1968.924, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.14, 1901.946, 1923.064, 1904.061, 1907.391, 
    1923.767, 1905.074, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.773, 1874.989, 1884.355, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.876, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.028, 2079.233, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.518, 1872.306, 1888.469, 
    1899.93, 1894.877, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.746, 
    1936.524, 1946.646, 1954.987, 1965.806, 1966.983, 1973.487, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.671, 
    1971.109, 1889.622, 1905.814, 1908.155, 1901.816, 1945.624, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.571, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.083, 1963.301, 1984.896, 1990.287, 2016.643, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.428, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.069, 1944.782, 
    1931.565, 1969.709, 1984.165, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.540418, 4.558938, 4.555333, 4.570301, 4.561993, 4.571801, 4.544168, 
    4.559675, 4.54977, 4.542082, 4.59945, 4.57097, 4.629154, 4.610897, 
    4.65685, 4.62631, 4.663023, 4.655964, 4.677227, 4.671129, 4.6984, 
    4.680043, 4.712574, 4.69401, 4.696912, 4.679439, 4.576689, 4.595898, 
    4.575553, 4.578289, 4.577061, 4.562165, 4.554673, 4.539003, 4.541845, 
    4.553354, 4.579519, 4.570624, 4.59306, 4.592552, 4.617619, 4.606305, 
    4.648574, 4.636533, 4.671383, 4.662602, 4.670971, 4.668432, 4.671004, 
    4.658131, 4.663643, 4.652326, 4.608423, 4.621297, 4.582974, 4.56004, 
    4.544847, 4.534089, 4.535609, 4.538507, 4.553421, 4.567473, 4.578203, 
    4.58539, 4.592479, 4.613988, 4.625396, 4.651012, 4.64638, 4.654227, 
    4.661729, 4.674345, 4.672267, 4.677832, 4.654019, 4.669837, 4.643744, 
    4.650871, 4.594415, 4.573022, 4.563956, 4.556026, 4.536777, 4.550064, 
    4.544824, 4.557297, 4.565237, 4.561308, 4.585587, 4.576138, 4.626073, 
    4.604518, 4.660854, 4.647331, 4.664099, 4.655537, 4.670215, 4.657003, 
    4.679903, 4.6849, 4.681485, 4.694611, 4.656272, 4.670971, 4.561199, 
    4.561839, 4.564823, 4.551716, 4.550915, 4.538926, 4.549592, 4.55414, 
    4.565696, 4.572543, 4.579058, 4.593404, 4.609464, 4.631983, 4.648207, 
    4.659103, 4.652419, 4.65832, 4.651724, 4.648634, 4.683028, 4.663695, 
    4.692721, 4.691112, 4.677964, 4.691293, 4.562289, 4.558604, 4.545827, 
    4.555824, 4.537621, 4.547805, 4.553668, 4.576336, 4.581326, 4.585958, 
    4.595114, 4.606884, 4.627581, 4.64564, 4.662166, 4.660954, 4.66138, 
    4.665078, 4.655923, 4.666582, 4.668373, 4.663692, 4.690896, 4.683113, 
    4.691077, 4.686008, 4.559801, 4.566004, 4.562652, 4.568957, 4.564515, 
    4.584294, 4.590235, 4.618106, 4.606652, 4.624888, 4.608502, 4.611403, 
    4.625487, 4.609386, 4.644644, 4.620723, 4.665222, 4.641265, 4.666726, 
    4.662094, 4.669764, 4.67664, 4.6853, 4.701308, 4.697598, 4.711004, 
    4.575261, 4.583327, 4.582615, 4.591065, 4.597322, 4.6109, 4.632738, 
    4.624517, 4.639615, 4.64265, 4.619715, 4.633789, 4.58873, 4.595991, 
    4.591666, 4.575898, 4.626412, 4.600441, 4.648475, 4.634347, 4.67566, 
    4.655085, 4.695556, 4.712932, 4.729317, 4.748521, 4.587732, 4.582247, 
    4.59207, 4.605688, 4.618344, 4.635209, 4.636936, 4.640101, 4.648305, 
    4.655211, 4.641104, 4.656943, 4.597679, 4.628671, 4.580175, 4.594743, 
    4.604884, 4.600432, 4.623578, 4.629045, 4.651307, 4.639789, 4.708641, 
    4.678095, 4.763172, 4.739296, 4.580332, 4.587712, 4.613466, 4.6012, 
    4.636335, 4.645012, 4.652073, 4.661111, 4.662087, 4.667449, 4.658665, 
    4.667101, 4.635245, 4.649462, 4.610516, 4.619976, 4.615622, 4.61085, 
    4.625587, 4.641326, 4.64166, 4.646715, 4.660983, 4.636478, 4.712597, 
    4.665493, 4.59577, 4.61003, 4.612067, 4.606538, 4.644142, 4.630493, 
    4.667317, 4.657345, 4.673691, 4.665564, 4.664369, 4.653946, 4.647465, 
    4.631119, 4.617846, 4.607339, 4.609781, 4.621328, 4.642289, 4.662176, 
    4.657815, 4.672448, 4.633782, 4.64997, 4.643709, 4.660045, 4.624299, 
    4.654734, 4.616542, 4.619882, 4.630222, 4.651071, 4.655688, 4.660626, 
    4.657578, 4.642822, 4.640406, 4.629971, 4.627093, 4.619154, 4.61259, 
    4.618588, 4.624893, 4.642827, 4.65903, 4.676739, 4.681078, 4.701844, 
    4.684938, 4.712861, 4.689119, 4.730265, 4.656498, 4.688417, 4.630692, 
    4.636888, 4.648109, 4.673912, 4.659968, 4.676277, 4.640311, 4.621728, 
    4.616925, 4.607978, 4.61713, 4.616385, 4.625153, 4.622334, 4.643423, 
    4.632087, 4.66434, 4.676148, 4.709599, 4.730185, 4.751197, 4.760494, 
    4.763326, 4.76451,
  5.632165, 5.655428, 5.650899, 5.669704, 5.659266, 5.671589, 5.636874, 
    5.656354, 5.643912, 5.634254, 5.706334, 5.670544, 5.743674, 5.720722, 
    5.778503, 5.7401, 5.786269, 5.77739, 5.804135, 5.796464, 5.830776, 
    5.807679, 5.848615, 5.825253, 5.828904, 5.806918, 5.677731, 5.70187, 
    5.676303, 5.67974, 5.678197, 5.659482, 5.65007, 5.630388, 5.633957, 
    5.648414, 5.681286, 5.67011, 5.698303, 5.697665, 5.729172, 5.714951, 
    5.768095, 5.752953, 5.796784, 5.785739, 5.796266, 5.793072, 5.796307, 
    5.780114, 5.787048, 5.772813, 5.717612, 5.733796, 5.685629, 5.656814, 
    5.637728, 5.624216, 5.626124, 5.629765, 5.648499, 5.666152, 5.679633, 
    5.688664, 5.697573, 5.724609, 5.73895, 5.771161, 5.765337, 5.775205, 
    5.784641, 5.800511, 5.797896, 5.804896, 5.774943, 5.794838, 5.762021, 
    5.770984, 5.700006, 5.673123, 5.661733, 5.65177, 5.627593, 5.644281, 
    5.637698, 5.653367, 5.663341, 5.658406, 5.688911, 5.677038, 5.739801, 
    5.712705, 5.78354, 5.766531, 5.787621, 5.776852, 5.795314, 5.778697, 
    5.807503, 5.81379, 5.809493, 5.826008, 5.777777, 5.796266, 5.658268, 
    5.659073, 5.662822, 5.646356, 5.64535, 5.630291, 5.643688, 5.649401, 
    5.663919, 5.672521, 5.680707, 5.698735, 5.718921, 5.747232, 5.767633, 
    5.781338, 5.772931, 5.780353, 5.772057, 5.768171, 5.811434, 5.787113, 
    5.82363, 5.821605, 5.805063, 5.821833, 5.659638, 5.655008, 5.638959, 
    5.651516, 5.628653, 5.641443, 5.648808, 5.677288, 5.683557, 5.689378, 
    5.700884, 5.715678, 5.741697, 5.764405, 5.78519, 5.783665, 5.784202, 
    5.788853, 5.777339, 5.790744, 5.792997, 5.787109, 5.821334, 5.811541, 
    5.821562, 5.815184, 5.656513, 5.664305, 5.660094, 5.668016, 5.662435, 
    5.687286, 5.694753, 5.729785, 5.715387, 5.738312, 5.717712, 5.721359, 
    5.739065, 5.718823, 5.763153, 5.733075, 5.789033, 5.758903, 5.790926, 
    5.7851, 5.794747, 5.803398, 5.814292, 5.834435, 5.829766, 5.846639, 
    5.675937, 5.686072, 5.685177, 5.695796, 5.703659, 5.720726, 5.748181, 
    5.737845, 5.756828, 5.760645, 5.731808, 5.749503, 5.692862, 5.701987, 
    5.696551, 5.676736, 5.740228, 5.70758, 5.767971, 5.750205, 5.802164, 
    5.776284, 5.827198, 5.849065, 5.86969, 5.893868, 5.691607, 5.684714, 
    5.697059, 5.714175, 5.730084, 5.751288, 5.753459, 5.75744, 5.767757, 
    5.776443, 5.7587, 5.778621, 5.704108, 5.743067, 5.682111, 5.700418, 
    5.713164, 5.707569, 5.736664, 5.743538, 5.771533, 5.757048, 5.843664, 
    5.805229, 5.912319, 5.882254, 5.682308, 5.691583, 5.723952, 5.708534, 
    5.752705, 5.763616, 5.772495, 5.783864, 5.78509, 5.791834, 5.780787, 
    5.791397, 5.751333, 5.769212, 5.720243, 5.732135, 5.726662, 5.720664, 
    5.739191, 5.75898, 5.7594, 5.765757, 5.783702, 5.752884, 5.848643, 
    5.789376, 5.70171, 5.719633, 5.722193, 5.715244, 5.762521, 5.745358, 
    5.791669, 5.779126, 5.799688, 5.789464, 5.787961, 5.774851, 5.766701, 
    5.746145, 5.729459, 5.716251, 5.71932, 5.733836, 5.760191, 5.785203, 
    5.779718, 5.798123, 5.749494, 5.76985, 5.761977, 5.782522, 5.737571, 
    5.775842, 5.727819, 5.732018, 5.745018, 5.771235, 5.777042, 5.783253, 
    5.77942, 5.760861, 5.757823, 5.744701, 5.741084, 5.731103, 5.722851, 
    5.730391, 5.738317, 5.760868, 5.781246, 5.803521, 5.808981, 5.83511, 
    5.813838, 5.848975, 5.819098, 5.870883, 5.778061, 5.818215, 5.745609, 
    5.753399, 5.767511, 5.799966, 5.782425, 5.802941, 5.757704, 5.734338, 
    5.728301, 5.717054, 5.728558, 5.727622, 5.738644, 5.7351, 5.761617, 
    5.747362, 5.787924, 5.802778, 5.84487, 5.870782, 5.897238, 5.908946, 
    5.912512, 5.914004,
  8.097893, 8.132092, 8.125433, 8.153086, 8.137735, 8.155857, 8.104815, 
    8.133452, 8.115161, 8.100965, 8.206972, 8.154321, 8.26194, 8.228148, 
    8.313241, 8.256677, 8.324682, 8.311601, 8.351015, 8.339708, 8.390292, 
    8.356237, 8.416603, 8.382147, 8.387531, 8.355117, 8.164891, 8.200403, 
    8.162791, 8.167847, 8.165577, 8.138053, 8.124214, 8.095282, 8.100527, 
    8.121778, 8.17012, 8.153682, 8.195155, 8.194217, 8.240587, 8.219654, 
    8.297907, 8.275604, 8.340179, 8.323902, 8.339416, 8.334708, 8.339477, 
    8.315614, 8.325831, 8.304857, 8.223572, 8.247396, 8.176509, 8.134129, 
    8.10607, 8.086209, 8.089015, 8.094366, 8.121903, 8.147861, 8.167689, 
    8.180975, 8.194082, 8.233871, 8.254984, 8.302424, 8.293843, 8.308381, 
    8.322285, 8.345673, 8.341819, 8.352137, 8.307995, 8.337312, 8.28896, 
    8.302162, 8.197661, 8.158113, 8.141362, 8.126713, 8.091172, 8.115704, 
    8.106026, 8.129061, 8.143727, 8.136471, 8.181338, 8.163872, 8.256237, 
    8.216349, 8.320662, 8.295604, 8.326676, 8.310808, 8.338013, 8.313526, 
    8.355978, 8.365247, 8.358912, 8.383261, 8.31217, 8.339417, 8.136268, 
    8.137451, 8.142964, 8.118753, 8.117273, 8.095138, 8.114831, 8.12323, 
    8.144577, 8.157228, 8.169269, 8.195791, 8.225497, 8.267179, 8.297226, 
    8.317417, 8.305031, 8.315966, 8.303743, 8.298018, 8.361773, 8.325928, 
    8.379756, 8.376769, 8.352383, 8.377106, 8.138282, 8.131474, 8.10788, 
    8.12634, 8.092731, 8.111531, 8.122358, 8.164239, 8.173461, 8.182024, 
    8.198954, 8.220724, 8.259028, 8.292471, 8.323093, 8.320847, 8.321637, 
    8.328491, 8.311524, 8.331279, 8.334599, 8.325922, 8.376369, 8.361932, 
    8.376706, 8.367303, 8.133686, 8.145145, 8.138952, 8.150602, 8.142394, 
    8.178947, 8.189933, 8.24149, 8.220296, 8.254045, 8.223718, 8.229086, 
    8.255153, 8.225354, 8.290627, 8.246333, 8.328757, 8.284368, 8.331546, 
    8.322961, 8.337177, 8.349927, 8.365988, 8.39569, 8.388803, 8.413689, 
    8.162251, 8.17716, 8.175845, 8.191467, 8.203036, 8.228156, 8.268576, 
    8.253357, 8.281311, 8.286933, 8.244469, 8.270523, 8.187149, 8.200576, 
    8.192577, 8.163428, 8.256866, 8.208807, 8.297724, 8.271557, 8.348109, 
    8.309971, 8.385015, 8.417268, 8.447699, 8.483386, 8.185304, 8.175163, 
    8.193326, 8.218513, 8.241931, 8.273151, 8.27635, 8.282212, 8.297409, 
    8.310205, 8.284069, 8.313415, 8.203697, 8.261046, 8.171334, 8.198269, 
    8.217025, 8.208791, 8.251618, 8.261739, 8.302971, 8.281634, 8.409301, 
    8.352626, 8.510629, 8.46624, 8.171623, 8.185268, 8.232903, 8.210211, 
    8.275238, 8.291309, 8.30439, 8.321138, 8.322947, 8.332885, 8.316605, 
    8.33224, 8.273218, 8.299552, 8.227445, 8.24495, 8.236893, 8.228063, 
    8.255338, 8.28448, 8.2851, 8.294463, 8.320901, 8.275502, 8.416645, 
    8.329261, 8.200168, 8.226546, 8.230315, 8.220085, 8.289697, 8.26442, 
    8.332642, 8.314158, 8.34446, 8.329391, 8.327177, 8.30786, 8.295853, 
    8.265578, 8.24101, 8.221568, 8.226085, 8.247454, 8.286264, 8.323112, 
    8.31503, 8.342154, 8.270509, 8.300493, 8.288895, 8.319162, 8.252954, 
    8.309319, 8.238597, 8.244778, 8.263919, 8.302532, 8.311089, 8.32024, 
    8.314591, 8.287251, 8.282777, 8.263453, 8.258125, 8.243431, 8.231283, 
    8.242383, 8.254052, 8.287261, 8.317282, 8.35011, 8.358157, 8.396684, 
    8.365316, 8.417134, 8.373072, 8.449458, 8.312589, 8.371771, 8.26479, 
    8.276261, 8.297047, 8.344869, 8.319019, 8.349255, 8.282601, 8.248194, 
    8.239305, 8.22275, 8.239683, 8.238305, 8.254533, 8.249315, 8.288365, 
    8.267371, 8.327123, 8.349014, 8.411079, 8.44931, 8.48836, 8.505648, 
    8.510915, 8.513118,
  12.66457, 12.72004, 12.70923, 12.7541, 12.72919, 12.7586, 12.6758, 
    12.72224, 12.69257, 12.66955, 12.8416, 12.75611, 12.93095, 12.87601, 
    13.01443, 12.92239, 13.03306, 13.01176, 13.07595, 13.05753, 13.13997, 
    13.08446, 13.18288, 13.12669, 13.13547, 13.08263, 12.77326, 12.83093, 
    12.76986, 12.77806, 12.77438, 12.72971, 12.70726, 12.66034, 12.66884, 
    12.70331, 12.78175, 12.75507, 12.82241, 12.82088, 12.89623, 12.86221, 
    12.98947, 12.95318, 13.0583, 13.03179, 13.05705, 13.04939, 13.05715, 
    13.0183, 13.03493, 13.00078, 12.86858, 12.9073, 12.79212, 12.72334, 
    12.67783, 12.64563, 12.65018, 12.65885, 12.70351, 12.74562, 12.77781, 
    12.79938, 12.82066, 12.88531, 12.91964, 12.99682, 12.98286, 13.00652, 
    13.02916, 13.06725, 13.06097, 13.07778, 13.00589, 13.05363, 12.97491, 
    12.9964, 12.82648, 12.76226, 12.73508, 12.71131, 12.65368, 12.69345, 
    12.67776, 12.71512, 12.73892, 12.72714, 12.79997, 12.77161, 12.92168, 
    12.85684, 13.02651, 12.98572, 13.03631, 13.01047, 13.05477, 13.01489, 
    13.08404, 13.09914, 13.08882, 13.12851, 13.01269, 13.05706, 12.72681, 
    12.72873, 12.73768, 12.6984, 12.696, 12.66011, 12.69204, 12.70566, 
    12.74029, 12.76083, 12.78037, 12.82344, 12.87171, 12.93947, 12.98836, 
    13.02123, 13.00107, 13.01887, 12.99897, 12.98965, 13.09348, 13.03509, 
    13.12279, 13.11792, 13.07818, 13.11847, 12.73008, 12.71903, 12.68077, 
    12.71071, 12.6562, 12.68669, 12.70425, 12.77221, 12.78718, 12.80108, 
    12.82858, 12.86395, 12.92622, 12.98062, 13.03047, 13.02681, 13.0281, 
    13.03926, 13.01164, 13.0438, 13.04921, 13.03508, 13.11727, 13.09374, 
    13.11782, 13.10249, 12.72262, 12.74122, 12.73117, 12.75007, 12.73675, 
    12.79608, 12.81392, 12.8977, 12.86325, 12.91811, 12.86881, 12.87754, 
    12.91992, 12.87147, 12.97762, 12.90557, 13.0397, 12.96744, 13.04424, 
    13.03026, 13.05341, 13.07418, 13.10035, 13.14877, 13.13754, 13.17813, 
    12.76898, 12.79318, 12.79105, 12.81642, 12.83521, 12.87603, 12.94175, 
    12.917, 12.96247, 12.97161, 12.90254, 12.94491, 12.8094, 12.83121, 
    12.81822, 12.77089, 12.9227, 12.84458, 12.98917, 12.9466, 13.07122, 
    13.00911, 13.13137, 13.18397, 13.23363, 13.29191, 12.80641, 12.78994, 
    12.81944, 12.86035, 12.89842, 12.94919, 12.95439, 12.96393, 12.98866, 
    13.00949, 12.96695, 13.01471, 12.83628, 12.9295, 12.78372, 12.82746, 
    12.85794, 12.84456, 12.91417, 12.93063, 12.99771, 12.96299, 13.17097, 
    13.07858, 13.33643, 13.2639, 12.78419, 12.80635, 12.88374, 12.84686, 
    12.95258, 12.97873, 13.00002, 13.02729, 13.03023, 13.04642, 13.01991, 
    13.04537, 12.9493, 12.99215, 12.87487, 12.90333, 12.89023, 12.87588, 
    12.92022, 12.96762, 12.96863, 12.98387, 13.0269, 12.95301, 13.18295, 
    13.04052, 12.83055, 12.87341, 12.87953, 12.86291, 12.97611, 12.93499, 
    13.04602, 13.01593, 13.06527, 13.04073, 13.03712, 13.00567, 12.98613, 
    12.93687, 12.89692, 12.86532, 12.87266, 12.9074, 12.97052, 13.0305, 
    13.01734, 13.06151, 12.94489, 12.99368, 12.9748, 13.02407, 12.91634, 
    13.00805, 12.893, 12.90305, 12.93417, 12.997, 13.01093, 13.02583, 
    13.01663, 12.97213, 12.96485, 12.93341, 12.92475, 12.90086, 12.88111, 
    12.89915, 12.91813, 12.97215, 13.02101, 13.07448, 13.08759, 13.15039, 
    13.09926, 13.18375, 13.1119, 13.2365, 13.01337, 13.10977, 12.93559, 
    12.95425, 12.98807, 13.06594, 13.02384, 13.07308, 12.96456, 12.9086, 
    12.89415, 12.86724, 12.89476, 12.89252, 12.91891, 12.91042, 12.97394, 
    12.93979, 13.03703, 13.07269, 13.17387, 13.23626, 13.30004, 13.32829, 
    13.33689, 13.34049,
  20.59555, 20.6916, 20.67289, 20.75065, 20.70747, 20.75845, 20.61498, 
    20.69543, 20.64403, 20.60417, 20.90253, 20.75413, 21.05791, 20.96234, 
    21.20336, 21.04301, 21.23585, 21.1987, 21.31072, 21.27856, 21.4226, 
    21.32558, 21.49769, 21.39938, 21.41473, 21.32239, 20.78389, 20.88399, 
    20.77798, 20.79221, 20.78582, 20.70836, 20.66946, 20.58822, 20.60294, 
    20.66262, 20.79862, 20.75233, 20.86919, 20.86654, 20.9975, 20.93834, 
    21.15984, 21.09661, 21.2799, 21.23364, 21.27773, 21.26435, 21.2779, 
    21.2101, 21.23912, 21.17956, 20.9494, 21.01675, 20.81661, 20.69733, 
    20.6185, 20.56278, 20.57064, 20.58566, 20.66297, 20.73595, 20.79177, 
    20.8292, 20.86616, 20.9785, 21.03822, 21.17266, 21.14831, 21.18956, 
    21.22904, 21.29552, 21.28456, 21.31391, 21.18847, 21.27175, 21.13446, 
    21.17191, 20.87625, 20.7648, 20.71767, 20.67648, 20.5767, 20.64555, 
    20.61838, 20.68308, 20.72432, 20.70391, 20.83022, 20.78102, 21.04177, 
    20.929, 21.22443, 21.15331, 21.24152, 21.19645, 21.27374, 21.20417, 
    21.32484, 21.35123, 21.3332, 21.40255, 21.20032, 21.27773, 20.70334, 
    20.70667, 20.72218, 20.65412, 20.64996, 20.58782, 20.6431, 20.66669, 
    20.72671, 20.76231, 20.79622, 20.87098, 20.95484, 21.07274, 21.15791, 
    21.21522, 21.18005, 21.21109, 21.1764, 21.16016, 21.34134, 21.23939, 
    21.39256, 21.38405, 21.31461, 21.38501, 20.70901, 20.68987, 20.62358, 
    20.67544, 20.58107, 20.63383, 20.66425, 20.78205, 20.80803, 20.83216, 
    20.8799, 20.94136, 21.04967, 21.14442, 21.23134, 21.22495, 21.2272, 
    21.24667, 21.19848, 21.2546, 21.26403, 21.23937, 21.38291, 21.34179, 
    21.38387, 21.35708, 20.69608, 20.72831, 20.71089, 20.74366, 20.72057, 
    20.82349, 20.85446, 21.00005, 20.94015, 21.03556, 20.94982, 20.96498, 
    21.0387, 20.95444, 21.13919, 21.01375, 21.24743, 21.12144, 21.25536, 
    21.23096, 21.27136, 21.30763, 21.35334, 21.43799, 21.41836, 21.48936, 
    20.77645, 20.81845, 20.81474, 20.85878, 20.89142, 20.96235, 21.0767, 
    21.03362, 21.11278, 21.12872, 21.00847, 21.08222, 20.84661, 20.88448, 
    20.86192, 20.77977, 21.04355, 20.90771, 21.15932, 21.08515, 21.30245, 
    21.19407, 21.40755, 21.49958, 21.58658, 21.68879, 20.84141, 20.81282, 
    20.86403, 20.93511, 21.0013, 21.08966, 21.09872, 21.11534, 21.15843, 
    21.19474, 21.1206, 21.20385, 20.89328, 21.05538, 20.80204, 20.87797, 
    20.93091, 20.90766, 21.0287, 21.05734, 21.17421, 21.1137, 21.47684, 
    21.3153, 21.76696, 21.63965, 20.80285, 20.8413, 20.97577, 20.91167, 
    21.09557, 21.14113, 21.17823, 21.22579, 21.23092, 21.25916, 21.21291, 
    21.25733, 21.08985, 21.16451, 20.96035, 21.00983, 20.98705, 20.96209, 
    21.03922, 21.12177, 21.12352, 21.15007, 21.22511, 21.09632, 21.4978, 
    21.24886, 20.88333, 20.95781, 20.96846, 20.93955, 21.13655, 21.06493, 
    21.25847, 21.20597, 21.29207, 21.24924, 21.24294, 21.18808, 21.15401, 
    21.06821, 20.99869, 20.94374, 20.9565, 21.01692, 21.12682, 21.23139, 
    21.20844, 21.28551, 21.08218, 21.16718, 21.13428, 21.22017, 21.03248, 
    21.19222, 20.99187, 21.00935, 21.06351, 21.17296, 21.19725, 21.22323, 
    21.20719, 21.12962, 21.11694, 21.06219, 21.04711, 21.00554, 20.9712, 
    21.00257, 21.03559, 21.12965, 21.21483, 21.30815, 21.33105, 21.44083, 
    21.35143, 21.4992, 21.37352, 21.59161, 21.20151, 21.36981, 21.06598, 
    21.09847, 21.1574, 21.29324, 21.21977, 21.30571, 21.11644, 21.01901, 
    20.99387, 20.94708, 20.99494, 20.99104, 21.03695, 21.02218, 21.13278, 
    21.07329, 21.24279, 21.30503, 21.48191, 21.59119, 21.70305, 21.75266, 
    21.76778, 21.77411,
  34.63898, 34.81974, 34.78448, 34.93107, 34.84964, 34.94579, 34.67551, 
    34.82695, 34.73016, 34.65519, 35.21814, 34.93763, 35.51294, 35.33147, 
    35.78992, 35.48462, 35.85194, 35.78104, 35.99503, 35.93353, 36.20937, 
    36.02347, 36.35357, 36.16483, 36.19426, 36.01736, 34.9938, 35.18304, 
    34.98264, 35.00952, 34.99745, 34.85132, 34.77803, 34.62521, 34.65288, 
    34.76515, 35.02161, 34.93423, 35.15502, 35.15001, 35.39818, 35.28597, 
    35.70694, 35.58654, 35.93609, 35.84771, 35.93194, 35.90636, 35.93227, 
    35.80278, 35.85817, 35.74453, 35.30695, 35.43474, 35.05562, 34.83053, 
    34.68213, 34.5774, 34.59218, 34.62038, 34.76581, 34.90334, 35.00868, 
    35.07941, 35.1493, 35.36214, 35.47552, 35.73137, 35.68498, 35.7636, 
    35.83894, 35.96596, 35.945, 36.00114, 35.76151, 35.92051, 35.6586, 
    35.72995, 35.1684, 34.95778, 34.86886, 34.79126, 34.60355, 34.73302, 
    34.6819, 34.80369, 34.88141, 34.84294, 35.08134, 34.98838, 35.48226, 
    35.26828, 35.83014, 35.69449, 35.86276, 35.77674, 35.92432, 35.79146, 
    36.02205, 36.07257, 36.03804, 36.17092, 35.78412, 35.93194, 34.84186, 
    34.84813, 34.87736, 34.74915, 34.74133, 34.62445, 34.72841, 34.77283, 
    34.88592, 34.95307, 35.01708, 35.15842, 35.31726, 35.54114, 35.70326, 
    35.81255, 35.74547, 35.80468, 35.7385, 35.70755, 36.05363, 35.8587, 
    36.15176, 36.13545, 36.00248, 36.13729, 34.85254, 34.81647, 34.69169, 
    34.78928, 34.61176, 34.71098, 34.76822, 34.99033, 35.03939, 35.085, 
    35.1753, 35.2917, 35.49728, 35.67757, 35.84332, 35.83113, 35.83543, 
    35.8726, 35.78062, 35.88774, 35.90577, 35.85867, 36.13327, 36.05449, 
    36.1351, 36.08378, 34.82819, 34.88893, 34.85609, 34.91788, 34.87434, 
    35.0686, 35.12716, 35.40303, 35.28941, 35.47047, 35.30774, 35.33649, 
    35.47643, 35.3165, 35.6676, 35.42903, 35.87405, 35.6338, 35.88919, 
    35.8426, 35.91978, 35.98911, 36.07661, 36.23891, 36.20123, 36.33757, 
    34.97977, 35.05909, 35.05208, 35.13534, 35.19711, 35.33151, 35.54867, 
    35.46677, 35.61732, 35.64766, 35.41902, 35.55915, 35.11231, 35.18396, 
    35.14127, 34.98602, 35.48564, 35.22794, 35.70595, 35.56473, 35.97921, 
    35.77221, 36.18051, 36.35721, 36.52464, 36.72184, 35.10248, 35.04845, 
    35.14526, 35.27986, 35.4054, 35.57332, 35.59056, 35.62218, 35.70425, 
    35.77348, 35.63219, 35.79086, 35.20063, 35.50813, 35.02807, 35.17164, 
    35.2719, 35.22786, 35.45743, 35.51186, 35.73433, 35.61906, 36.31349, 
    36.0038, 36.87302, 36.62698, 35.02961, 35.10229, 35.35696, 35.23545, 
    35.58456, 35.67129, 35.742, 35.83272, 35.84253, 35.89646, 35.80815, 
    35.89296, 35.57368, 35.71584, 35.3277, 35.4216, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63776, 35.68833, 35.83143, 35.58599, 36.35379, 
    35.87679, 35.18179, 35.32288, 35.34308, 35.28828, 35.66258, 35.52629, 
    35.89514, 35.79489, 35.95936, 35.87749, 35.86547, 35.76078, 35.69584, 
    35.53252, 35.40045, 35.29622, 35.32042, 35.43505, 35.64405, 35.84343, 
    35.79961, 35.94682, 35.55908, 35.72092, 35.65825, 35.82201, 35.4646, 
    35.76868, 35.3875, 35.42068, 35.52359, 35.73195, 35.77826, 35.82785, 
    35.79724, 35.64937, 35.62523, 35.52108, 35.49241, 35.41345, 35.34827, 
    35.40782, 35.47051, 35.64943, 35.81181, 35.9901, 36.03392, 36.24435, 
    36.07294, 36.35648, 36.11526, 36.53433, 35.78639, 36.10815, 35.52828, 
    35.59008, 35.70229, 35.96159, 35.82123, 35.98545, 35.62428, 35.43902, 
    35.3913, 35.30255, 35.39333, 35.38593, 35.4731, 35.44505, 35.65539, 
    35.54218, 35.86518, 35.98414, 36.32325, 36.53352, 36.7494, 36.84534, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34589, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59598, 62.19373, 
    63.21417, 62.53307, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73952, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13967, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47564, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13955, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25315, 61.48349, 
    61.63854, 61.79207, 62.26156, 62.51286, 63.08306, 62.97935, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.6428, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73633, 63.85044, 63.77242, 64.07315, 63.20119, 63.5332, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36182, 61.5019, 61.81213, 62.16233, 62.65869, 63.02021, 
    63.26492, 63.11462, 63.24727, 63.09903, 63.02979, 63.80764, 63.36849, 
    64.02972, 63.99276, 63.69214, 63.99692, 61.14231, 61.06372, 60.79243, 
    61.00454, 60.61915, 60.8343, 60.95869, 61.44333, 61.55079, 61.65081, 
    61.84928, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31625, 
    63.39974, 63.19335, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18986, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40972, 63.40299, 62.86511, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59398, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49344, 62.82833, 62.89602, 62.38752, 62.69877, 61.71079, 61.86834, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.09491, 64.49689, 64.87986, 65.33361, 61.68919, 61.57066, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86152, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75535, 62.94876, 63.10686, 63.31018, 63.33219, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29745, 62.19272, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86355, 62.17475, 62.2194, 62.09832, 62.92932, 62.62566, 
    63.4504, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00362, 
    62.63952, 62.34638, 62.11584, 62.16929, 62.42306, 62.88795, 63.3342, 
    63.23591, 63.5667, 62.69861, 63.0597, 62.91965, 63.28613, 62.48863, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26327, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65374, 62.84386, 62.43187, 
    62.3261, 62.12982, 62.33061, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38306, 63.65079, 64.41946, 64.90024, 65.39728, 65.61928, 
    65.68716, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7406, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02022763, -0.01989731, -0.01996107, -0.01969795, -0.01984346, 
    -0.01967183, -0.0201602, -0.0198843, -0.02005997, -0.02019767, 
    -0.01919786, -0.01968631, -0.01870443, -0.01900581, -0.01825852, 
    -0.01875097, -0.01816094, -0.01827257, -0.0179389, -0.01803381, 
    -0.01761414, -0.01789527, -0.01740083, -0.01768086, -0.01763672, 
    -0.01790462, -0.01958698, -0.01925795, -0.01960665, -0.01955932, 
    -0.01958055, -0.01984043, -0.01997278, -0.02025314, -0.02020193, 
    -0.01999618, -0.01953807, -0.01969233, -0.01930613, -0.01931476, 
    -0.01889415, -0.01908256, -0.01839036, -0.01858431, -0.01802984, 
    -0.01816757, -0.01803628, -0.01807598, -0.01803576, -0.01823822, 
    -0.01815118, -0.01833045, -0.01904711, -0.01883339, -0.01947855, 
    -0.01987785, -0.02014801, -0.02034208, -0.02031452, -0.02026209, 
    -0.01999498, -0.01974732, -0.01956079, -0.01943707, -0.019316, 
    -0.01895435, -0.01876597, -0.01835139, -0.0184255, -0.01830017, 
    -0.01818134, -0.01798366, -0.01801604, -0.01792951, -0.01830349, 
    -0.018054, -0.01846785, -0.01835365, -0.0192831, -0.01965059, 
    -0.01980896, -0.0199488, -0.02029336, -0.02005473, -0.02014843, 
    -0.01992629, -0.0197865, -0.01985551, -0.0194337, -0.01959653, 
    -0.01875486, -0.01911253, -0.01819515, -0.01841027, -0.018144, 
    -0.01827935, -0.01804809, -0.01825608, -0.01789743, -0.01782034, 
    -0.01787298, -0.01767172, -0.01826769, -0.01803627, -0.01985744, 
    -0.01984617, -0.01979374, -0.02002531, -0.02003957, -0.02025454, 
    -0.02006315, -0.01998223, -0.01977843, -0.01965892, -0.01954603, 
    -0.01930028, -0.01902972, -0.01865826, -0.01839624, -0.01822283, 
    -0.01832896, -0.01823522, -0.01834004, -0.01838939, -0.01784918, 
    -0.01815036, -0.01770052, -0.01772509, -0.01792746, -0.01772232, 
    -0.01983825, -0.0199032, -0.02013044, -0.01995237, -0.0202781, 
    -0.02009506, -0.01999061, -0.01959308, -0.01950692, -0.01942735, 
    -0.01927124, -0.01907286, -0.01873015, -0.01843739, -0.01817445, 
    -0.01819358, -0.01818684, -0.01812861, -0.01827322, -0.01810499, 
    -0.01807691, -0.01815041, -0.01772839, -0.01784786, -0.01772562, 
    -0.0178033, -0.01988207, -0.01977305, -0.01983188, -0.0197214, 
    -0.01979915, -0.01945589, -0.01935422, -0.01888608, -0.01907674, 
    -0.0187743, -0.01904579, -0.01899737, -0.01876447, -0.01903102, 
    -0.01845338, -0.01884285, -0.01812635, -0.01850779, -0.01810273, 
    -0.01817558, -0.01805514, -0.017948, -0.0178142, -0.01757011, 
    -0.01762631, -0.01742429, -0.01961172, -0.01947249, -0.01948472, 
    -0.01934007, -0.01923384, -0.01900575, -0.01864597, -0.0187804, 
    -0.01853443, -0.01848546, -0.01885948, -0.01862886, -0.01937992, 
    -0.01925637, -0.01932984, -0.01960068, -0.0187493, -0.01918113, 
    -0.01839194, -0.01861978, -0.01796323, -0.01828654, -0.01765733, 
    -0.01739548, -0.01715298, -0.01687412, -0.01939697, -0.01949106, 
    -0.01932296, -0.0190929, -0.01888214, -0.01860579, -0.01857778, 
    -0.01852657, -0.01839466, -0.01828453, -0.01851039, -0.01825704, 
    -0.0192278, -0.01871232, -0.01952674, -0.01927753, -0.01910639, 
    -0.01918128, -0.01879583, -0.0187062, -0.01834668, -0.01853161, 
    -0.0174597, -0.01792542, -0.01666516, -0.01700736, -0.01952405, 
    -0.01939731, -0.01896303, -0.01916834, -0.01858751, -0.01844746, 
    -0.01833447, -0.01819109, -0.0181757, -0.0180914, -0.01822976, 
    -0.01809685, -0.01860521, -0.01837615, -0.01901216, -0.01885519, 
    -0.01892723, -0.01900658, -0.01876283, -0.0185068, -0.01850141, 
    -0.01842014, -0.01819312, -0.0185852, -0.01740049, -0.01812208, 
    -0.01926011, -0.01902026, -0.01898631, -0.01907865, -0.01846145, 
    -0.01868255, -0.01809345, -0.01825067, -0.01799385, -0.01812097, 
    -0.01813975, -0.01830464, -0.01840811, -0.01867235, -0.01889037, 
    -0.01906523, -0.01902442, -0.01883288, -0.01849127, -0.01817429, 
    -0.01824322, -0.01801323, -0.01862898, -0.01836804, -0.01846841, 
    -0.01820794, -0.01878398, -0.01829212, -0.01891197, -0.01885673, 
    -0.01868697, -0.01835046, -0.01827695, -0.01819875, -0.01824697, 
    -0.0184827, -0.01852164, -0.01869109, -0.01873815, -0.01886874, 
    -0.01897759, -0.01887811, -0.01877423, -0.01848261, -0.01822398, 
    -0.01794647, -0.01787927, -0.01756201, -0.01781976, -0.01739655, 
    -0.01775558, -0.01713909, -0.0182641, -0.01776633, -0.0186793, 
    -0.01857856, -0.01839779, -0.01799041, -0.01820915, -0.01795363, 
    -0.01852318, -0.01882629, -0.01890563, -0.01905454, -0.01890224, 
    -0.01891458, -0.01876996, -0.01881631, -0.01847301, -0.01865657, 
    -0.01814022, -0.01795564, -0.01744533, -0.01714026, -0.01683571, 
    -0.01670311, -0.01666298, -0.01664624,
  -0.05397912, -0.05293612, -0.05313723, -0.0523081, -0.05276638, 
    -0.05222589, -0.05376598, -0.05289511, -0.05344935, -0.05388441, 
    -0.05073763, -0.05227144, -0.04919505, -0.05013639, -0.04780718, 
    -0.04934024, -0.04750423, -0.0478508, -0.04681598, -0.04711, -0.04581207, 
    -0.04668094, -0.04515439, -0.04601805, -0.04588176, -0.04670988, 
    -0.05195899, -0.05092593, -0.05202086, -0.05187203, -0.05193878, 
    -0.05275683, -0.05317415, -0.0540598, -0.05389789, -0.053248, 
    -0.05180525, -0.05229039, -0.05107701, -0.05110408, -0.04978732, 
    -0.05037652, -0.04821691, -0.04882059, -0.04709769, -0.04752481, 
    -0.04711764, -0.04724073, -0.04711604, -0.04774414, -0.04747394, 
    -0.04803064, -0.0502656, -0.04959753, -0.05161822, -0.05287476, 
    -0.05372744, -0.05434122, -0.054254, -0.05408812, -0.05324422, 
    -0.05246353, -0.05187666, -0.05148795, -0.05110798, -0.04997546, 
    -0.04938704, -0.04809575, -0.04832621, -0.04793655, -0.04756754, 
    -0.04695462, -0.04705494, -0.04678693, -0.04794686, -0.04717259, 
    -0.04845798, -0.04810276, -0.05100481, -0.05215906, -0.05265765, 
    -0.0530985, -0.05418704, -0.0534328, -0.05372879, -0.05302753, 
    -0.05258689, -0.05280435, -0.05147737, -0.05198902, -0.0493524, 
    -0.05047034, -0.04761042, -0.04827882, -0.04745169, -0.04787188, 
    -0.04715426, -0.04779959, -0.04668763, -0.04644912, -0.04661196, 
    -0.04598982, -0.04783563, -0.04711761, -0.05281045, -0.05277491, 
    -0.05260972, -0.05333992, -0.05338496, -0.05406423, -0.05345941, 
    -0.05320399, -0.0525615, -0.05218526, -0.05183026, -0.05105866, 
    -0.05021119, -0.04905107, -0.04823519, -0.04769632, -0.04802601, 
    -0.04773481, -0.04806045, -0.0482139, -0.04653831, -0.04747141, 
    -0.04607876, -0.04615469, -0.04678057, -0.04614612, -0.05274997, 
    -0.05295471, -0.05367194, -0.05310978, -0.05413876, -0.05356017, 
    -0.05323042, -0.05197819, -0.05170734, -0.05145741, -0.05096762, 
    -0.05034618, -0.04927529, -0.04836318, -0.04754617, -0.04760554, 
    -0.04758463, -0.04740393, -0.04785282, -0.04733067, -0.04724359, 
    -0.04747156, -0.04616486, -0.04653425, -0.0461563, -0.04639642, 
    -0.05288808, -0.05254453, -0.05272987, -0.0523819, -0.05262677, 
    -0.05154703, -0.05122788, -0.0497621, -0.05035832, -0.04941304, 
    -0.05026146, -0.05010999, -0.04938237, -0.05021525, -0.04841293, 
    -0.04962708, -0.04739692, -0.04858228, -0.04732366, -0.04754968, 
    -0.04717612, -0.04684416, -0.04643012, -0.04567619, -0.04584963, 
    -0.04522666, -0.05203679, -0.05159917, -0.05163762, -0.0511835, 
    -0.05085035, -0.0501362, -0.04901276, -0.04943209, -0.04866523, 
    -0.04851278, -0.04967902, -0.04895943, -0.05130852, -0.050921, 
    -0.05115141, -0.05200208, -0.04933503, -0.0506852, -0.04822181, 
    -0.04893113, -0.04689133, -0.04789419, -0.04594538, -0.04513793, 
    -0.04439203, -0.04353658, -0.05136206, -0.05165754, -0.0511298, 
    -0.05040889, -0.0497498, -0.04888754, -0.04880025, -0.04864076, 
    -0.04823028, -0.04788796, -0.04859038, -0.04780256, -0.05083142, 
    -0.04921967, -0.05176964, -0.05098733, -0.05045112, -0.05068567, 
    -0.04948027, -0.04920058, -0.04808111, -0.04865645, -0.04533575, 
    -0.04677427, -0.04289719, -0.04394502, -0.05176118, -0.05136311, 
    -0.0500026, -0.05064513, -0.04883058, -0.04839453, -0.04804315, 
    -0.0475978, -0.04755003, -0.04728852, -0.04771785, -0.04730542, 
    -0.04888572, -0.04817273, -0.05015624, -0.04966561, -0.04989071, 
    -0.05013881, -0.04937725, -0.04857922, -0.04856243, -0.04830951, 
    -0.04760409, -0.04882337, -0.04515333, -0.04738366, -0.05093271, 
    -0.05018158, -0.05007539, -0.05036429, -0.04843806, -0.04912683, 
    -0.04729489, -0.04778278, -0.04698617, -0.04738024, -0.0474385, 
    -0.04795045, -0.04827211, -0.049095, -0.04977551, -0.05032229, 
    -0.0501946, -0.04959593, -0.04853088, -0.04754566, -0.04775963, 
    -0.04704622, -0.04895981, -0.0481475, -0.04845972, -0.0476501, 
    -0.04944326, -0.04791154, -0.04984299, -0.04967042, -0.04914061, 
    -0.04809285, -0.04786441, -0.04762158, -0.04777129, -0.04850418, 
    -0.04862543, -0.04915344, -0.04930023, -0.04970795, -0.05004814, 
    -0.0497372, -0.04941282, -0.04850391, -0.04769991, -0.04683944, 
    -0.04663142, -0.0456512, -0.04644732, -0.04514121, -0.0462489, 
    -0.04434937, -0.04782449, -0.04628212, -0.04911667, -0.04880268, 
    -0.04824001, -0.04697552, -0.04765387, -0.04686161, -0.04863019, 
    -0.04957535, -0.04982318, -0.05028885, -0.04981259, -0.04985115, 
    -0.04939951, -0.04954418, -0.04847404, -0.0490458, -0.04743994, 
    -0.04686784, -0.04529148, -0.04435296, -0.04341895, -0.04301323, 
    -0.04289054, -0.04283937,
  -0.07871142, -0.07706042, -0.07737859, -0.07606745, -0.07679196, 
    -0.07593752, -0.07837384, -0.07699556, -0.07787254, -0.0785614, 
    -0.0735881, -0.07600951, -0.07115819, -0.07264037, -0.06897667, 
    -0.07138666, -0.06850109, -0.06904516, -0.06742147, -0.06788254, 
    -0.06584877, -0.06720977, -0.06481982, -0.06617125, -0.06595786, 
    -0.06725515, -0.07551583, -0.0738851, -0.07561357, -0.07537846, 
    -0.0754839, -0.07677686, -0.07743701, -0.07883923, -0.07858275, 
    -0.07755386, -0.07527298, -0.07603946, -0.07412342, -0.07416613, 
    -0.0720905, -0.07301879, -0.06962023, -0.07056914, -0.06786323, 
    -0.0685334, -0.06789453, -0.06808762, -0.06789202, -0.06887769, 
    -0.06845356, -0.06932762, -0.07284396, -0.07179166, -0.07497764, 
    -0.07696337, -0.07831282, -0.07928513, -0.07914691, -0.07888409, 
    -0.07754788, -0.07631312, -0.07538578, -0.07477198, -0.07417228, 
    -0.07238684, -0.07146032, -0.06942989, -0.06979197, -0.06917983, 
    -0.06860045, -0.06763885, -0.06779617, -0.06737594, -0.06919602, 
    -0.06798072, -0.06999906, -0.06944089, -0.07400952, -0.07583191, 
    -0.07662003, -0.0773173, -0.0790408, -0.07784636, -0.07831495, 
    -0.07720502, -0.07650815, -0.07685202, -0.07475527, -0.07556327, 
    -0.07140579, -0.07316667, -0.06866777, -0.0697175, -0.06841863, 
    -0.06907827, -0.06795198, -0.06896476, -0.06722026, -0.06684647, 
    -0.06710166, -0.06612704, -0.06902135, -0.06789448, -0.07686165, 
    -0.07680544, -0.07654424, -0.07769934, -0.07777062, -0.07884624, 
    -0.07788846, -0.07748422, -0.076468, -0.07587332, -0.07531249, 
    -0.07409448, -0.07275823, -0.07093167, -0.06964895, -0.06880262, 
    -0.06932034, -0.06886305, -0.06937443, -0.0696155, -0.06698624, 
    -0.06844959, -0.06626631, -0.06638522, -0.06736595, -0.06637181, 
    -0.07676601, -0.07708983, -0.07822493, -0.07733515, -0.07896432, 
    -0.07804798, -0.07752604, -0.07554615, -0.07511837, -0.07472376, 
    -0.07395084, -0.07297097, -0.07128445, -0.06985006, -0.06856692, 
    -0.06866011, -0.06862728, -0.06834368, -0.06904834, -0.06822872, 
    -0.06809211, -0.06844983, -0.06640116, -0.06697986, -0.06638775, 
    -0.06676389, -0.07698443, -0.07644118, -0.07673422, -0.07618409, 
    -0.07657119, -0.07486524, -0.0743615, -0.07205078, -0.0729901, 
    -0.07150124, -0.07283745, -0.07259877, -0.07145297, -0.07276462, 
    -0.06992826, -0.07183819, -0.06833269, -0.07019445, -0.06821773, 
    -0.06857242, -0.06798626, -0.06746566, -0.0668167, -0.0656361, 
    -0.06590756, -0.06493283, -0.07563873, -0.07494757, -0.07500827, 
    -0.07429145, -0.07376588, -0.07264006, -0.07087139, -0.07153121, 
    -0.07032485, -0.07008519, -0.07191996, -0.0707875, -0.07448875, 
    -0.0738773, -0.07424081, -0.0755839, -0.07137845, -0.07350542, 
    -0.06962793, -0.07074299, -0.06753962, -0.06911331, -0.06605747, 
    -0.06479409, -0.06362849, -0.06229345, -0.07457325, -0.07503971, 
    -0.07420672, -0.07306981, -0.07203142, -0.07067443, -0.07053716, 
    -0.07028639, -0.06964124, -0.06910352, -0.07020719, -0.06896942, 
    -0.07373603, -0.07119692, -0.07521676, -0.07398194, -0.07313637, 
    -0.07350617, -0.07160706, -0.07116689, -0.06940689, -0.07031105, 
    -0.06510346, -0.06735608, -0.06129685, -0.06293062, -0.07520338, 
    -0.0745749, -0.07242958, -0.07344224, -0.07058486, -0.06989934, 
    -0.06934726, -0.06864797, -0.06857298, -0.06816259, -0.06883642, 
    -0.06818912, -0.07067157, -0.06955081, -0.07267164, -0.07189884, 
    -0.07225333, -0.07264418, -0.0714449, -0.07018964, -0.07016324, 
    -0.06976573, -0.06865785, -0.07057352, -0.06481819, -0.06831189, 
    -0.07389577, -0.07271158, -0.07254426, -0.07299951, -0.06996775, 
    -0.07105084, -0.06817259, -0.06893835, -0.06768834, -0.06830651, 
    -0.06839794, -0.06920166, -0.06970696, -0.07100077, -0.07207191, 
    -0.07293332, -0.07273208, -0.07178913, -0.07011364, -0.06856612, 
    -0.06890202, -0.06778251, -0.07078809, -0.06951118, -0.07000179, 
    -0.06873005, -0.0715488, -0.06914055, -0.07217818, -0.07190642, 
    -0.07107252, -0.06942532, -0.06906655, -0.06868529, -0.06892032, 
    -0.07007167, -0.07026228, -0.07109271, -0.07132369, -0.07196551, 
    -0.07250132, -0.07201157, -0.07150089, -0.07007126, -0.06880826, 
    -0.06745825, -0.06713215, -0.06559701, -0.06684365, -0.06479923, 
    -0.06653281, -0.06356186, -0.06900387, -0.06658484, -0.07103487, 
    -0.07054098, -0.06965654, -0.06767163, -0.06873597, -0.06749302, 
    -0.07026977, -0.07175674, -0.07214698, -0.07288061, -0.0721303, 
    -0.07219103, -0.07147994, -0.07170767, -0.0700243, -0.07092337, 
    -0.06840019, -0.06750278, -0.06503422, -0.06356747, -0.06211002, 
    -0.06147763, -0.0612865, -0.06120677,
  -0.08618353, -0.08427349, -0.08464147, -0.0831254, -0.08396304, 
    -0.08297521, -0.08579286, -0.08419848, -0.08521285, -0.08600991, 
    -0.08026101, -0.08305842, -0.07745696, -0.07916695, -0.07494241, 
    -0.07772047, -0.07439461, -0.07502131, -0.07315151, -0.07368231, 
    -0.07134196, -0.07290784, -0.07015888, -0.07171289, -0.07146743, 
    -0.07296006, -0.08248782, -0.08060396, -0.08260078, -0.08232907, 
    -0.08245092, -0.08394558, -0.08470904, -0.08633143, -0.08603461, 
    -0.0848442, -0.0822072, -0.08309303, -0.08087917, -0.0809285, 
    -0.07853242, -0.07960373, -0.07568392, -0.07677772, -0.07366008, 
    -0.07443181, -0.07369611, -0.07391843, -0.07369322, -0.07482839, 
    -0.07433986, -0.07534675, -0.07940193, -0.07818764, -0.08186593, 
    -0.08416127, -0.08572226, -0.08684757, -0.08668757, -0.08638337, 
    -0.08483729, -0.08340939, -0.08233754, -0.08162832, -0.0809356, 
    -0.07887437, -0.07780542, -0.07546459, -0.07588185, -0.07517647, 
    -0.07450904, -0.07340175, -0.07358287, -0.07309909, -0.07519511, 
    -0.07379535, -0.07612053, -0.07547726, -0.08074765, -0.08285314, 
    -0.08376424, -0.08457059, -0.08656475, -0.08518256, -0.08572473, 
    -0.08444072, -0.08363488, -0.08403248, -0.08160901, -0.08254264, 
    -0.07774253, -0.07977444, -0.07458658, -0.07579603, -0.07429963, 
    -0.07505945, -0.07376225, -0.07492869, -0.07291992, -0.07248974, 
    -0.07278342, -0.07166202, -0.07499388, -0.07369605, -0.08404361, 
    -0.08397863, -0.0836766, -0.08501249, -0.08509494, -0.08633956, 
    -0.08523127, -0.08476365, -0.08358846, -0.08290099, -0.08225284, 
    -0.08084575, -0.07930298, -0.07719573, -0.07571702, -0.07474191, 
    -0.07533836, -0.07481152, -0.07540068, -0.07567847, -0.07265058, 
    -0.07433528, -0.07182223, -0.07195903, -0.0730876, -0.0719436, 
    -0.08393303, -0.08430749, -0.08562056, -0.08459122, -0.08647621, 
    -0.08541582, -0.08481202, -0.08252287, -0.08202853, -0.08157261, 
    -0.08067986, -0.07954854, -0.07760257, -0.0759488, -0.07447042, 
    -0.07457776, -0.07453994, -0.07421332, -0.07502497, -0.07408092, 
    -0.07392361, -0.07433555, -0.07197737, -0.07264324, -0.07196194, 
    -0.07239471, -0.08418561, -0.08355745, -0.08389628, -0.08326023, 
    -0.08370776, -0.08173608, -0.08115415, -0.0784866, -0.07957061, 
    -0.07785263, -0.07939442, -0.07911894, -0.07779696, -0.07931035, 
    -0.07603893, -0.07824133, -0.07420065, -0.07634576, -0.07406826, 
    -0.07447675, -0.07380173, -0.07320237, -0.07245547, -0.07109738, 
    -0.07140958, -0.07028879, -0.08262986, -0.08183119, -0.08190131, 
    -0.08107325, -0.08046627, -0.0791666, -0.07712621, -0.0778872, 
    -0.07649607, -0.0762198, -0.07833565, -0.07702949, -0.08130115, 
    -0.08059495, -0.08101475, -0.08256649, -0.077711, -0.08016553, 
    -0.0756928, -0.07697816, -0.07328751, -0.07509983, -0.071582, 
    -0.07012931, -0.06878995, -0.06725701, -0.08139874, -0.08193765, 
    -0.08097537, -0.07966264, -0.07846425, -0.07689911, -0.07674084, 
    -0.07645173, -0.07570814, -0.07508855, -0.07636043, -0.07493406, 
    -0.08043181, -0.07750162, -0.08214222, -0.08071578, -0.07973947, 
    -0.08016639, -0.07797468, -0.07746699, -0.07543809, -0.07648016, 
    -0.07048495, -0.07307625, -0.06611346, -0.06798849, -0.08212676, 
    -0.08140065, -0.07892369, -0.08009258, -0.07679582, -0.07600559, 
    -0.07536938, -0.07456376, -0.0744774, -0.07400478, -0.07478084, 
    -0.07403532, -0.07689581, -0.07560393, -0.07920305, -0.07831129, 
    -0.0787203, -0.07917134, -0.07778763, -0.07634021, -0.07630978, 
    -0.07585161, -0.07457516, -0.07678276, -0.07015703, -0.07417672, 
    -0.08061627, -0.07924914, -0.07905603, -0.07958147, -0.07608444, 
    -0.07733315, -0.07401628, -0.07489827, -0.07345872, -0.0741705, 
    -0.0742758, -0.07520162, -0.07578388, -0.07727541, -0.07851098, 
    -0.07950507, -0.0792728, -0.07818472, -0.07625261, -0.0744695, 
    -0.07485642, -0.07356714, -0.07703017, -0.07555826, -0.07612368, 
    -0.07465832, -0.07790748, -0.07513123, -0.07863358, -0.07832003, 
    -0.07735815, -0.07545933, -0.07504595, -0.07460675, -0.07487749, 
    -0.07620423, -0.07642394, -0.07738143, -0.07764784, -0.07838821, 
    -0.07900649, -0.07844134, -0.07785222, -0.07620375, -0.0747484, 
    -0.07319385, -0.07281851, -0.07105243, -0.0724865, -0.07013524, 
    -0.07212884, -0.06871344, -0.07497375, -0.07218871, -0.07731473, 
    -0.07674524, -0.07572577, -0.07343949, -0.07466514, -0.07323387, 
    -0.07643258, -0.07814736, -0.07859759, -0.07944423, -0.07857834, 
    -0.07864842, -0.07782806, -0.07809074, -0.07614963, -0.07718615, 
    -0.07427839, -0.07324512, -0.07040534, -0.06871986, -0.06704647, 
    -0.06632084, -0.06610157, -0.06601012,
  -0.06731972, -0.06577227, -0.0660704, -0.06484208, -0.06552074, 
    -0.06472041, -0.06700322, -0.0657115, -0.06653332, -0.06717907, 
    -0.06252129, -0.06478783, -0.06024929, -0.06163482, -0.05821183, 
    -0.0604628, -0.05776796, -0.05827576, -0.05676073, -0.05719081, 
    -0.05529455, -0.0565633, -0.05433598, -0.05559508, -0.05539621, 
    -0.05660561, -0.06432551, -0.06279916, -0.06441703, -0.0641969, 
    -0.06429562, -0.0655066, -0.06612515, -0.06743955, -0.06719907, 
    -0.06623465, -0.06409815, -0.06481586, -0.06302214, -0.06306212, 
    -0.06112069, -0.06198872, -0.05881265, -0.05969892, -0.0571728, 
    -0.0577981, -0.057202, -0.05738214, -0.05719965, -0.05811943, -0.0577236, 
    -0.05853945, -0.06182522, -0.06084133, -0.06382164, -0.06568135, 
    -0.06694602, -0.06785769, -0.06772807, -0.06748162, -0.06622905, 
    -0.06507218, -0.06420375, -0.06362913, -0.06306786, -0.06139776, 
    -0.06053163, -0.05863493, -0.05897302, -0.05840148, -0.05786068, 
    -0.05696348, -0.05711024, -0.05671826, -0.05841658, -0.05728241, 
    -0.05916642, -0.0586452, -0.06291559, -0.0646215, -0.06535968, 
    -0.06601297, -0.06762857, -0.06650878, -0.06694803, -0.06590775, 
    -0.06525487, -0.06557701, -0.06361348, -0.06436993, -0.06048067, 
    -0.06212704, -0.05792351, -0.05890349, -0.057691, -0.05830666, 
    -0.05725559, -0.05820071, -0.05657308, -0.05622452, -0.05646248, 
    -0.05555387, -0.05825353, -0.05720195, -0.06558603, -0.06553338, 
    -0.06528867, -0.06637099, -0.0664378, -0.06744613, -0.06654824, 
    -0.06616938, -0.06521726, -0.06466027, -0.06413513, -0.06299506, 
    -0.06174504, -0.06003761, -0.05883947, -0.05804937, -0.05853265, 
    -0.05810577, -0.05858315, -0.05880823, -0.05635485, -0.05771989, 
    -0.05568368, -0.05579452, -0.05670895, -0.05578202, -0.06549644, 
    -0.06579982, -0.06686363, -0.06602969, -0.06755684, -0.06669775, 
    -0.06620858, -0.06435391, -0.06395338, -0.06358399, -0.06286065, 
    -0.061944, -0.06036727, -0.05902728, -0.05782939, -0.05791636, 
    -0.05788572, -0.05762107, -0.05827872, -0.0575138, -0.05738633, 
    -0.05772011, -0.05580937, -0.0563489, -0.05579688, -0.05614753, 
    -0.06570107, -0.06519213, -0.06546665, -0.06495133, -0.06531392, 
    -0.06371644, -0.06324494, -0.06108356, -0.06196189, -0.06056988, 
    -0.06181912, -0.06159592, -0.06052478, -0.06175101, -0.05910031, 
    -0.06088483, -0.05761081, -0.05934892, -0.05750354, -0.05783452, 
    -0.05728757, -0.05680194, -0.05619676, -0.05509637, -0.05534932, 
    -0.05444123, -0.06444059, -0.0637935, -0.06385031, -0.06317939, 
    -0.06268759, -0.06163453, -0.05998129, -0.06059789, -0.05947071, 
    -0.05924686, -0.06096125, -0.05990292, -0.06336404, -0.06279185, 
    -0.063132, -0.06438926, -0.06045512, -0.06244392, -0.05881985, 
    -0.05986133, -0.05687093, -0.05833939, -0.05548903, -0.05431202, 
    -0.05322686, -0.05198491, -0.06344312, -0.06387975, -0.06310008, 
    -0.06203645, -0.06106545, -0.05979728, -0.05966903, -0.05943478, 
    -0.05883227, -0.05833024, -0.05936081, -0.05820506, -0.06265968, 
    -0.06028548, -0.0640455, -0.06288976, -0.0620987, -0.06244462, 
    -0.06066878, -0.06025741, -0.05861346, -0.05945782, -0.05460016, 
    -0.05669975, -0.05105847, -0.05257753, -0.06403297, -0.06344466, 
    -0.06143772, -0.06238481, -0.05971359, -0.05907329, -0.05855779, 
    -0.05790503, -0.05783505, -0.05745209, -0.05808092, -0.05747684, 
    -0.05979461, -0.05874784, -0.06166407, -0.06094152, -0.06127292, 
    -0.06163838, -0.06051721, -0.05934442, -0.05931976, -0.05894853, 
    -0.05791427, -0.059703, -0.05433448, -0.05759142, -0.06280912, 
    -0.06170142, -0.06154495, -0.06197068, -0.05913718, -0.06014897, 
    -0.05746142, -0.05817606, -0.05700965, -0.05758637, -0.05767169, 
    -0.05842186, -0.05889364, -0.06010218, -0.06110331, -0.06190878, 
    -0.06172059, -0.06083897, -0.05927344, -0.05782864, -0.05814215, 
    -0.05709749, -0.05990347, -0.05871083, -0.05916898, -0.05798164, 
    -0.06061433, -0.05836483, -0.06120265, -0.0609486, -0.06016922, 
    -0.05863068, -0.05829572, -0.05793986, -0.05815922, -0.05923424, 
    -0.05941226, -0.06018809, -0.06040395, -0.06100384, -0.0615048, 
    -0.06104689, -0.06056955, -0.05923385, -0.05805463, -0.05679503, 
    -0.05649091, -0.05505996, -0.05622191, -0.05431682, -0.05593212, 
    -0.05316487, -0.05823722, -0.05598062, -0.06013404, -0.05967261, 
    -0.05884656, -0.05699407, -0.05798716, -0.05682747, -0.05941926, 
    -0.06080869, -0.06117349, -0.06185949, -0.0611579, -0.06121467, 
    -0.06054997, -0.06076281, -0.05919, -0.06002986, -0.0576738, -0.05683658, 
    -0.05453566, -0.05317008, -0.05181434, -0.05122647, -0.05104884, 
    -0.05097476,
  -0.06391447, -0.06222167, -0.06254755, -0.06120564, -0.06194681, 
    -0.06107282, -0.06356799, -0.06215525, -0.0630538, -0.06376047, 
    -0.05867587, -0.06114641, -0.05620678, -0.0577116, -0.0539992, 
    -0.05643849, -0.05351913, -0.05406837, -0.05243094, -0.05289539, 
    -0.05084988, -0.05221782, -0.04981819, -0.05117367, -0.05095939, 
    -0.05226349, -0.0606419, -0.05897837, -0.06074176, -0.06050161, 
    -0.06060929, -0.06193136, -0.06260741, -0.06404568, -0.06378238, 
    -0.06272715, -0.0603939, -0.06117702, -0.05922118, -0.05926472, 
    -0.05715287, -0.05809643, -0.05464952, -0.05560982, -0.05287593, 
    -0.05355172, -0.05290747, -0.0531021, -0.05290494, -0.05389925, 
    -0.05347117, -0.05435374, -0.05791861, -0.05684945, -0.06009239, 
    -0.0621223, -0.06350539, -0.0645037, -0.0643617, -0.06409176, 
    -0.06272102, -0.06145686, -0.06050908, -0.05988252, -0.05927098, 
    -0.05745393, -0.05651321, -0.0544571, -0.0548232, -0.05420442, 
    -0.05361939, -0.05264986, -0.05280836, -0.05238508, -0.05422076, 
    -0.05299434, -0.0550327, -0.05446822, -0.05910514, -0.06096487, 
    -0.06177086, -0.06248477, -0.0642527, -0.06302696, -0.06350757, 
    -0.06236975, -0.06165637, -0.06200828, -0.05986547, -0.06069036, 
    -0.05645789, -0.05824688, -0.05368733, -0.05474789, -0.05343593, 
    -0.05410181, -0.05296537, -0.05398717, -0.05222838, -0.0518523, 
    -0.05210903, -0.05112926, -0.05404432, -0.05290742, -0.06201814, 
    -0.06196061, -0.06169329, -0.06287625, -0.06294932, -0.06405289, 
    -0.06307013, -0.06265578, -0.0616153, -0.06100719, -0.06043423, 
    -0.05919169, -0.05783143, -0.05597714, -0.05467856, -0.05382345, 
    -0.05434638, -0.05388446, -0.05440104, -0.05464473, -0.05199289, 
    -0.05346716, -0.05126915, -0.05138862, -0.05237504, -0.05137515, 
    -0.06192025, -0.06225177, -0.06341521, -0.06250305, -0.06417414, 
    -0.0632337, -0.06269864, -0.06067289, -0.06023603, -0.05983333, 
    -0.05904532, -0.05804779, -0.05633481, -0.05488196, -0.05358555, 
    -0.0536796, -0.05364647, -0.05336033, -0.05407158, -0.05324438, 
    -0.05310663, -0.0534674, -0.05140464, -0.05198648, -0.05139116, 
    -0.05176925, -0.06214385, -0.06158786, -0.06188772, -0.06132491, 
    -0.06172087, -0.0599777, -0.05946387, -0.05711254, -0.05806725, 
    -0.05655472, -0.05791198, -0.05766932, -0.05650576, -0.05783793, 
    -0.05496107, -0.05689669, -0.05334923, -0.05523045, -0.0532333, 
    -0.0535911, -0.05299992, -0.05247543, -0.05182235, -0.05063646, 
    -0.05090889, -0.04993139, -0.06076746, -0.0600617, -0.06012364, 
    -0.05939246, -0.0588569, -0.05771129, -0.05591604, -0.05658513, 
    -0.05536243, -0.05511985, -0.05697969, -0.05583104, -0.05959363, 
    -0.05897041, -0.05934083, -0.06071145, -0.05643016, -0.05859167, 
    -0.05465731, -0.05578594, -0.05254991, -0.05413722, -0.0510594, 
    -0.04979242, -0.04862646, -0.04729465, -0.0596798, -0.06015574, 
    -0.05930608, -0.05814834, -0.05709287, -0.05571648, -0.05557742, 
    -0.05532349, -0.05467076, -0.05412732, -0.05524332, -0.05399187, 
    -0.05882651, -0.05624605, -0.06033648, -0.05907702, -0.05821606, 
    -0.05859243, -0.05666208, -0.05621559, -0.05443385, -0.05534846, 
    -0.05010237, -0.05236511, -0.04630303, -0.0479298, -0.06032282, 
    -0.05968149, -0.05749736, -0.05852734, -0.05562573, -0.05493181, 
    -0.05437359, -0.05366734, -0.05359167, -0.0531777, -0.05385758, 
    -0.05320444, -0.05571358, -0.05457934, -0.0577434, -0.05695825, 
    -0.05731827, -0.05771548, -0.05649755, -0.05522557, -0.05519884, 
    -0.05479667, -0.05367734, -0.05561425, -0.04981658, -0.05332828, 
    -0.05898922, -0.05778401, -0.05761391, -0.05807681, -0.05500102, 
    -0.05609794, -0.05318778, -0.0539605, -0.05269971, -0.05332283, 
    -0.05341506, -0.05422647, -0.05473723, -0.05604718, -0.05713399, 
    -0.05800948, -0.05780485, -0.05684688, -0.05514865, -0.05358474, 
    -0.05392382, -0.05279458, -0.05583163, -0.05453927, -0.05503546, 
    -0.05375019, -0.05660297, -0.05416476, -0.05724192, -0.05696595, 
    -0.05611991, -0.05445249, -0.05408997, -0.05370501, -0.05394229, 
    -0.05510618, -0.05529909, -0.05614038, -0.05637461, -0.05702594, 
    -0.05757027, -0.05707271, -0.05655436, -0.05510575, -0.05382914, 
    -0.05246797, -0.05213971, -0.05059725, -0.05184948, -0.04979759, 
    -0.05153696, -0.04855993, -0.05402667, -0.05158925, -0.05608174, 
    -0.0555813, -0.05468624, -0.05268289, -0.05375617, -0.05250299, 
    -0.05530667, -0.056814, -0.05721024, -0.05795588, -0.05719329, 
    -0.05725498, -0.0565331, -0.05676418, -0.05505824, -0.05596872, 
    -0.05341733, -0.05251282, -0.05003298, -0.04856551, -0.04711195, 
    -0.04648273, -0.04629274, -0.04621351,
  -0.04035198, -0.03907359, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009016, -0.03902347, -0.03970177, -0.0402356, 
    -0.03640241, -0.03826259, -0.03454811, -0.03567765, -0.03289467, 
    -0.03472191, -0.0325357, -0.03294641, -0.03172283, -0.03206963, 
    -0.03054395, -0.03156378, -0.02977613, -0.03078516, -0.03062552, 
    -0.03159786, -0.03788236, -0.03662992, -0.0379576, -0.03777665, 
    -0.03785779, -0.03885455, -0.03936473, -0.04045115, -0.04025215, 
    -0.03945512, -0.03769551, -0.03828567, -0.0368126, -0.03684536, 
    -0.03525804, -0.0359668, -0.03338129, -0.03410057, -0.03205509, 
    -0.03256006, -0.03207865, -0.03222404, -0.03207676, -0.03281991, 
    -0.03249985, -0.03315991, -0.03583318, -0.03503027, -0.03746841, 
    -0.03899861, -0.04004287, -0.0407974, -0.04069003, -0.04048597, 
    -0.0394505, -0.03849666, -0.03778228, -0.03731038, -0.03685007, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351131, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306041, 
    -0.03214354, -0.03366819, -0.03324559, -0.03672529, -0.03812575, 
    -0.03873348, -0.03927216, -0.04060763, -0.0396815, -0.04004452, 
    -0.03918534, -0.03864712, -0.03891259, -0.03729754, -0.03791887, 
    -0.03473647, -0.03607988, -0.03266144, -0.03345493, -0.0324735, 
    -0.03297142, -0.0321219, -0.03288567, -0.03157166, -0.03129108, 
    -0.0314826, -0.03075207, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887662, -0.03867497, -0.0395677, -0.03962287, -0.04045659, 
    -0.0397141, -0.03940124, -0.03861614, -0.03815764, -0.03772589, 
    -0.03679041, -0.03576767, -0.03437591, -0.03340303, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319531, -0.03337771, -0.03139596, 
    -0.03249685, -0.03085631, -0.03094536, -0.03168111, -0.03093531, 
    -0.03884617, -0.03909631, -0.03997475, -0.03928595, -0.04054824, 
    -0.03983764, -0.0394336, -0.03790571, -0.0375766, -0.03727334, 
    -0.03668029, -0.03593025, -0.03464414, -0.03355532, -0.03258535, 
    -0.03265566, -0.03263089, -0.032417, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249703, -0.03095729, -0.03139117, -0.03094725, 
    -0.03122914, -0.03901487, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869577, -0.03738204, -0.03699523, -0.03522776, -0.03594487, 
    -0.03480911, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240871, -0.03381631, -0.03232207, 
    -0.0325895, -0.03214771, -0.03175604, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797697, -0.0374453, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567741, -0.03433011, -0.03483192, 
    -0.03391519, -0.03373347, -0.03512803, -0.03426639, -0.0370929, 
    -0.03662394, -0.03690264, -0.03793476, -0.03471566, -0.03633909, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299791, -0.03070002, 
    -0.02975696, -0.02889069, -0.02790317, -0.03715776, -0.03751612, 
    -0.03687648, -0.03600582, -0.03521299, -0.03418051, -0.03407629, 
    -0.03388602, -0.03339719, -0.03299051, -0.03382596, -0.03288919, 
    -0.0365157, -0.03457757, -0.03765226, -0.03670414, -0.03605671, 
    -0.03633966, -0.03488967, -0.03455472, -0.03321987, -0.03390472, 
    -0.02998751, -0.0316737, -0.02716934, -0.02837385, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629072, -0.03411249, -0.03359264, 
    -0.03317476, -0.0326465, -0.03258992, -0.03228053, -0.03278875, 
    -0.03230051, -0.03417834, -0.03332876, -0.03570153, -0.03511194, 
    -0.03538223, -0.03568055, -0.03476622, -0.03381266, -0.03379264, 
    -0.03349145, -0.03265397, -0.03410389, -0.02977493, -0.03239306, 
    -0.03663808, -0.03573204, -0.03560426, -0.03595205, -0.03364447, 
    -0.03446649, -0.03228806, -0.03286572, -0.03192349, -0.03238898, 
    -0.03245791, -0.03306468, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199434, -0.03426683, -0.03329876, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301851, -0.0353249, -0.03511771, 
    -0.03448297, -0.03323382, -0.03296256, -0.03267466, -0.0328521, 
    -0.03372323, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480884, -0.03372291, -0.03276749, 
    -0.03175048, -0.03150549, -0.03035583, -0.03128898, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.03407919, -0.03340878, -0.03191093, -0.03271292, -0.03177662, 
    -0.03387342, -0.03500367, -0.03530111, -0.03586118, -0.03528839, 
    -0.0353347, -0.03479289, -0.03496628, -0.03368732, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993588, -0.02884545, -0.02776788, 
    -0.02730223, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.0189572, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277074, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459348, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927695, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  297.7961, 299.0511, 298.8069, 299.8214, 299.2584, 299.9231, 298.0503, 
    299.101, 298.4299, 297.909, 301.7971, 299.8668, 303.7903, 302.5721, 
    305.638, 303.6005, 306.0502, 305.5793, 306.9988, 306.5916, 308.4124, 
    307.1869, 309.36, 308.1195, 308.3132, 307.1465, 300.2548, 301.5568, 
    300.1777, 300.3631, 300.2799, 299.2699, 298.7618, 297.7005, 297.8929, 
    298.6727, 300.4465, 299.8435, 301.3653, 301.3309, 303.0214, 302.2617, 
    305.0861, 304.2829, 306.6086, 306.0224, 306.581, 306.4116, 306.5832, 
    305.7238, 306.0918, 305.3365, 302.4048, 303.2665, 300.6809, 299.1254, 
    298.0963, 297.3675, 297.4704, 297.6667, 298.6772, 299.6299, 300.3575, 
    300.845, 301.3259, 302.7787, 303.5397, 305.2486, 304.9398, 305.4632, 
    305.9641, 306.8063, 306.6676, 307.0391, 305.4495, 306.5052, 304.764, 
    305.2394, 301.4561, 300.0061, 299.3909, 298.8538, 297.5496, 298.4497, 
    298.0946, 298.9401, 299.4783, 299.212, 300.8583, 300.2174, 303.5848, 
    302.1407, 305.9057, 305.0032, 306.1223, 305.5509, 306.5305, 305.6487, 
    307.1775, 307.511, 307.283, 308.1599, 305.5999, 306.581, 299.2046, 
    299.248, 299.4503, 298.5616, 298.5074, 297.6952, 298.4178, 298.726, 
    299.5095, 299.9736, 300.4154, 301.3885, 302.4751, 303.9791, 305.0616, 
    305.7889, 305.3428, 305.7366, 305.2964, 305.0903, 307.386, 306.0952, 
    308.0336, 307.9261, 307.0479, 307.9382, 299.2784, 299.0287, 298.1627, 
    298.8403, 297.6068, 298.2967, 298.6938, 300.2307, 300.5693, 300.8834, 
    301.5046, 302.3008, 303.6856, 304.8903, 305.9933, 305.9124, 305.9409, 
    306.1876, 305.5766, 306.288, 306.4075, 306.0951, 307.9117, 307.3919, 
    307.9238, 307.5853, 299.1099, 299.5303, 299.3031, 299.7305, 299.4293, 
    300.7703, 301.1732, 303.0536, 302.2851, 303.506, 302.4103, 302.6064, 
    303.5454, 302.4701, 304.8236, 303.2279, 306.1972, 304.5979, 306.2976, 
    305.9885, 306.5005, 306.9595, 307.5379, 308.6071, 308.3593, 309.2552, 
    300.158, 300.7048, 300.6568, 301.2299, 301.6541, 302.5725, 304.0296, 
    303.4815, 304.4885, 304.6909, 303.1614, 304.0996, 301.0714, 301.5637, 
    301.2706, 300.201, 303.6075, 301.8648, 305.0795, 304.1371, 306.894, 
    305.5204, 308.2229, 309.3835, 310.4796, 311.7636, 301.0038, 300.6318, 
    301.2982, 302.2197, 303.0698, 304.1945, 304.3098, 304.5209, 305.0683, 
    305.5291, 304.5875, 305.6447, 301.6775, 303.7583, 300.4911, 301.479, 
    302.1654, 301.8644, 303.4189, 303.7835, 305.2684, 304.5002, 309.0966, 
    307.0564, 312.7444, 311.1466, 300.5019, 301.0025, 302.7445, 301.9164, 
    304.2697, 304.8485, 305.3197, 305.9228, 305.988, 306.3458, 305.7596, 
    306.3227, 304.1969, 305.1454, 302.5466, 303.1786, 302.8885, 302.5692, 
    303.5529, 304.6023, 304.6249, 304.962, 305.913, 304.2793, 309.3604, 
    306.2142, 301.5492, 302.5133, 302.6514, 302.2776, 304.7904, 303.88, 
    306.3371, 305.6715, 306.7627, 306.2201, 306.1403, 305.4447, 305.0122, 
    303.9216, 303.0366, 302.3318, 302.4969, 303.2687, 304.6666, 305.9938, 
    305.7027, 306.6797, 304.0994, 305.1792, 304.7614, 305.8517, 303.4669, 
    305.4961, 302.9499, 303.1725, 303.8619, 305.2523, 305.561, 305.8904, 
    305.6871, 304.7022, 304.5412, 303.8452, 303.6531, 303.124, 302.6864, 
    303.0862, 303.5064, 304.7027, 305.7838, 306.966, 307.256, 308.6423, 
    307.5131, 309.3779, 307.7915, 310.5419, 305.6143, 307.7453, 303.8934, 
    304.3066, 305.0549, 306.7769, 305.8465, 306.935, 304.5349, 303.2952, 
    302.9753, 302.3749, 302.989, 302.9393, 303.524, 303.336, 304.7425, 
    303.9864, 306.1382, 306.9265, 309.1612, 310.5372, 311.9432, 312.5654, 
    312.7549, 312.8342 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.356944e-08, 6.384899e-08, 6.379465e-08, 6.402013e-08, 6.389505e-08, 
    6.404269e-08, 6.362611e-08, 6.38601e-08, 6.371073e-08, 6.359461e-08, 
    6.445772e-08, 6.403019e-08, 6.490177e-08, 6.462912e-08, 6.531402e-08, 
    6.485934e-08, 6.540569e-08, 6.53009e-08, 6.56163e-08, 6.552594e-08, 
    6.592938e-08, 6.565801e-08, 6.61385e-08, 6.586457e-08, 6.590742e-08, 
    6.564905e-08, 6.411622e-08, 6.44045e-08, 6.409914e-08, 6.414025e-08, 
    6.41218e-08, 6.389764e-08, 6.378468e-08, 6.354806e-08, 6.359102e-08, 
    6.376479e-08, 6.415873e-08, 6.4025e-08, 6.436202e-08, 6.435441e-08, 
    6.47296e-08, 6.456043e-08, 6.519103e-08, 6.50118e-08, 6.552971e-08, 
    6.539947e-08, 6.552359e-08, 6.548596e-08, 6.552408e-08, 6.533306e-08, 
    6.541491e-08, 6.524682e-08, 6.459211e-08, 6.478453e-08, 6.421065e-08, 
    6.386559e-08, 6.363638e-08, 6.347373e-08, 6.349672e-08, 6.354056e-08, 
    6.376582e-08, 6.397759e-08, 6.413898e-08, 6.424694e-08, 6.435332e-08, 
    6.467531e-08, 6.484571e-08, 6.522728e-08, 6.515841e-08, 6.527507e-08, 
    6.538651e-08, 6.557362e-08, 6.554281e-08, 6.562525e-08, 6.527198e-08, 
    6.550677e-08, 6.511919e-08, 6.522519e-08, 6.438226e-08, 6.406108e-08, 
    6.392459e-08, 6.38051e-08, 6.351441e-08, 6.371515e-08, 6.363602e-08, 
    6.382428e-08, 6.394391e-08, 6.388474e-08, 6.42499e-08, 6.410793e-08, 
    6.485581e-08, 6.453368e-08, 6.537351e-08, 6.517254e-08, 6.542168e-08, 
    6.529455e-08, 6.551238e-08, 6.531634e-08, 6.565593e-08, 6.572988e-08, 
    6.567934e-08, 6.587345e-08, 6.530546e-08, 6.55236e-08, 6.388309e-08, 
    6.389273e-08, 6.393769e-08, 6.374008e-08, 6.372799e-08, 6.354689e-08, 
    6.370803e-08, 6.377665e-08, 6.395084e-08, 6.405388e-08, 6.415182e-08, 
    6.436717e-08, 6.460768e-08, 6.494398e-08, 6.518557e-08, 6.534752e-08, 
    6.524822e-08, 6.533589e-08, 6.523788e-08, 6.519194e-08, 6.570217e-08, 
    6.541567e-08, 6.584553e-08, 6.582174e-08, 6.562721e-08, 6.582443e-08, 
    6.389951e-08, 6.384398e-08, 6.365119e-08, 6.380206e-08, 6.352717e-08, 
    6.368104e-08, 6.376953e-08, 6.411091e-08, 6.41859e-08, 6.425545e-08, 
    6.439281e-08, 6.456909e-08, 6.487833e-08, 6.514738e-08, 6.539299e-08, 
    6.537499e-08, 6.538133e-08, 6.54362e-08, 6.530028e-08, 6.545852e-08, 
    6.548507e-08, 6.541563e-08, 6.581856e-08, 6.570345e-08, 6.582124e-08, 
    6.574629e-08, 6.386203e-08, 6.395546e-08, 6.390498e-08, 6.399992e-08, 
    6.393303e-08, 6.423046e-08, 6.431962e-08, 6.473687e-08, 6.456563e-08, 
    6.483815e-08, 6.45933e-08, 6.463669e-08, 6.484705e-08, 6.460653e-08, 
    6.513255e-08, 6.477594e-08, 6.543834e-08, 6.508223e-08, 6.546065e-08, 
    6.539193e-08, 6.55057e-08, 6.560761e-08, 6.57358e-08, 6.597234e-08, 
    6.591757e-08, 6.611538e-08, 6.409476e-08, 6.421595e-08, 6.420527e-08, 
    6.43321e-08, 6.44259e-08, 6.462918e-08, 6.495523e-08, 6.483262e-08, 
    6.505771e-08, 6.51029e-08, 6.476093e-08, 6.49709e-08, 6.429705e-08, 
    6.440593e-08, 6.43411e-08, 6.410432e-08, 6.486088e-08, 6.447262e-08, 
    6.518957e-08, 6.497923e-08, 6.559308e-08, 6.528781e-08, 6.588741e-08, 
    6.614376e-08, 6.638498e-08, 6.666692e-08, 6.428208e-08, 6.419974e-08, 
    6.434718e-08, 6.455118e-08, 6.474044e-08, 6.499207e-08, 6.501781e-08, 
    6.506495e-08, 6.518705e-08, 6.52897e-08, 6.507986e-08, 6.531544e-08, 
    6.443119e-08, 6.489459e-08, 6.416861e-08, 6.438723e-08, 6.453915e-08, 
    6.44725e-08, 6.481861e-08, 6.490018e-08, 6.523167e-08, 6.506031e-08, 
    6.60805e-08, 6.562914e-08, 6.688157e-08, 6.653157e-08, 6.417097e-08, 
    6.42818e-08, 6.466754e-08, 6.448401e-08, 6.500886e-08, 6.513805e-08, 
    6.524307e-08, 6.537733e-08, 6.539182e-08, 6.547136e-08, 6.534101e-08, 
    6.546621e-08, 6.49926e-08, 6.520425e-08, 6.462344e-08, 6.476481e-08, 
    6.469977e-08, 6.462844e-08, 6.48486e-08, 6.508316e-08, 6.508817e-08, 
    6.516338e-08, 6.537534e-08, 6.501099e-08, 6.613876e-08, 6.544229e-08, 
    6.440266e-08, 6.461615e-08, 6.464663e-08, 6.456393e-08, 6.51251e-08, 
    6.492177e-08, 6.546942e-08, 6.532141e-08, 6.556392e-08, 6.544342e-08, 
    6.542568e-08, 6.52709e-08, 6.517455e-08, 6.493109e-08, 6.473301e-08, 
    6.457592e-08, 6.461245e-08, 6.4785e-08, 6.509751e-08, 6.539313e-08, 
    6.532837e-08, 6.554549e-08, 6.497081e-08, 6.521179e-08, 6.511865e-08, 
    6.53615e-08, 6.482936e-08, 6.528253e-08, 6.471353e-08, 6.476342e-08, 
    6.491774e-08, 6.522814e-08, 6.52968e-08, 6.537012e-08, 6.532488e-08, 
    6.510544e-08, 6.506949e-08, 6.491398e-08, 6.487105e-08, 6.475256e-08, 
    6.465446e-08, 6.474409e-08, 6.483822e-08, 6.510553e-08, 6.534642e-08, 
    6.560906e-08, 6.567333e-08, 6.598021e-08, 6.57304e-08, 6.614265e-08, 
    6.579219e-08, 6.639884e-08, 6.530878e-08, 6.578186e-08, 6.492476e-08, 
    6.501709e-08, 6.518411e-08, 6.556716e-08, 6.536035e-08, 6.560221e-08, 
    6.506808e-08, 6.479096e-08, 6.471925e-08, 6.458548e-08, 6.472231e-08, 
    6.471118e-08, 6.484211e-08, 6.480003e-08, 6.511441e-08, 6.494554e-08, 
    6.542524e-08, 6.56003e-08, 6.609465e-08, 6.639771e-08, 6.670619e-08, 
    6.684238e-08, 6.688383e-08, 6.690116e-08 ;

 SOM_C_LEACHED =
  4.172668e-20, 2.750924e-20, 1.189856e-20, 5.877486e-20, 1.04472e-19, 
    7.595438e-20, -1.635496e-20, -2.524378e-20, 1.315887e-20, -7.086818e-20, 
    -3.005919e-20, -1.023792e-19, -2.966874e-21, 2.93304e-20, -3.208455e-20, 
    -2.74681e-20, -5.555858e-20, 4.373168e-20, 6.147027e-20, 2.085321e-20, 
    6.732506e-20, 8.391944e-21, 5.604515e-21, 5.394327e-20, 1.094892e-20, 
    2.900356e-20, -1.885039e-20, -1.031215e-20, 1.552561e-20, 3.55774e-20, 
    -1.223806e-20, 7.750026e-21, -4.404338e-20, -2.459556e-20, 1.970379e-20, 
    3.755412e-20, 2.910186e-20, 8.141574e-21, -7.174193e-20, 5.145777e-20, 
    -1.367022e-21, -3.922405e-20, 8.366962e-21, 4.858215e-20, 4.323555e-20, 
    2.469052e-20, 3.834084e-21, -1.609749e-20, 4.217389e-20, -8.919628e-21, 
    7.582116e-20, -4.021469e-21, 8.149819e-21, -6.389564e-21, 3.456095e-20, 
    -2.103239e-20, -1.489926e-20, 5.460325e-23, -2.397492e-20, 7.973549e-20, 
    5.996887e-21, -1.480831e-20, 4.735051e-22, -2.777373e-20, 5.037259e-20, 
    -4.140785e-20, 3.253018e-20, -3.195561e-20, 3.450796e-20, 4.85205e-20, 
    6.316777e-20, 9.925612e-20, -1.046742e-20, 8.196196e-20, 9.608168e-21, 
    -7.883415e-21, -1.297238e-21, -9.049799e-21, 2.963135e-21, -1.41671e-20, 
    -6.016175e-20, -3.400418e-20, 7.242881e-20, 5.559413e-20, 4.252663e-20, 
    1.64607e-20, -9.053774e-20, -5.937541e-22, -2.577919e-21, -2.428117e-20, 
    5.215131e-20, -2.961324e-20, -2.106327e-20, -5.935776e-20, 2.248151e-20, 
    -7.484787e-21, -3.752421e-20, 2.228632e-21, -1.13765e-20, 2.207038e-20, 
    -4.233705e-20, -2.018524e-20, -1.691586e-20, -3.85045e-21, -1.093293e-19, 
    5.257411e-20, -4.543077e-20, 3.517366e-20, -5.736715e-22, -2.204317e-20, 
    -1.129458e-20, 1.3584e-20, -4.788669e-20, -1.562811e-20, 7.505953e-20, 
    -1.123332e-20, -1.347956e-20, 2.587378e-20, 4.413468e-20, 2.409851e-20, 
    -1.011631e-20, 4.157261e-20, 6.496429e-20, -3.645009e-20, 8.231101e-21, 
    -5.323883e-20, 5.427689e-21, -2.074143e-20, -3.860831e-20, 1.753372e-20, 
    -4.24374e-20, 8.776877e-21, 5.410728e-21, -1.577525e-20, 3.539826e-20, 
    -3.676122e-20, -1.592459e-20, 1.700578e-20, 5.121628e-20, -2.525126e-20, 
    3.457789e-20, 3.207219e-20, -1.920387e-20, 2.602557e-21, 1.060548e-20, 
    5.255014e-22, -9.707794e-21, -5.04028e-20, -3.015215e-20, -1.01393e-20, 
    1.442175e-21, 5.917158e-20, 1.424551e-20, -2.539252e-20, 1.641216e-20, 
    -6.262229e-20, -4.447895e-20, 3.28543e-21, -2.590308e-21, 1.639659e-20, 
    1.166497e-20, 6.476177e-20, 2.270967e-20, 4.128278e-20, -1.149501e-22, 
    1.700327e-20, -9.521291e-21, -1.583039e-20, -2.73022e-21, -2.980284e-20, 
    -3.758554e-20, -1.85731e-21, -4.02884e-20, 4.670748e-22, 2.886346e-20, 
    3.714719e-20, -2.826952e-20, 3.79997e-20, 2.886894e-20, -5.724151e-21, 
    1.556024e-20, 1.090364e-19, -2.6666e-20, -7.188293e-20, -8.097746e-20, 
    -5.872302e-20, -1.506031e-20, -3.347449e-20, 5.232739e-21, 3.782222e-20, 
    1.075344e-20, 5.132369e-20, 1.447743e-20, -2.343941e-20, -4.250769e-20, 
    -1.386484e-20, 7.246628e-20, -1.671663e-20, 1.844126e-20, 1.977562e-20, 
    1.654558e-20, 8.592811e-21, -1.251593e-21, 7.52828e-21, -6.895e-20, 
    -3.305883e-20, -3.642677e-20, -8.46843e-20, 2.6309e-20, 3.328043e-21, 
    2.654006e-20, -1.044463e-20, 5.255487e-20, -3.816505e-21, -2.589256e-20, 
    -1.236298e-20, -4.291771e-20, 3.232525e-20, -9.940696e-21, 6.598884e-20, 
    3.51118e-20, 6.090281e-20, -2.853647e-21, -1.365004e-20, -9.115278e-21, 
    -8.486373e-21, 1.400518e-20, 9.476893e-21, 1.007898e-20, 4.424205e-20, 
    -5.134629e-20, -1.249332e-20, -1.989729e-20, 2.219033e-20, -4.991932e-20, 
    -2.421973e-20, -8.659539e-21, -8.849324e-21, 1.884872e-20, -5.408064e-20, 
    4.05214e-20, -2.537309e-20, -3.665104e-20, 5.892696e-20, -3.81124e-20, 
    -4.122564e-20, -1.352265e-20, -5.326275e-22, 2.939215e-20, -9.573474e-21, 
    9.048784e-21, 1.553833e-20, -7.860888e-21, 2.79622e-20, 4.648168e-20, 
    2.493775e-21, 3.398325e-20, -1.908337e-21, 6.375722e-21, 2.624556e-20, 
    -1.957796e-20, -1.312708e-20, -1.331018e-20, -3.777352e-20, 1.440295e-21, 
    -1.289033e-19, 1.875867e-20, 2.946462e-20, 3.798789e-21, -8.383429e-21, 
    -3.608149e-20, -2.491612e-20, 4.968096e-20, -1.619991e-21, -1.27387e-21, 
    -8.408436e-21, 6.378686e-21, -7.344179e-20, 6.416423e-21, 1.114509e-20, 
    3.877672e-20, -1.922895e-20, -1.929254e-20, 2.231761e-20, -3.206176e-20, 
    6.168897e-21, 9.163176e-21, -4.424281e-20, 5.219425e-20, 4.15561e-21, 
    3.558458e-20, -3.775072e-20, -4.765597e-21, 3.198314e-20, 7.519157e-20, 
    -2.418048e-20, -7.119145e-20, -6.650131e-21, 1.297459e-19, -4.372501e-20, 
    -4.240972e-20, -1.749503e-20, 6.619747e-21, -7.926776e-21, -7.936027e-20, 
    9.453118e-21, -2.243319e-21, -7.206351e-21, -2.686602e-20, 4.994185e-20, 
    5.297528e-20, 4.045616e-20, -6.77559e-20, 3.06663e-20, 2.962996e-20, 
    -2.709473e-20, 6.383182e-21, -4.979682e-21, 2.434642e-21, 1.237569e-19, 
    -5.390203e-20, -1.740731e-20, 1.875514e-20, 3.5526e-20, 4.745443e-21, 
    -3.231266e-20, -6.287616e-20, 1.874415e-20, 2.354357e-20, 8.409056e-20, 
    9.987844e-21, 4.267954e-21, 1.878327e-20, -6.977782e-20, 4.80332e-20, 
    4.91432e-20, -2.179538e-20, -1.701671e-20 ;

 SR =
  6.35703e-08, 6.384985e-08, 6.379551e-08, 6.402099e-08, 6.389591e-08, 
    6.404356e-08, 6.362697e-08, 6.386096e-08, 6.371158e-08, 6.359546e-08, 
    6.445858e-08, 6.403105e-08, 6.490264e-08, 6.462999e-08, 6.531489e-08, 
    6.486022e-08, 6.540657e-08, 6.530176e-08, 6.561717e-08, 6.552681e-08, 
    6.593026e-08, 6.565888e-08, 6.613939e-08, 6.586544e-08, 6.59083e-08, 
    6.564993e-08, 6.411708e-08, 6.440536e-08, 6.410001e-08, 6.414111e-08, 
    6.412267e-08, 6.38985e-08, 6.378554e-08, 6.354892e-08, 6.359188e-08, 
    6.376565e-08, 6.41596e-08, 6.402587e-08, 6.436288e-08, 6.435527e-08, 
    6.473046e-08, 6.45613e-08, 6.519191e-08, 6.501268e-08, 6.553059e-08, 
    6.540034e-08, 6.552447e-08, 6.548683e-08, 6.552496e-08, 6.533394e-08, 
    6.541578e-08, 6.524769e-08, 6.459298e-08, 6.47854e-08, 6.421152e-08, 
    6.386645e-08, 6.363724e-08, 6.347459e-08, 6.349758e-08, 6.354141e-08, 
    6.376668e-08, 6.397845e-08, 6.413985e-08, 6.424781e-08, 6.435418e-08, 
    6.467617e-08, 6.484658e-08, 6.522815e-08, 6.515928e-08, 6.527594e-08, 
    6.538738e-08, 6.557449e-08, 6.554369e-08, 6.562612e-08, 6.527286e-08, 
    6.550764e-08, 6.512006e-08, 6.522607e-08, 6.438312e-08, 6.406194e-08, 
    6.392545e-08, 6.380596e-08, 6.351526e-08, 6.371601e-08, 6.363688e-08, 
    6.382514e-08, 6.394477e-08, 6.38856e-08, 6.425076e-08, 6.41088e-08, 
    6.485669e-08, 6.453455e-08, 6.537438e-08, 6.517342e-08, 6.542255e-08, 
    6.529542e-08, 6.551326e-08, 6.531721e-08, 6.565681e-08, 6.573075e-08, 
    6.568022e-08, 6.587433e-08, 6.530634e-08, 6.552447e-08, 6.388395e-08, 
    6.389359e-08, 6.393855e-08, 6.374094e-08, 6.372885e-08, 6.354775e-08, 
    6.370889e-08, 6.377751e-08, 6.39517e-08, 6.405474e-08, 6.415268e-08, 
    6.436803e-08, 6.460854e-08, 6.494484e-08, 6.518644e-08, 6.53484e-08, 
    6.524908e-08, 6.533676e-08, 6.523875e-08, 6.519281e-08, 6.570305e-08, 
    6.541654e-08, 6.584641e-08, 6.582263e-08, 6.562809e-08, 6.58253e-08, 
    6.390037e-08, 6.384484e-08, 6.365205e-08, 6.380292e-08, 6.352803e-08, 
    6.36819e-08, 6.377039e-08, 6.411177e-08, 6.418676e-08, 6.425632e-08, 
    6.439367e-08, 6.456996e-08, 6.48792e-08, 6.514825e-08, 6.539386e-08, 
    6.537586e-08, 6.53822e-08, 6.543707e-08, 6.530116e-08, 6.545939e-08, 
    6.548594e-08, 6.541651e-08, 6.581944e-08, 6.570433e-08, 6.582212e-08, 
    6.574717e-08, 6.386289e-08, 6.395633e-08, 6.390584e-08, 6.400078e-08, 
    6.39339e-08, 6.423132e-08, 6.432049e-08, 6.473773e-08, 6.456649e-08, 
    6.483902e-08, 6.459417e-08, 6.463756e-08, 6.484792e-08, 6.46074e-08, 
    6.513343e-08, 6.477681e-08, 6.543921e-08, 6.508311e-08, 6.546152e-08, 
    6.53928e-08, 6.550658e-08, 6.560848e-08, 6.573668e-08, 6.597322e-08, 
    6.591844e-08, 6.611626e-08, 6.409562e-08, 6.421681e-08, 6.420614e-08, 
    6.433297e-08, 6.442676e-08, 6.463005e-08, 6.49561e-08, 6.483349e-08, 
    6.505858e-08, 6.510377e-08, 6.47618e-08, 6.497177e-08, 6.429792e-08, 
    6.44068e-08, 6.434197e-08, 6.410518e-08, 6.486175e-08, 6.447348e-08, 
    6.519043e-08, 6.498011e-08, 6.559395e-08, 6.528868e-08, 6.588829e-08, 
    6.614464e-08, 6.638587e-08, 6.66678e-08, 6.428295e-08, 6.42006e-08, 
    6.434804e-08, 6.455205e-08, 6.474131e-08, 6.499293e-08, 6.501867e-08, 
    6.506582e-08, 6.518791e-08, 6.529058e-08, 6.508073e-08, 6.531631e-08, 
    6.443206e-08, 6.489545e-08, 6.416948e-08, 6.438809e-08, 6.454002e-08, 
    6.447337e-08, 6.481947e-08, 6.490105e-08, 6.523254e-08, 6.506118e-08, 
    6.608137e-08, 6.563001e-08, 6.688245e-08, 6.653246e-08, 6.417183e-08, 
    6.428267e-08, 6.466841e-08, 6.448487e-08, 6.500973e-08, 6.513893e-08, 
    6.524394e-08, 6.53782e-08, 6.539269e-08, 6.547224e-08, 6.534189e-08, 
    6.546708e-08, 6.499347e-08, 6.520511e-08, 6.462431e-08, 6.476568e-08, 
    6.470064e-08, 6.46293e-08, 6.484947e-08, 6.508403e-08, 6.508903e-08, 
    6.516425e-08, 6.537621e-08, 6.501185e-08, 6.613964e-08, 6.544317e-08, 
    6.440352e-08, 6.461701e-08, 6.464749e-08, 6.456479e-08, 6.512597e-08, 
    6.492264e-08, 6.54703e-08, 6.532228e-08, 6.55648e-08, 6.544429e-08, 
    6.542655e-08, 6.527178e-08, 6.517542e-08, 6.493197e-08, 6.473388e-08, 
    6.457679e-08, 6.461332e-08, 6.478587e-08, 6.509838e-08, 6.5394e-08, 
    6.532925e-08, 6.554637e-08, 6.497167e-08, 6.521266e-08, 6.511952e-08, 
    6.536237e-08, 6.483023e-08, 6.528341e-08, 6.471441e-08, 6.476429e-08, 
    6.49186e-08, 6.522901e-08, 6.529767e-08, 6.5371e-08, 6.532575e-08, 
    6.510631e-08, 6.507035e-08, 6.491485e-08, 6.487192e-08, 6.475343e-08, 
    6.465533e-08, 6.474496e-08, 6.483909e-08, 6.51064e-08, 6.534729e-08, 
    6.560993e-08, 6.56742e-08, 6.598109e-08, 6.573129e-08, 6.614352e-08, 
    6.579306e-08, 6.639972e-08, 6.530966e-08, 6.578274e-08, 6.492562e-08, 
    6.501796e-08, 6.518498e-08, 6.556804e-08, 6.536123e-08, 6.560308e-08, 
    6.506895e-08, 6.479183e-08, 6.472012e-08, 6.458635e-08, 6.472317e-08, 
    6.471205e-08, 6.484298e-08, 6.480091e-08, 6.511527e-08, 6.494641e-08, 
    6.542611e-08, 6.560117e-08, 6.609553e-08, 6.639859e-08, 6.670707e-08, 
    6.684326e-08, 6.688472e-08, 6.690204e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 0.9999933, 
    0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999935, 0.9999933, 0.9999934, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 
    0.9999933, 0.9999933, 0.9999933, 0.9999932, 0.9999932, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999932, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 
    0.9999935, 0.9999935, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999934, 0.9999935, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999935, 0.9999936, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999932, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 
    0.9999936, 0.9999936, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999933, 0.9999934, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999933, 0.9999933, 
    0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999936, 0.9999935, 0.9999937, 0.9999936, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999935, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999937 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.147706, -0.1477211, -0.1477182, -0.1477302, -0.1477237, -0.1477314, 
    -0.1477091, -0.1477216, -0.1477137, -0.1477075, -0.1477518, -0.1477308, 
    -0.1477674, -0.1477586, -0.1477914, -0.1477659, -0.1477943, -0.1477912, 
    -0.147801, -0.1477982, -0.1478104, -0.1478023, -0.147817, -0.1478086, 
    -0.1478099, -0.147802, -0.1477353, -0.1477491, -0.1477344, -0.1477364, 
    -0.1477355, -0.1477237, -0.1477174, -0.147705, -0.1477073, -0.1477165, 
    -0.1477373, -0.1477307, -0.1477477, -0.1477474, -0.1477619, -0.1477563, 
    -0.1477878, -0.1477709, -0.1477984, -0.1477943, -0.1477981, -0.147797, 
    -0.1477982, -0.1477922, -0.1477947, -0.1477896, -0.1477574, -0.1477636, 
    -0.14774, -0.1477216, -0.1477097, -0.1477009, -0.1477022, -0.1477045, 
    -0.1477166, -0.1477281, -0.1477365, -0.1477419, -0.1477473, -0.1477598, 
    -0.1477655, -0.1477888, -0.1477868, -0.1477903, -0.1477939, -0.1477997, 
    -0.1477987, -0.1478013, -0.1477903, -0.1477975, -0.1477742, -0.1477889, 
    -0.1477479, -0.1477325, -0.1477249, -0.1477187, -0.1477031, -0.1477139, 
    -0.1477096, -0.1477199, -0.1477263, -0.1477232, -0.1477421, -0.1477349, 
    -0.1477659, -0.1477552, -0.1477935, -0.1477872, -0.147795, -0.1477911, 
    -0.1477977, -0.1477917, -0.1478022, -0.1478044, -0.1478029, -0.147809, 
    -0.1477914, -0.1477981, -0.147723, -0.1477236, -0.147726, -0.1477152, 
    -0.1477146, -0.1477049, -0.1477136, -0.1477172, -0.1477268, -0.1477321, 
    -0.1477371, -0.1477479, -0.1477578, -0.1477688, -0.1477876, -0.1477927, 
    -0.1477896, -0.1477923, -0.1477893, -0.1477879, -0.1478036, -0.1477947, 
    -0.1478081, -0.1478074, -0.1478013, -0.1478075, -0.1477239, -0.147721, 
    -0.1477105, -0.1477187, -0.1477038, -0.1477121, -0.1477167, -0.1477348, 
    -0.1477388, -0.1477423, -0.1477492, -0.1477566, -0.1477667, -0.1477864, 
    -0.1477941, -0.1477936, -0.1477938, -0.1477954, -0.1477912, -0.1477961, 
    -0.1477969, -0.1477948, -0.1478073, -0.1478037, -0.1478074, -0.1478051, 
    -0.147722, -0.147727, -0.1477242, -0.1477293, -0.1477257, -0.1477408, 
    -0.1477453, -0.147762, -0.1477564, -0.1477654, -0.1477574, -0.1477588, 
    -0.1477654, -0.1477579, -0.1477744, -0.1477632, -0.1477955, -0.1477727, 
    -0.1477962, -0.1477941, -0.1477976, -0.1478007, -0.1478047, -0.1478119, 
    -0.1478103, -0.1478164, -0.1477342, -0.1477402, -0.1477398, -0.1477462, 
    -0.1477508, -0.1477586, -0.1477692, -0.1477653, -0.1477723, -0.1477736, 
    -0.147763, -0.1477696, -0.1477443, -0.1477496, -0.1477466, -0.1477346, 
    -0.1477661, -0.1477529, -0.1477877, -0.1477699, -0.1478003, -0.1477907, 
    -0.1478094, -0.147817, -0.1478248, -0.1478333, -0.1477436, -0.1477395, 
    -0.147747, -0.1477558, -0.1477622, -0.1477703, -0.1477711, -0.1477725, 
    -0.1477877, -0.1477909, -0.1477728, -0.1477917, -0.1477505, -0.1477672, 
    -0.1477379, -0.1477486, -0.1477554, -0.147753, -0.1477649, -0.1477675, 
    -0.147789, -0.1477724, -0.1478151, -0.1478012, -0.1478401, -0.1478292, 
    -0.1477381, -0.1477437, -0.1477598, -0.1477534, -0.1477708, -0.1477747, 
    -0.1477895, -0.1477935, -0.1477941, -0.1477965, -0.1477925, -0.1477964, 
    -0.1477703, -0.1477882, -0.1477585, -0.147763, -0.147761, -0.1477586, 
    -0.1477658, -0.1477729, -0.1477732, -0.1477869, -0.1477929, -0.1477709, 
    -0.1478165, -0.1477951, -0.1477498, -0.147758, -0.1477592, -0.1477565, 
    -0.1477743, -0.1477682, -0.1477965, -0.1477919, -0.1477994, -0.1477957, 
    -0.1477951, -0.1477903, -0.1477873, -0.1477684, -0.147762, -0.1477569, 
    -0.1477581, -0.1477637, -0.1477734, -0.147794, -0.147792, -0.1477988, 
    -0.1477697, -0.1477884, -0.147774, -0.1477931, -0.1477652, -0.1477901, 
    -0.1477614, -0.1477631, -0.1477681, -0.1477888, -0.1477911, -0.1477933, 
    -0.147792, -0.1477736, -0.1477726, -0.147768, -0.1477665, -0.1477627, 
    -0.1477595, -0.1477624, -0.1477654, -0.1477737, -0.1477926, -0.1478007, 
    -0.1478028, -0.1478119, -0.1478042, -0.1478166, -0.1478057, -0.1478247, 
    -0.1477912, -0.1478058, -0.1477683, -0.1477711, -0.1477875, -0.1477993, 
    -0.1477931, -0.1478004, -0.1477726, -0.1477638, -0.1477616, -0.1477572, 
    -0.1477617, -0.1477613, -0.1477657, -0.1477643, -0.147774, -0.1477689, 
    -0.147795, -0.1478004, -0.1478157, -0.147825, -0.1478347, -0.1478389, 
    -0.1478402, -0.1478408 ;

 TAUY =
  -0.147706, -0.1477211, -0.1477182, -0.1477302, -0.1477237, -0.1477314, 
    -0.1477091, -0.1477216, -0.1477137, -0.1477075, -0.1477518, -0.1477308, 
    -0.1477674, -0.1477586, -0.1477914, -0.1477659, -0.1477943, -0.1477912, 
    -0.147801, -0.1477982, -0.1478104, -0.1478023, -0.147817, -0.1478086, 
    -0.1478099, -0.147802, -0.1477353, -0.1477491, -0.1477344, -0.1477364, 
    -0.1477355, -0.1477237, -0.1477174, -0.147705, -0.1477073, -0.1477165, 
    -0.1477373, -0.1477307, -0.1477477, -0.1477474, -0.1477619, -0.1477563, 
    -0.1477878, -0.1477709, -0.1477984, -0.1477943, -0.1477981, -0.147797, 
    -0.1477982, -0.1477922, -0.1477947, -0.1477896, -0.1477574, -0.1477636, 
    -0.14774, -0.1477216, -0.1477097, -0.1477009, -0.1477022, -0.1477045, 
    -0.1477166, -0.1477281, -0.1477365, -0.1477419, -0.1477473, -0.1477598, 
    -0.1477655, -0.1477888, -0.1477868, -0.1477903, -0.1477939, -0.1477997, 
    -0.1477987, -0.1478013, -0.1477903, -0.1477975, -0.1477742, -0.1477889, 
    -0.1477479, -0.1477325, -0.1477249, -0.1477187, -0.1477031, -0.1477139, 
    -0.1477096, -0.1477199, -0.1477263, -0.1477232, -0.1477421, -0.1477349, 
    -0.1477659, -0.1477552, -0.1477935, -0.1477872, -0.147795, -0.1477911, 
    -0.1477977, -0.1477917, -0.1478022, -0.1478044, -0.1478029, -0.147809, 
    -0.1477914, -0.1477981, -0.147723, -0.1477236, -0.147726, -0.1477152, 
    -0.1477146, -0.1477049, -0.1477136, -0.1477172, -0.1477268, -0.1477321, 
    -0.1477371, -0.1477479, -0.1477578, -0.1477688, -0.1477876, -0.1477927, 
    -0.1477896, -0.1477923, -0.1477893, -0.1477879, -0.1478036, -0.1477947, 
    -0.1478081, -0.1478074, -0.1478013, -0.1478075, -0.1477239, -0.147721, 
    -0.1477105, -0.1477187, -0.1477038, -0.1477121, -0.1477167, -0.1477348, 
    -0.1477388, -0.1477423, -0.1477492, -0.1477566, -0.1477667, -0.1477864, 
    -0.1477941, -0.1477936, -0.1477938, -0.1477954, -0.1477912, -0.1477961, 
    -0.1477969, -0.1477948, -0.1478073, -0.1478037, -0.1478074, -0.1478051, 
    -0.147722, -0.147727, -0.1477242, -0.1477293, -0.1477257, -0.1477408, 
    -0.1477453, -0.147762, -0.1477564, -0.1477654, -0.1477574, -0.1477588, 
    -0.1477654, -0.1477579, -0.1477744, -0.1477632, -0.1477955, -0.1477727, 
    -0.1477962, -0.1477941, -0.1477976, -0.1478007, -0.1478047, -0.1478119, 
    -0.1478103, -0.1478164, -0.1477342, -0.1477402, -0.1477398, -0.1477462, 
    -0.1477508, -0.1477586, -0.1477692, -0.1477653, -0.1477723, -0.1477736, 
    -0.147763, -0.1477696, -0.1477443, -0.1477496, -0.1477466, -0.1477346, 
    -0.1477661, -0.1477529, -0.1477877, -0.1477699, -0.1478003, -0.1477907, 
    -0.1478094, -0.147817, -0.1478248, -0.1478333, -0.1477436, -0.1477395, 
    -0.147747, -0.1477558, -0.1477622, -0.1477703, -0.1477711, -0.1477725, 
    -0.1477877, -0.1477909, -0.1477728, -0.1477917, -0.1477505, -0.1477672, 
    -0.1477379, -0.1477486, -0.1477554, -0.147753, -0.1477649, -0.1477675, 
    -0.147789, -0.1477724, -0.1478151, -0.1478012, -0.1478401, -0.1478292, 
    -0.1477381, -0.1477437, -0.1477598, -0.1477534, -0.1477708, -0.1477747, 
    -0.1477895, -0.1477935, -0.1477941, -0.1477965, -0.1477925, -0.1477964, 
    -0.1477703, -0.1477882, -0.1477585, -0.147763, -0.147761, -0.1477586, 
    -0.1477658, -0.1477729, -0.1477732, -0.1477869, -0.1477929, -0.1477709, 
    -0.1478165, -0.1477951, -0.1477498, -0.147758, -0.1477592, -0.1477565, 
    -0.1477743, -0.1477682, -0.1477965, -0.1477919, -0.1477994, -0.1477957, 
    -0.1477951, -0.1477903, -0.1477873, -0.1477684, -0.147762, -0.1477569, 
    -0.1477581, -0.1477637, -0.1477734, -0.147794, -0.147792, -0.1477988, 
    -0.1477697, -0.1477884, -0.147774, -0.1477931, -0.1477652, -0.1477901, 
    -0.1477614, -0.1477631, -0.1477681, -0.1477888, -0.1477911, -0.1477933, 
    -0.147792, -0.1477736, -0.1477726, -0.147768, -0.1477665, -0.1477627, 
    -0.1477595, -0.1477624, -0.1477654, -0.1477737, -0.1477926, -0.1478007, 
    -0.1478028, -0.1478119, -0.1478042, -0.1478166, -0.1478057, -0.1478247, 
    -0.1477912, -0.1478058, -0.1477683, -0.1477711, -0.1477875, -0.1477993, 
    -0.1477931, -0.1478004, -0.1477726, -0.1477638, -0.1477616, -0.1477572, 
    -0.1477617, -0.1477613, -0.1477657, -0.1477643, -0.147774, -0.1477689, 
    -0.147795, -0.1478004, -0.1478157, -0.147825, -0.1478347, -0.1478389, 
    -0.1478402, -0.1478408 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  262.7671, 262.781, 262.7783, 262.7896, 262.7833, 262.7907, 262.7699, 
    262.7816, 262.7741, 262.7684, 262.8113, 262.79, 262.8337, 262.82, 
    262.8542, 262.8315, 262.8589, 262.8536, 262.8695, 262.8649, 262.8852, 
    262.8716, 262.8957, 262.8819, 262.8841, 262.8711, 262.7943, 262.8087, 
    262.7935, 262.7955, 262.7946, 262.7834, 262.7778, 262.7661, 262.7682, 
    262.7768, 262.7965, 262.7898, 262.8066, 262.8062, 262.825, 262.8166, 
    262.8481, 262.8392, 262.8651, 262.8586, 262.8648, 262.8629, 262.8648, 
    262.8552, 262.8593, 262.8509, 262.8181, 262.8278, 262.7991, 262.7818, 
    262.7704, 262.7624, 262.7635, 262.7657, 262.7769, 262.7874, 262.7955, 
    262.8009, 262.8062, 262.8223, 262.8308, 262.8499, 262.8465, 262.8523, 
    262.8579, 262.8673, 262.8658, 262.8699, 262.8522, 262.864, 262.8446, 
    262.8498, 262.8076, 262.7916, 262.7848, 262.7788, 262.7644, 262.7744, 
    262.7704, 262.7798, 262.7858, 262.7828, 262.801, 262.7939, 262.8314, 
    262.8152, 262.8573, 262.8472, 262.8597, 262.8533, 262.8642, 262.8544, 
    262.8715, 262.8752, 262.8726, 262.8824, 262.8539, 262.8648, 262.7827, 
    262.7832, 262.7855, 262.7756, 262.775, 262.766, 262.774, 262.7774, 
    262.7861, 262.7913, 262.7961, 262.8069, 262.8189, 262.8358, 262.8478, 
    262.856, 262.851, 262.8554, 262.8505, 262.8481, 262.8738, 262.8594, 
    262.881, 262.8798, 262.87, 262.8799, 262.7835, 262.7808, 262.7712, 
    262.7787, 262.765, 262.7727, 262.7771, 262.7941, 262.7979, 262.8013, 
    262.8082, 262.817, 262.8325, 262.8459, 262.8582, 262.8573, 262.8577, 
    262.8604, 262.8536, 262.8615, 262.8629, 262.8594, 262.8796, 262.8738, 
    262.8798, 262.876, 262.7817, 262.7863, 262.7838, 262.7885, 262.7852, 
    262.8, 262.8045, 262.8254, 262.8168, 262.8305, 262.8182, 262.8204, 
    262.8309, 262.8189, 262.8453, 262.8273, 262.8605, 262.8427, 262.8616, 
    262.8582, 262.8639, 262.869, 262.8755, 262.8874, 262.8846, 262.8946, 
    262.7933, 262.7993, 262.7988, 262.8051, 262.8098, 262.82, 262.8364, 
    262.8302, 262.8415, 262.8438, 262.8266, 262.8372, 262.8034, 262.8088, 
    262.8056, 262.7938, 262.8316, 262.8121, 262.848, 262.8376, 262.8683, 
    262.8529, 262.8831, 262.8959, 262.9081, 262.9222, 262.8026, 262.7985, 
    262.8059, 262.8161, 262.8256, 262.8382, 262.8395, 262.8419, 262.8479, 
    262.8531, 262.8426, 262.8543, 262.81, 262.8333, 262.797, 262.8079, 
    262.8155, 262.8121, 262.8295, 262.8336, 262.8501, 262.8417, 262.8928, 
    262.8701, 262.9331, 262.9155, 262.7971, 262.8026, 262.8219, 262.8127, 
    262.8391, 262.8456, 262.8507, 262.8575, 262.8582, 262.8622, 262.8556, 
    262.8619, 262.8383, 262.8488, 262.8197, 262.8268, 262.8235, 262.82, 
    262.831, 262.8428, 262.843, 262.8467, 262.8573, 262.8392, 262.8956, 
    262.8607, 262.8087, 262.8193, 262.8209, 262.8167, 262.8449, 262.8347, 
    262.8621, 262.8546, 262.8669, 262.8608, 262.8599, 262.8521, 262.8473, 
    262.8351, 262.8252, 262.8174, 262.8192, 262.8278, 262.8435, 262.8582, 
    262.855, 262.8659, 262.8372, 262.8491, 262.8446, 262.8567, 262.83, 
    262.8526, 262.8242, 262.8268, 262.8345, 262.8499, 262.8534, 262.8571, 
    262.8548, 262.8439, 262.8421, 262.8343, 262.8322, 262.8262, 262.8213, 
    262.8258, 262.8305, 262.8439, 262.8559, 262.8691, 262.8723, 262.8877, 
    262.8752, 262.8958, 262.8782, 262.9088, 262.854, 262.8777, 262.8348, 
    262.8395, 262.8477, 262.867, 262.8566, 262.8687, 262.842, 262.8281, 
    262.8245, 262.8178, 262.8247, 262.8241, 262.8307, 262.8286, 262.8444, 
    262.8359, 262.8599, 262.8687, 262.8935, 262.9087, 262.9243, 262.9311, 
    262.9332, 262.9341 ;

 TG_R =
  262.7671, 262.781, 262.7783, 262.7896, 262.7833, 262.7907, 262.7699, 
    262.7816, 262.7741, 262.7684, 262.8113, 262.79, 262.8337, 262.82, 
    262.8542, 262.8315, 262.8589, 262.8536, 262.8695, 262.8649, 262.8852, 
    262.8716, 262.8957, 262.8819, 262.8841, 262.8711, 262.7943, 262.8087, 
    262.7935, 262.7955, 262.7946, 262.7834, 262.7778, 262.7661, 262.7682, 
    262.7768, 262.7965, 262.7898, 262.8066, 262.8062, 262.825, 262.8166, 
    262.8481, 262.8392, 262.8651, 262.8586, 262.8648, 262.8629, 262.8648, 
    262.8552, 262.8593, 262.8509, 262.8181, 262.8278, 262.7991, 262.7818, 
    262.7704, 262.7624, 262.7635, 262.7657, 262.7769, 262.7874, 262.7955, 
    262.8009, 262.8062, 262.8223, 262.8308, 262.8499, 262.8465, 262.8523, 
    262.8579, 262.8673, 262.8658, 262.8699, 262.8522, 262.864, 262.8446, 
    262.8498, 262.8076, 262.7916, 262.7848, 262.7788, 262.7644, 262.7744, 
    262.7704, 262.7798, 262.7858, 262.7828, 262.801, 262.7939, 262.8314, 
    262.8152, 262.8573, 262.8472, 262.8597, 262.8533, 262.8642, 262.8544, 
    262.8715, 262.8752, 262.8726, 262.8824, 262.8539, 262.8648, 262.7827, 
    262.7832, 262.7855, 262.7756, 262.775, 262.766, 262.774, 262.7774, 
    262.7861, 262.7913, 262.7961, 262.8069, 262.8189, 262.8358, 262.8478, 
    262.856, 262.851, 262.8554, 262.8505, 262.8481, 262.8738, 262.8594, 
    262.881, 262.8798, 262.87, 262.8799, 262.7835, 262.7808, 262.7712, 
    262.7787, 262.765, 262.7727, 262.7771, 262.7941, 262.7979, 262.8013, 
    262.8082, 262.817, 262.8325, 262.8459, 262.8582, 262.8573, 262.8577, 
    262.8604, 262.8536, 262.8615, 262.8629, 262.8594, 262.8796, 262.8738, 
    262.8798, 262.876, 262.7817, 262.7863, 262.7838, 262.7885, 262.7852, 
    262.8, 262.8045, 262.8254, 262.8168, 262.8305, 262.8182, 262.8204, 
    262.8309, 262.8189, 262.8453, 262.8273, 262.8605, 262.8427, 262.8616, 
    262.8582, 262.8639, 262.869, 262.8755, 262.8874, 262.8846, 262.8946, 
    262.7933, 262.7993, 262.7988, 262.8051, 262.8098, 262.82, 262.8364, 
    262.8302, 262.8415, 262.8438, 262.8266, 262.8372, 262.8034, 262.8088, 
    262.8056, 262.7938, 262.8316, 262.8121, 262.848, 262.8376, 262.8683, 
    262.8529, 262.8831, 262.8959, 262.9081, 262.9222, 262.8026, 262.7985, 
    262.8059, 262.8161, 262.8256, 262.8382, 262.8395, 262.8419, 262.8479, 
    262.8531, 262.8426, 262.8543, 262.81, 262.8333, 262.797, 262.8079, 
    262.8155, 262.8121, 262.8295, 262.8336, 262.8501, 262.8417, 262.8928, 
    262.8701, 262.9331, 262.9155, 262.7971, 262.8026, 262.8219, 262.8127, 
    262.8391, 262.8456, 262.8507, 262.8575, 262.8582, 262.8622, 262.8556, 
    262.8619, 262.8383, 262.8488, 262.8197, 262.8268, 262.8235, 262.82, 
    262.831, 262.8428, 262.843, 262.8467, 262.8573, 262.8392, 262.8956, 
    262.8607, 262.8087, 262.8193, 262.8209, 262.8167, 262.8449, 262.8347, 
    262.8621, 262.8546, 262.8669, 262.8608, 262.8599, 262.8521, 262.8473, 
    262.8351, 262.8252, 262.8174, 262.8192, 262.8278, 262.8435, 262.8582, 
    262.855, 262.8659, 262.8372, 262.8491, 262.8446, 262.8567, 262.83, 
    262.8526, 262.8242, 262.8268, 262.8345, 262.8499, 262.8534, 262.8571, 
    262.8548, 262.8439, 262.8421, 262.8343, 262.8322, 262.8262, 262.8213, 
    262.8258, 262.8305, 262.8439, 262.8559, 262.8691, 262.8723, 262.8877, 
    262.8752, 262.8958, 262.8782, 262.9088, 262.854, 262.8777, 262.8348, 
    262.8395, 262.8477, 262.867, 262.8566, 262.8687, 262.842, 262.8281, 
    262.8245, 262.8178, 262.8247, 262.8241, 262.8307, 262.8286, 262.8444, 
    262.8359, 262.8599, 262.8687, 262.8935, 262.9087, 262.9243, 262.9311, 
    262.9332, 262.9341 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  255.001, 255.0005, 255.0006, 255.0003, 255.0005, 255.0002, 255.0009, 
    255.0005, 255.0008, 255.0009, 254.9996, 255.0003, 254.999, 254.9994, 
    254.9985, 254.9991, 254.9984, 254.9985, 254.9981, 254.9982, 254.9977, 
    254.9981, 254.9975, 254.9978, 254.9977, 254.9981, 255.0001, 254.9997, 
    255.0002, 255.0001, 255.0001, 255.0005, 255.0006, 255.001, 255.0009, 
    255.0007, 255.0001, 255.0003, 254.9998, 254.9998, 254.9993, 254.9995, 
    254.9986, 254.9989, 254.9982, 254.9984, 254.9982, 254.9983, 254.9982, 
    254.9985, 254.9984, 254.9986, 254.9995, 254.9992, 255, 255.0005, 
    255.0009, 255.0011, 255.0011, 255.001, 255.0007, 255.0004, 255.0001, 255, 
    254.9998, 254.9993, 254.9991, 254.9986, 254.9987, 254.9985, 254.9984, 
    254.9982, 254.9982, 254.9981, 254.9985, 254.9982, 254.9987, 254.9986, 
    254.9997, 255.0002, 255.0004, 255.0006, 255.0011, 255.0007, 255.0009, 
    255.0006, 255.0004, 255.0005, 255, 255.0002, 254.9991, 254.9995, 
    254.9984, 254.9987, 254.9984, 254.9985, 254.9982, 254.9985, 254.9981, 
    254.998, 254.998, 254.9978, 254.9985, 254.9982, 255.0005, 255.0005, 
    255.0004, 255.0007, 255.0007, 255.001, 255.0008, 255.0007, 255.0004, 
    255.0002, 255.0001, 254.9998, 254.9994, 254.999, 254.9986, 254.9984, 
    254.9986, 254.9985, 254.9986, 254.9986, 254.998, 254.9984, 254.9978, 
    254.9978, 254.9981, 254.9978, 255.0005, 255.0006, 255.0009, 255.0006, 
    255.0011, 255.0008, 255.0007, 255.0001, 255, 254.9999, 254.9997, 
    254.9995, 254.9991, 254.9987, 254.9984, 254.9984, 254.9984, 254.9983, 
    254.9985, 254.9983, 254.9983, 254.9984, 254.9979, 254.998, 254.9978, 
    254.998, 255.0005, 255.0004, 255.0005, 255.0003, 255.0004, 255, 254.9998, 
    254.9992, 254.9995, 254.9991, 254.9995, 254.9994, 254.9991, 254.9994, 
    254.9987, 254.9992, 254.9983, 254.9988, 254.9983, 254.9984, 254.9982, 
    254.9981, 254.998, 254.9977, 254.9977, 254.9975, 255.0002, 255, 255, 
    254.9998, 254.9997, 254.9994, 254.999, 254.9991, 254.9988, 254.9988, 
    254.9992, 254.9989, 254.9999, 254.9997, 254.9998, 255.0002, 254.9991, 
    254.9996, 254.9986, 254.9989, 254.9981, 254.9985, 254.9978, 254.9974, 
    254.9972, 254.9968, 254.9999, 255, 254.9998, 254.9995, 254.9993, 
    254.9989, 254.9989, 254.9988, 254.9986, 254.9985, 254.9988, 254.9985, 
    254.9996, 254.999, 255.0001, 254.9997, 254.9995, 254.9996, 254.9991, 
    254.999, 254.9986, 254.9988, 254.9975, 254.9981, 254.9966, 254.997, 
    255.0001, 254.9999, 254.9993, 254.9996, 254.9989, 254.9987, 254.9986, 
    254.9984, 254.9984, 254.9983, 254.9985, 254.9983, 254.9989, 254.9986, 
    254.9994, 254.9992, 254.9993, 254.9994, 254.9991, 254.9988, 254.9988, 
    254.9987, 254.9983, 254.9989, 254.9974, 254.9983, 254.9997, 254.9994, 
    254.9994, 254.9995, 254.9987, 254.999, 254.9983, 254.9985, 254.9982, 
    254.9983, 254.9983, 254.9985, 254.9987, 254.999, 254.9993, 254.9995, 
    254.9994, 254.9992, 254.9988, 254.9984, 254.9985, 254.9982, 254.9989, 
    254.9986, 254.9987, 254.9984, 254.9991, 254.9985, 254.9993, 254.9992, 
    254.999, 254.9986, 254.9985, 254.9984, 254.9985, 254.9988, 254.9988, 
    254.999, 254.9991, 254.9992, 254.9994, 254.9993, 254.9991, 254.9988, 
    254.9984, 254.9981, 254.998, 254.9976, 254.9979, 254.9974, 254.9978, 
    254.9971, 254.9985, 254.9979, 254.999, 254.9989, 254.9986, 254.9981, 
    254.9984, 254.9981, 254.9988, 254.9992, 254.9993, 254.9995, 254.9993, 
    254.9993, 254.9991, 254.9992, 254.9987, 254.999, 254.9983, 254.9981, 
    254.9975, 254.9971, 254.9968, 254.9966, 254.9966, 254.9966 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTCOLCH4 =
  1.384293e-05, 1.363263e-05, 1.367344e-05, 1.350439e-05, 1.359809e-05, 
    1.348751e-05, 1.380023e-05, 1.36243e-05, 1.373653e-05, 1.382397e-05, 
    1.31784e-05, 1.349687e-05, 1.285096e-05, 1.30516e-05, 1.263902e-05, 
    1.288208e-05, 1.256842e-05, 1.264917e-05, 1.240743e-05, 1.24763e-05, 
    1.217138e-05, 1.237576e-05, 1.201605e-05, 1.221992e-05, 1.218781e-05, 
    1.238255e-05, 1.343257e-05, 1.321788e-05, 1.344533e-05, 1.341462e-05, 
    1.34284e-05, 1.359615e-05, 1.368093e-05, 1.385905e-05, 1.382667e-05, 
    1.369587e-05, 1.340083e-05, 1.350075e-05, 1.324947e-05, 1.325513e-05, 
    1.29775e-05, 1.310237e-05, 1.273425e-05, 1.287398e-05, 1.247342e-05, 
    1.257321e-05, 1.247809e-05, 1.250687e-05, 1.247771e-05, 1.262434e-05, 
    1.256134e-05, 1.269099e-05, 1.307894e-05, 1.293706e-05, 1.336211e-05, 
    1.362017e-05, 1.379249e-05, 1.391515e-05, 1.389779e-05, 1.386471e-05, 
    1.369511e-05, 1.353624e-05, 1.341558e-05, 1.333508e-05, 1.325594e-05, 
    1.301749e-05, 1.289209e-05, 1.270612e-05, 1.27596e-05, 1.266912e-05, 
    1.258318e-05, 1.243992e-05, 1.246341e-05, 1.240063e-05, 1.267151e-05, 
    1.249094e-05, 1.279013e-05, 1.270775e-05, 1.323439e-05, 1.347377e-05, 
    1.357593e-05, 1.366559e-05, 1.388445e-05, 1.37332e-05, 1.379276e-05, 
    1.36512e-05, 1.356147e-05, 1.360583e-05, 1.333288e-05, 1.343876e-05, 
    1.288468e-05, 1.312216e-05, 1.259318e-05, 1.274861e-05, 1.255615e-05, 
    1.265407e-05, 1.248665e-05, 1.263725e-05, 1.237733e-05, 1.232133e-05, 
    1.235958e-05, 1.221327e-05, 1.264564e-05, 1.247808e-05, 1.360707e-05, 
    1.359983e-05, 1.356613e-05, 1.371445e-05, 1.372354e-05, 1.385994e-05, 
    1.373856e-05, 1.368696e-05, 1.355628e-05, 1.347916e-05, 1.340599e-05, 
    1.324564e-05, 1.306744e-05, 1.282004e-05, 1.273849e-05, 1.26132e-05, 
    1.268991e-05, 1.262216e-05, 1.269792e-05, 1.273355e-05, 1.234229e-05, 
    1.256075e-05, 1.223421e-05, 1.225209e-05, 1.239913e-05, 1.225007e-05, 
    1.359475e-05, 1.363641e-05, 1.378134e-05, 1.366788e-05, 1.387482e-05, 
    1.375886e-05, 1.369231e-05, 1.343653e-05, 1.338057e-05, 1.332873e-05, 
    1.32266e-05, 1.309596e-05, 1.286816e-05, 1.276817e-05, 1.257819e-05, 
    1.259204e-05, 1.258716e-05, 1.2545e-05, 1.264964e-05, 1.252789e-05, 
    1.250754e-05, 1.256079e-05, 1.225448e-05, 1.234133e-05, 1.225247e-05, 
    1.230894e-05, 1.362286e-05, 1.355281e-05, 1.359065e-05, 1.351952e-05, 
    1.356961e-05, 1.334735e-05, 1.328097e-05, 1.297213e-05, 1.309853e-05, 
    1.289765e-05, 1.307806e-05, 1.304601e-05, 1.28911e-05, 1.306829e-05, 
    1.27797e-05, 1.294337e-05, 1.254336e-05, 1.281891e-05, 1.252625e-05, 
    1.257901e-05, 1.249176e-05, 1.241404e-05, 1.231687e-05, 1.213933e-05, 
    1.218023e-05, 1.203314e-05, 1.344861e-05, 1.335816e-05, 1.336613e-05, 
    1.327171e-05, 1.320204e-05, 1.305156e-05, 1.28118e-05, 1.290172e-05, 
    1.283809e-05, 1.280282e-05, 1.295443e-05, 1.280033e-05, 1.329777e-05, 
    1.321684e-05, 1.326501e-05, 1.344146e-05, 1.288096e-05, 1.316738e-05, 
    1.273539e-05, 1.279423e-05, 1.24251e-05, 1.265927e-05, 1.22028e-05, 
    1.201216e-05, 1.183549e-05, 1.163243e-05, 1.330891e-05, 1.337025e-05, 
    1.32605e-05, 1.31092e-05, 1.296951e-05, 1.278485e-05, 1.286928e-05, 
    1.283243e-05, 1.273735e-05, 1.265782e-05, 1.282078e-05, 1.263794e-05, 
    1.319808e-05, 1.285624e-05, 1.339346e-05, 1.323073e-05, 1.311811e-05, 
    1.316747e-05, 1.291202e-05, 1.285214e-05, 1.270272e-05, 1.283606e-05, 
    1.205894e-05, 1.239766e-05, 1.14805e-05, 1.172943e-05, 1.339171e-05, 
    1.330912e-05, 1.302324e-05, 1.315895e-05, 1.287628e-05, 1.277543e-05, 
    1.26939e-05, 1.259024e-05, 1.25791e-05, 1.251804e-05, 1.261821e-05, 
    1.252199e-05, 1.278446e-05, 1.272399e-05, 1.30558e-05, 1.295158e-05, 
    1.299948e-05, 1.305211e-05, 1.288999e-05, 1.28182e-05, 1.281431e-05, 
    1.275573e-05, 1.259172e-05, 1.287462e-05, 1.201582e-05, 1.254029e-05, 
    1.321929e-05, 1.306117e-05, 1.303868e-05, 1.309978e-05, 1.278552e-05, 
    1.283631e-05, 1.251953e-05, 1.263333e-05, 1.244731e-05, 1.253947e-05, 
    1.255307e-05, 1.267235e-05, 1.274705e-05, 1.282948e-05, 1.297499e-05, 
    1.309092e-05, 1.306392e-05, 1.293672e-05, 1.280701e-05, 1.257808e-05, 
    1.262795e-05, 1.246137e-05, 1.280041e-05, 1.271814e-05, 1.279054e-05, 
    1.260243e-05, 1.290411e-05, 1.266332e-05, 1.298934e-05, 1.29526e-05, 
    1.283927e-05, 1.270545e-05, 1.265234e-05, 1.259578e-05, 1.263066e-05, 
    1.280083e-05, 1.282888e-05, 1.284202e-05, 1.28735e-05, 1.29606e-05, 
    1.30329e-05, 1.296683e-05, 1.28976e-05, 1.280077e-05, 1.261404e-05, 
    1.241294e-05, 1.236414e-05, 1.213344e-05, 1.232092e-05, 1.201295e-05, 
    1.227428e-05, 1.182538e-05, 1.264306e-05, 1.228209e-05, 1.283413e-05, 
    1.286984e-05, 1.273961e-05, 1.244483e-05, 1.260331e-05, 1.241814e-05, 
    1.282999e-05, 1.293233e-05, 1.298513e-05, 1.308385e-05, 1.298287e-05, 
    1.299107e-05, 1.289475e-05, 1.292567e-05, 1.279385e-05, 1.28189e-05, 
    1.255341e-05, 1.24196e-05, 1.204847e-05, 1.182623e-05, 1.160448e-05, 
    1.150807e-05, 1.147892e-05, 1.146675e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976207e-05, 5.976193e-05, 5.976195e-05, 5.976183e-05, 5.97619e-05, 
    5.976182e-05, 5.976204e-05, 5.976192e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976183e-05, 5.976138e-05, 5.976152e-05, 5.976116e-05, 
    5.97614e-05, 5.976111e-05, 5.976117e-05, 5.976101e-05, 5.976105e-05, 
    5.976085e-05, 5.976098e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976178e-05, 5.976163e-05, 5.976179e-05, 5.976177e-05, 
    5.976178e-05, 5.97619e-05, 5.976196e-05, 5.976208e-05, 5.976206e-05, 
    5.976197e-05, 5.976176e-05, 5.976183e-05, 5.976166e-05, 5.976166e-05, 
    5.976147e-05, 5.976155e-05, 5.976123e-05, 5.976132e-05, 5.976105e-05, 
    5.976112e-05, 5.976105e-05, 5.976107e-05, 5.976105e-05, 5.976115e-05, 
    5.976111e-05, 5.97612e-05, 5.976154e-05, 5.976144e-05, 5.976174e-05, 
    5.976191e-05, 5.976203e-05, 5.976212e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976177e-05, 5.976172e-05, 5.976166e-05, 
    5.976149e-05, 5.976141e-05, 5.976121e-05, 5.976124e-05, 5.976118e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.9761e-05, 5.976118e-05, 
    5.976106e-05, 5.976126e-05, 5.976121e-05, 5.976165e-05, 5.976181e-05, 
    5.976189e-05, 5.976195e-05, 5.97621e-05, 5.976199e-05, 5.976203e-05, 
    5.976194e-05, 5.976187e-05, 5.976191e-05, 5.976171e-05, 5.976179e-05, 
    5.97614e-05, 5.976157e-05, 5.976113e-05, 5.976123e-05, 5.976111e-05, 
    5.976117e-05, 5.976106e-05, 5.976116e-05, 5.976098e-05, 5.976095e-05, 
    5.976097e-05, 5.976087e-05, 5.976117e-05, 5.976105e-05, 5.976191e-05, 
    5.97619e-05, 5.976188e-05, 5.976198e-05, 5.976199e-05, 5.976208e-05, 
    5.9762e-05, 5.976196e-05, 5.976187e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976153e-05, 5.976135e-05, 5.976123e-05, 5.976114e-05, 
    5.97612e-05, 5.976115e-05, 5.97612e-05, 5.976123e-05, 5.976096e-05, 
    5.976111e-05, 5.976089e-05, 5.97609e-05, 5.9761e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976171e-05, 
    5.976164e-05, 5.976155e-05, 5.976139e-05, 5.976125e-05, 5.976112e-05, 
    5.976113e-05, 5.976113e-05, 5.97611e-05, 5.976117e-05, 5.976109e-05, 
    5.976107e-05, 5.976111e-05, 5.97609e-05, 5.976096e-05, 5.97609e-05, 
    5.976094e-05, 5.976192e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976188e-05, 5.976173e-05, 5.976168e-05, 5.976146e-05, 5.976155e-05, 
    5.976141e-05, 5.976154e-05, 5.976151e-05, 5.976141e-05, 5.976153e-05, 
    5.976126e-05, 5.976144e-05, 5.97611e-05, 5.976128e-05, 5.976109e-05, 
    5.976112e-05, 5.976106e-05, 5.976101e-05, 5.976094e-05, 5.976082e-05, 
    5.976085e-05, 5.976075e-05, 5.97618e-05, 5.976173e-05, 5.976174e-05, 
    5.976167e-05, 5.976162e-05, 5.976152e-05, 5.976135e-05, 5.976141e-05, 
    5.97613e-05, 5.976127e-05, 5.976145e-05, 5.976134e-05, 5.976169e-05, 
    5.976163e-05, 5.976167e-05, 5.976179e-05, 5.97614e-05, 5.97616e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976073e-05, 5.976061e-05, 5.976046e-05, 5.97617e-05, 5.976174e-05, 
    5.976166e-05, 5.976156e-05, 5.976146e-05, 5.976133e-05, 5.976131e-05, 
    5.976129e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976116e-05, 
    5.976162e-05, 5.976138e-05, 5.976176e-05, 5.976165e-05, 5.976157e-05, 
    5.97616e-05, 5.976142e-05, 5.976138e-05, 5.976121e-05, 5.976129e-05, 
    5.976076e-05, 5.9761e-05, 5.976035e-05, 5.976053e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.976159e-05, 5.976132e-05, 5.976125e-05, 
    5.97612e-05, 5.976113e-05, 5.976112e-05, 5.976108e-05, 5.976115e-05, 
    5.976109e-05, 5.976133e-05, 5.976122e-05, 5.976152e-05, 5.976145e-05, 
    5.976148e-05, 5.976152e-05, 5.976141e-05, 5.976128e-05, 5.976128e-05, 
    5.976124e-05, 5.976113e-05, 5.976132e-05, 5.976074e-05, 5.97611e-05, 
    5.976163e-05, 5.976153e-05, 5.976151e-05, 5.976155e-05, 5.976126e-05, 
    5.976137e-05, 5.976108e-05, 5.976116e-05, 5.976103e-05, 5.97611e-05, 
    5.97611e-05, 5.976118e-05, 5.976123e-05, 5.976136e-05, 5.976146e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976127e-05, 5.976112e-05, 
    5.976115e-05, 5.976104e-05, 5.976134e-05, 5.976122e-05, 5.976126e-05, 
    5.976114e-05, 5.976141e-05, 5.976118e-05, 5.976147e-05, 5.976145e-05, 
    5.976137e-05, 5.976121e-05, 5.976117e-05, 5.976113e-05, 5.976116e-05, 
    5.976127e-05, 5.976129e-05, 5.976137e-05, 5.976139e-05, 5.976145e-05, 
    5.97615e-05, 5.976146e-05, 5.976141e-05, 5.976127e-05, 5.976115e-05, 
    5.976101e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976073e-05, 
    5.976091e-05, 5.97606e-05, 5.976117e-05, 5.976092e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976103e-05, 5.976114e-05, 5.976101e-05, 
    5.976129e-05, 5.976143e-05, 5.976147e-05, 5.976154e-05, 5.976147e-05, 
    5.976147e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976135e-05, 
    5.97611e-05, 5.976101e-05, 5.976076e-05, 5.97606e-05, 5.976044e-05, 
    5.976037e-05, 5.976035e-05, 5.976034e-05 ;

 TOTLITC_1m =
  5.976207e-05, 5.976193e-05, 5.976195e-05, 5.976183e-05, 5.97619e-05, 
    5.976182e-05, 5.976204e-05, 5.976192e-05, 5.9762e-05, 5.976206e-05, 
    5.976161e-05, 5.976183e-05, 5.976138e-05, 5.976152e-05, 5.976116e-05, 
    5.97614e-05, 5.976111e-05, 5.976117e-05, 5.976101e-05, 5.976105e-05, 
    5.976085e-05, 5.976098e-05, 5.976074e-05, 5.976088e-05, 5.976086e-05, 
    5.976099e-05, 5.976178e-05, 5.976163e-05, 5.976179e-05, 5.976177e-05, 
    5.976178e-05, 5.97619e-05, 5.976196e-05, 5.976208e-05, 5.976206e-05, 
    5.976197e-05, 5.976176e-05, 5.976183e-05, 5.976166e-05, 5.976166e-05, 
    5.976147e-05, 5.976155e-05, 5.976123e-05, 5.976132e-05, 5.976105e-05, 
    5.976112e-05, 5.976105e-05, 5.976107e-05, 5.976105e-05, 5.976115e-05, 
    5.976111e-05, 5.97612e-05, 5.976154e-05, 5.976144e-05, 5.976174e-05, 
    5.976191e-05, 5.976203e-05, 5.976212e-05, 5.976211e-05, 5.976209e-05, 
    5.976197e-05, 5.976186e-05, 5.976177e-05, 5.976172e-05, 5.976166e-05, 
    5.976149e-05, 5.976141e-05, 5.976121e-05, 5.976124e-05, 5.976118e-05, 
    5.976113e-05, 5.976103e-05, 5.976105e-05, 5.9761e-05, 5.976118e-05, 
    5.976106e-05, 5.976126e-05, 5.976121e-05, 5.976165e-05, 5.976181e-05, 
    5.976189e-05, 5.976195e-05, 5.97621e-05, 5.976199e-05, 5.976203e-05, 
    5.976194e-05, 5.976187e-05, 5.976191e-05, 5.976171e-05, 5.976179e-05, 
    5.97614e-05, 5.976157e-05, 5.976113e-05, 5.976123e-05, 5.976111e-05, 
    5.976117e-05, 5.976106e-05, 5.976116e-05, 5.976098e-05, 5.976095e-05, 
    5.976097e-05, 5.976087e-05, 5.976117e-05, 5.976105e-05, 5.976191e-05, 
    5.97619e-05, 5.976188e-05, 5.976198e-05, 5.976199e-05, 5.976208e-05, 
    5.9762e-05, 5.976196e-05, 5.976187e-05, 5.976182e-05, 5.976177e-05, 
    5.976166e-05, 5.976153e-05, 5.976135e-05, 5.976123e-05, 5.976114e-05, 
    5.97612e-05, 5.976115e-05, 5.97612e-05, 5.976123e-05, 5.976096e-05, 
    5.976111e-05, 5.976089e-05, 5.97609e-05, 5.9761e-05, 5.97609e-05, 
    5.97619e-05, 5.976193e-05, 5.976203e-05, 5.976195e-05, 5.976209e-05, 
    5.976201e-05, 5.976197e-05, 5.976179e-05, 5.976175e-05, 5.976171e-05, 
    5.976164e-05, 5.976155e-05, 5.976139e-05, 5.976125e-05, 5.976112e-05, 
    5.976113e-05, 5.976113e-05, 5.97611e-05, 5.976117e-05, 5.976109e-05, 
    5.976107e-05, 5.976111e-05, 5.97609e-05, 5.976096e-05, 5.97609e-05, 
    5.976094e-05, 5.976192e-05, 5.976187e-05, 5.97619e-05, 5.976185e-05, 
    5.976188e-05, 5.976173e-05, 5.976168e-05, 5.976146e-05, 5.976155e-05, 
    5.976141e-05, 5.976154e-05, 5.976151e-05, 5.976141e-05, 5.976153e-05, 
    5.976126e-05, 5.976144e-05, 5.97611e-05, 5.976128e-05, 5.976109e-05, 
    5.976112e-05, 5.976106e-05, 5.976101e-05, 5.976094e-05, 5.976082e-05, 
    5.976085e-05, 5.976075e-05, 5.97618e-05, 5.976173e-05, 5.976174e-05, 
    5.976167e-05, 5.976162e-05, 5.976152e-05, 5.976135e-05, 5.976141e-05, 
    5.97613e-05, 5.976127e-05, 5.976145e-05, 5.976134e-05, 5.976169e-05, 
    5.976163e-05, 5.976167e-05, 5.976179e-05, 5.97614e-05, 5.97616e-05, 
    5.976123e-05, 5.976134e-05, 5.976102e-05, 5.976118e-05, 5.976087e-05, 
    5.976073e-05, 5.976061e-05, 5.976046e-05, 5.97617e-05, 5.976174e-05, 
    5.976166e-05, 5.976156e-05, 5.976146e-05, 5.976133e-05, 5.976131e-05, 
    5.976129e-05, 5.976123e-05, 5.976118e-05, 5.976129e-05, 5.976116e-05, 
    5.976162e-05, 5.976138e-05, 5.976176e-05, 5.976165e-05, 5.976157e-05, 
    5.97616e-05, 5.976142e-05, 5.976138e-05, 5.976121e-05, 5.976129e-05, 
    5.976076e-05, 5.9761e-05, 5.976035e-05, 5.976053e-05, 5.976176e-05, 
    5.97617e-05, 5.97615e-05, 5.976159e-05, 5.976132e-05, 5.976125e-05, 
    5.97612e-05, 5.976113e-05, 5.976112e-05, 5.976108e-05, 5.976115e-05, 
    5.976109e-05, 5.976133e-05, 5.976122e-05, 5.976152e-05, 5.976145e-05, 
    5.976148e-05, 5.976152e-05, 5.976141e-05, 5.976128e-05, 5.976128e-05, 
    5.976124e-05, 5.976113e-05, 5.976132e-05, 5.976074e-05, 5.97611e-05, 
    5.976163e-05, 5.976153e-05, 5.976151e-05, 5.976155e-05, 5.976126e-05, 
    5.976137e-05, 5.976108e-05, 5.976116e-05, 5.976103e-05, 5.97611e-05, 
    5.97611e-05, 5.976118e-05, 5.976123e-05, 5.976136e-05, 5.976146e-05, 
    5.976155e-05, 5.976153e-05, 5.976144e-05, 5.976127e-05, 5.976112e-05, 
    5.976115e-05, 5.976104e-05, 5.976134e-05, 5.976122e-05, 5.976126e-05, 
    5.976114e-05, 5.976141e-05, 5.976118e-05, 5.976147e-05, 5.976145e-05, 
    5.976137e-05, 5.976121e-05, 5.976117e-05, 5.976113e-05, 5.976116e-05, 
    5.976127e-05, 5.976129e-05, 5.976137e-05, 5.976139e-05, 5.976145e-05, 
    5.97615e-05, 5.976146e-05, 5.976141e-05, 5.976127e-05, 5.976115e-05, 
    5.976101e-05, 5.976098e-05, 5.976082e-05, 5.976095e-05, 5.976073e-05, 
    5.976091e-05, 5.97606e-05, 5.976117e-05, 5.976092e-05, 5.976137e-05, 
    5.976132e-05, 5.976123e-05, 5.976103e-05, 5.976114e-05, 5.976101e-05, 
    5.976129e-05, 5.976143e-05, 5.976147e-05, 5.976154e-05, 5.976147e-05, 
    5.976147e-05, 5.976141e-05, 5.976143e-05, 5.976127e-05, 5.976135e-05, 
    5.97611e-05, 5.976101e-05, 5.976076e-05, 5.97606e-05, 5.976044e-05, 
    5.976037e-05, 5.976035e-05, 5.976034e-05 ;

 TOTLITN =
  1.37593e-06, 1.375926e-06, 1.375927e-06, 1.375923e-06, 1.375925e-06, 
    1.375923e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 1.37593e-06, 
    1.375917e-06, 1.375923e-06, 1.375911e-06, 1.375915e-06, 1.375905e-06, 
    1.375911e-06, 1.375903e-06, 1.375905e-06, 1.3759e-06, 1.375902e-06, 
    1.375896e-06, 1.3759e-06, 1.375893e-06, 1.375897e-06, 1.375896e-06, 
    1.3759e-06, 1.375922e-06, 1.375918e-06, 1.375922e-06, 1.375922e-06, 
    1.375922e-06, 1.375925e-06, 1.375927e-06, 1.37593e-06, 1.37593e-06, 
    1.375927e-06, 1.375922e-06, 1.375923e-06, 1.375918e-06, 1.375919e-06, 
    1.375913e-06, 1.375916e-06, 1.375906e-06, 1.375909e-06, 1.375901e-06, 
    1.375903e-06, 1.375902e-06, 1.375902e-06, 1.375902e-06, 1.375904e-06, 
    1.375903e-06, 1.375906e-06, 1.375915e-06, 1.375912e-06, 1.375921e-06, 
    1.375926e-06, 1.375929e-06, 1.375932e-06, 1.375931e-06, 1.375931e-06, 
    1.375927e-06, 1.375924e-06, 1.375922e-06, 1.37592e-06, 1.375919e-06, 
    1.375914e-06, 1.375911e-06, 1.375906e-06, 1.375907e-06, 1.375905e-06, 
    1.375903e-06, 1.375901e-06, 1.375901e-06, 1.3759e-06, 1.375905e-06, 
    1.375902e-06, 1.375907e-06, 1.375906e-06, 1.375918e-06, 1.375923e-06, 
    1.375925e-06, 1.375927e-06, 1.375931e-06, 1.375928e-06, 1.375929e-06, 
    1.375926e-06, 1.375925e-06, 1.375926e-06, 1.37592e-06, 1.375922e-06, 
    1.375911e-06, 1.375916e-06, 1.375904e-06, 1.375907e-06, 1.375903e-06, 
    1.375905e-06, 1.375902e-06, 1.375905e-06, 1.3759e-06, 1.375898e-06, 
    1.375899e-06, 1.375896e-06, 1.375905e-06, 1.375902e-06, 1.375926e-06, 
    1.375925e-06, 1.375925e-06, 1.375928e-06, 1.375928e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.375922e-06, 
    1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375906e-06, 1.375904e-06, 
    1.375906e-06, 1.375904e-06, 1.375906e-06, 1.375906e-06, 1.375899e-06, 
    1.375903e-06, 1.375897e-06, 1.375897e-06, 1.3759e-06, 1.375897e-06, 
    1.375925e-06, 1.375926e-06, 1.375929e-06, 1.375927e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375922e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375916e-06, 1.375911e-06, 1.375907e-06, 1.375903e-06, 
    1.375904e-06, 1.375904e-06, 1.375903e-06, 1.375905e-06, 1.375902e-06, 
    1.375902e-06, 1.375903e-06, 1.375897e-06, 1.375899e-06, 1.375897e-06, 
    1.375898e-06, 1.375926e-06, 1.375925e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.37592e-06, 1.375919e-06, 1.375913e-06, 1.375916e-06, 
    1.375912e-06, 1.375915e-06, 1.375915e-06, 1.375911e-06, 1.375915e-06, 
    1.375907e-06, 1.375912e-06, 1.375903e-06, 1.375908e-06, 1.375902e-06, 
    1.375903e-06, 1.375902e-06, 1.3759e-06, 1.375898e-06, 1.375895e-06, 
    1.375896e-06, 1.375893e-06, 1.375922e-06, 1.375921e-06, 1.375921e-06, 
    1.375919e-06, 1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375912e-06, 
    1.375908e-06, 1.375908e-06, 1.375913e-06, 1.37591e-06, 1.37592e-06, 
    1.375918e-06, 1.375919e-06, 1.375922e-06, 1.375911e-06, 1.375917e-06, 
    1.375906e-06, 1.37591e-06, 1.375901e-06, 1.375905e-06, 1.375896e-06, 
    1.375892e-06, 1.375889e-06, 1.375885e-06, 1.37592e-06, 1.375921e-06, 
    1.375919e-06, 1.375916e-06, 1.375913e-06, 1.375909e-06, 1.375909e-06, 
    1.375908e-06, 1.375906e-06, 1.375905e-06, 1.375908e-06, 1.375905e-06, 
    1.375917e-06, 1.375911e-06, 1.375921e-06, 1.375918e-06, 1.375916e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375893e-06, 1.3759e-06, 1.375882e-06, 1.375887e-06, 1.375921e-06, 
    1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 1.375907e-06, 
    1.375906e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375904e-06, 
    1.375902e-06, 1.375909e-06, 1.375906e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375915e-06, 1.375911e-06, 1.375908e-06, 1.375908e-06, 
    1.375907e-06, 1.375904e-06, 1.375909e-06, 1.375893e-06, 1.375903e-06, 
    1.375918e-06, 1.375915e-06, 1.375914e-06, 1.375916e-06, 1.375907e-06, 
    1.37591e-06, 1.375902e-06, 1.375905e-06, 1.375901e-06, 1.375903e-06, 
    1.375903e-06, 1.375905e-06, 1.375907e-06, 1.37591e-06, 1.375913e-06, 
    1.375915e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375903e-06, 
    1.375904e-06, 1.375901e-06, 1.37591e-06, 1.375906e-06, 1.375907e-06, 
    1.375904e-06, 1.375912e-06, 1.375905e-06, 1.375913e-06, 1.375913e-06, 
    1.37591e-06, 1.375906e-06, 1.375905e-06, 1.375904e-06, 1.375904e-06, 
    1.375908e-06, 1.375908e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 
    1.375914e-06, 1.375913e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.3759e-06, 1.375899e-06, 1.375895e-06, 1.375898e-06, 1.375893e-06, 
    1.375898e-06, 1.375889e-06, 1.375905e-06, 1.375898e-06, 1.37591e-06, 
    1.375909e-06, 1.375906e-06, 1.375901e-06, 1.375904e-06, 1.3759e-06, 
    1.375908e-06, 1.375912e-06, 1.375913e-06, 1.375915e-06, 1.375913e-06, 
    1.375913e-06, 1.375911e-06, 1.375912e-06, 1.375907e-06, 1.37591e-06, 
    1.375903e-06, 1.3759e-06, 1.375893e-06, 1.375889e-06, 1.375884e-06, 
    1.375882e-06, 1.375882e-06, 1.375882e-06 ;

 TOTLITN_1m =
  1.37593e-06, 1.375926e-06, 1.375927e-06, 1.375923e-06, 1.375925e-06, 
    1.375923e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 1.37593e-06, 
    1.375917e-06, 1.375923e-06, 1.375911e-06, 1.375915e-06, 1.375905e-06, 
    1.375911e-06, 1.375903e-06, 1.375905e-06, 1.3759e-06, 1.375902e-06, 
    1.375896e-06, 1.3759e-06, 1.375893e-06, 1.375897e-06, 1.375896e-06, 
    1.3759e-06, 1.375922e-06, 1.375918e-06, 1.375922e-06, 1.375922e-06, 
    1.375922e-06, 1.375925e-06, 1.375927e-06, 1.37593e-06, 1.37593e-06, 
    1.375927e-06, 1.375922e-06, 1.375923e-06, 1.375918e-06, 1.375919e-06, 
    1.375913e-06, 1.375916e-06, 1.375906e-06, 1.375909e-06, 1.375901e-06, 
    1.375903e-06, 1.375902e-06, 1.375902e-06, 1.375902e-06, 1.375904e-06, 
    1.375903e-06, 1.375906e-06, 1.375915e-06, 1.375912e-06, 1.375921e-06, 
    1.375926e-06, 1.375929e-06, 1.375932e-06, 1.375931e-06, 1.375931e-06, 
    1.375927e-06, 1.375924e-06, 1.375922e-06, 1.37592e-06, 1.375919e-06, 
    1.375914e-06, 1.375911e-06, 1.375906e-06, 1.375907e-06, 1.375905e-06, 
    1.375903e-06, 1.375901e-06, 1.375901e-06, 1.3759e-06, 1.375905e-06, 
    1.375902e-06, 1.375907e-06, 1.375906e-06, 1.375918e-06, 1.375923e-06, 
    1.375925e-06, 1.375927e-06, 1.375931e-06, 1.375928e-06, 1.375929e-06, 
    1.375926e-06, 1.375925e-06, 1.375926e-06, 1.37592e-06, 1.375922e-06, 
    1.375911e-06, 1.375916e-06, 1.375904e-06, 1.375907e-06, 1.375903e-06, 
    1.375905e-06, 1.375902e-06, 1.375905e-06, 1.3759e-06, 1.375898e-06, 
    1.375899e-06, 1.375896e-06, 1.375905e-06, 1.375902e-06, 1.375926e-06, 
    1.375925e-06, 1.375925e-06, 1.375928e-06, 1.375928e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.375922e-06, 
    1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375906e-06, 1.375904e-06, 
    1.375906e-06, 1.375904e-06, 1.375906e-06, 1.375906e-06, 1.375899e-06, 
    1.375903e-06, 1.375897e-06, 1.375897e-06, 1.3759e-06, 1.375897e-06, 
    1.375925e-06, 1.375926e-06, 1.375929e-06, 1.375927e-06, 1.375931e-06, 
    1.375928e-06, 1.375927e-06, 1.375922e-06, 1.375921e-06, 1.37592e-06, 
    1.375918e-06, 1.375916e-06, 1.375911e-06, 1.375907e-06, 1.375903e-06, 
    1.375904e-06, 1.375904e-06, 1.375903e-06, 1.375905e-06, 1.375902e-06, 
    1.375902e-06, 1.375903e-06, 1.375897e-06, 1.375899e-06, 1.375897e-06, 
    1.375898e-06, 1.375926e-06, 1.375925e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.37592e-06, 1.375919e-06, 1.375913e-06, 1.375916e-06, 
    1.375912e-06, 1.375915e-06, 1.375915e-06, 1.375911e-06, 1.375915e-06, 
    1.375907e-06, 1.375912e-06, 1.375903e-06, 1.375908e-06, 1.375902e-06, 
    1.375903e-06, 1.375902e-06, 1.3759e-06, 1.375898e-06, 1.375895e-06, 
    1.375896e-06, 1.375893e-06, 1.375922e-06, 1.375921e-06, 1.375921e-06, 
    1.375919e-06, 1.375918e-06, 1.375915e-06, 1.37591e-06, 1.375912e-06, 
    1.375908e-06, 1.375908e-06, 1.375913e-06, 1.37591e-06, 1.37592e-06, 
    1.375918e-06, 1.375919e-06, 1.375922e-06, 1.375911e-06, 1.375917e-06, 
    1.375906e-06, 1.37591e-06, 1.375901e-06, 1.375905e-06, 1.375896e-06, 
    1.375892e-06, 1.375889e-06, 1.375885e-06, 1.37592e-06, 1.375921e-06, 
    1.375919e-06, 1.375916e-06, 1.375913e-06, 1.375909e-06, 1.375909e-06, 
    1.375908e-06, 1.375906e-06, 1.375905e-06, 1.375908e-06, 1.375905e-06, 
    1.375917e-06, 1.375911e-06, 1.375921e-06, 1.375918e-06, 1.375916e-06, 
    1.375917e-06, 1.375912e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375893e-06, 1.3759e-06, 1.375882e-06, 1.375887e-06, 1.375921e-06, 
    1.37592e-06, 1.375914e-06, 1.375917e-06, 1.375909e-06, 1.375907e-06, 
    1.375906e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375904e-06, 
    1.375902e-06, 1.375909e-06, 1.375906e-06, 1.375915e-06, 1.375913e-06, 
    1.375914e-06, 1.375915e-06, 1.375911e-06, 1.375908e-06, 1.375908e-06, 
    1.375907e-06, 1.375904e-06, 1.375909e-06, 1.375893e-06, 1.375903e-06, 
    1.375918e-06, 1.375915e-06, 1.375914e-06, 1.375916e-06, 1.375907e-06, 
    1.37591e-06, 1.375902e-06, 1.375905e-06, 1.375901e-06, 1.375903e-06, 
    1.375903e-06, 1.375905e-06, 1.375907e-06, 1.37591e-06, 1.375913e-06, 
    1.375915e-06, 1.375915e-06, 1.375912e-06, 1.375908e-06, 1.375903e-06, 
    1.375904e-06, 1.375901e-06, 1.37591e-06, 1.375906e-06, 1.375907e-06, 
    1.375904e-06, 1.375912e-06, 1.375905e-06, 1.375913e-06, 1.375913e-06, 
    1.37591e-06, 1.375906e-06, 1.375905e-06, 1.375904e-06, 1.375904e-06, 
    1.375908e-06, 1.375908e-06, 1.37591e-06, 1.375911e-06, 1.375913e-06, 
    1.375914e-06, 1.375913e-06, 1.375912e-06, 1.375908e-06, 1.375904e-06, 
    1.3759e-06, 1.375899e-06, 1.375895e-06, 1.375898e-06, 1.375893e-06, 
    1.375898e-06, 1.375889e-06, 1.375905e-06, 1.375898e-06, 1.37591e-06, 
    1.375909e-06, 1.375906e-06, 1.375901e-06, 1.375904e-06, 1.3759e-06, 
    1.375908e-06, 1.375912e-06, 1.375913e-06, 1.375915e-06, 1.375913e-06, 
    1.375913e-06, 1.375911e-06, 1.375912e-06, 1.375907e-06, 1.37591e-06, 
    1.375903e-06, 1.3759e-06, 1.375893e-06, 1.375889e-06, 1.375884e-06, 
    1.375882e-06, 1.375882e-06, 1.375882e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34458, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34452, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34454, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773745, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773748, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773737, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773745, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773748, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773737, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  243.0869, 243.0901, 243.0895, 243.0921, 243.0906, 243.0923, 243.0875, 
    243.0902, 243.0885, 243.0872, 243.097, 243.0922, 243.1021, 243.0991, 
    243.1068, 243.1016, 243.1079, 243.1067, 243.1103, 243.1093, 243.1137, 
    243.1108, 243.1161, 243.1131, 243.1135, 243.1107, 243.0932, 243.0963, 
    243.093, 243.0934, 243.0932, 243.0907, 243.0893, 243.0866, 243.0871, 
    243.0891, 243.0936, 243.0921, 243.096, 243.0959, 243.1002, 243.0983, 
    243.1055, 243.1034, 243.1093, 243.1078, 243.1092, 243.1088, 243.1092, 
    243.1071, 243.108, 243.1061, 243.0986, 243.1008, 243.0943, 243.0902, 
    243.0876, 243.0858, 243.086, 243.0865, 243.0891, 243.0916, 243.0935, 
    243.0947, 243.0959, 243.0995, 243.1015, 243.1059, 243.1051, 243.1064, 
    243.1077, 243.1098, 243.1095, 243.1104, 243.1064, 243.109, 243.1047, 
    243.1059, 243.0961, 243.0926, 243.0909, 243.0896, 243.0862, 243.0885, 
    243.0876, 243.0898, 243.0912, 243.0905, 243.0947, 243.0931, 243.1016, 
    243.098, 243.1075, 243.1053, 243.1081, 243.1067, 243.1091, 243.1069, 
    243.1107, 243.1115, 243.111, 243.1132, 243.1068, 243.1092, 243.0905, 
    243.0906, 243.0911, 243.0888, 243.0887, 243.0866, 243.0885, 243.0893, 
    243.0913, 243.0925, 243.0936, 243.0961, 243.0988, 243.1026, 243.1054, 
    243.1073, 243.1061, 243.1071, 243.106, 243.1055, 243.1112, 243.108, 
    243.1129, 243.1126, 243.1104, 243.1126, 243.0907, 243.0901, 243.0878, 
    243.0896, 243.0864, 243.0882, 243.0892, 243.0931, 243.094, 243.0948, 
    243.0964, 243.0984, 243.1019, 243.1049, 243.1078, 243.1076, 243.1076, 
    243.1082, 243.1067, 243.1085, 243.1088, 243.108, 243.1126, 243.1113, 
    243.1126, 243.1118, 243.0903, 243.0914, 243.0908, 243.0918, 243.0911, 
    243.0945, 243.0955, 243.1003, 243.0983, 243.1014, 243.0987, 243.0992, 
    243.1014, 243.0988, 243.1048, 243.1007, 243.1083, 243.1041, 243.1085, 
    243.1078, 243.1091, 243.1102, 243.1116, 243.1143, 243.1137, 243.1159, 
    243.093, 243.0943, 243.0942, 243.0957, 243.0967, 243.0991, 243.1028, 
    243.1014, 243.104, 243.1045, 243.1006, 243.103, 243.0953, 243.0965, 
    243.0958, 243.093, 243.1017, 243.0972, 243.1055, 243.1031, 243.11, 
    243.1065, 243.1133, 243.1161, 243.1189, 243.122, 243.0951, 243.0942, 
    243.0959, 243.0981, 243.1003, 243.1032, 243.1035, 243.104, 243.1054, 
    243.1066, 243.1042, 243.1069, 243.0967, 243.1021, 243.0938, 243.0962, 
    243.098, 243.0973, 243.1013, 243.1022, 243.1059, 243.104, 243.1154, 
    243.1104, 243.1244, 243.1205, 243.0938, 243.0951, 243.0995, 243.0974, 
    243.1034, 243.1049, 243.1061, 243.1076, 243.1078, 243.1086, 243.1072, 
    243.1086, 243.1032, 243.1056, 243.099, 243.1006, 243.0999, 243.0991, 
    243.1016, 243.1042, 243.1043, 243.1051, 243.1074, 243.1034, 243.1159, 
    243.1081, 243.0965, 243.0989, 243.0993, 243.0983, 243.1047, 243.1024, 
    243.1086, 243.107, 243.1097, 243.1083, 243.1081, 243.1064, 243.1053, 
    243.1025, 243.1003, 243.0985, 243.0989, 243.1008, 243.1044, 243.1077, 
    243.107, 243.1095, 243.103, 243.1057, 243.1046, 243.1074, 243.1013, 
    243.1063, 243.1001, 243.1006, 243.1024, 243.1058, 243.1067, 243.1075, 
    243.107, 243.1045, 243.1041, 243.1023, 243.1018, 243.1005, 243.0994, 
    243.1004, 243.1014, 243.1045, 243.1072, 243.1102, 243.1109, 243.1143, 
    243.1115, 243.116, 243.112, 243.1189, 243.1067, 243.112, 243.1025, 
    243.1035, 243.1053, 243.1097, 243.1074, 243.1101, 243.1041, 243.1009, 
    243.1001, 243.0986, 243.1002, 243.1, 243.1015, 243.101, 243.1046, 
    243.1027, 243.1081, 243.1101, 243.1156, 243.119, 243.1225, 243.124, 
    243.1245, 243.1246 ;

 TREFMNAV_R =
  243.0869, 243.0901, 243.0895, 243.0921, 243.0906, 243.0923, 243.0875, 
    243.0902, 243.0885, 243.0872, 243.097, 243.0922, 243.1021, 243.0991, 
    243.1068, 243.1016, 243.1079, 243.1067, 243.1103, 243.1093, 243.1137, 
    243.1108, 243.1161, 243.1131, 243.1135, 243.1107, 243.0932, 243.0963, 
    243.093, 243.0934, 243.0932, 243.0907, 243.0893, 243.0866, 243.0871, 
    243.0891, 243.0936, 243.0921, 243.096, 243.0959, 243.1002, 243.0983, 
    243.1055, 243.1034, 243.1093, 243.1078, 243.1092, 243.1088, 243.1092, 
    243.1071, 243.108, 243.1061, 243.0986, 243.1008, 243.0943, 243.0902, 
    243.0876, 243.0858, 243.086, 243.0865, 243.0891, 243.0916, 243.0935, 
    243.0947, 243.0959, 243.0995, 243.1015, 243.1059, 243.1051, 243.1064, 
    243.1077, 243.1098, 243.1095, 243.1104, 243.1064, 243.109, 243.1047, 
    243.1059, 243.0961, 243.0926, 243.0909, 243.0896, 243.0862, 243.0885, 
    243.0876, 243.0898, 243.0912, 243.0905, 243.0947, 243.0931, 243.1016, 
    243.098, 243.1075, 243.1053, 243.1081, 243.1067, 243.1091, 243.1069, 
    243.1107, 243.1115, 243.111, 243.1132, 243.1068, 243.1092, 243.0905, 
    243.0906, 243.0911, 243.0888, 243.0887, 243.0866, 243.0885, 243.0893, 
    243.0913, 243.0925, 243.0936, 243.0961, 243.0988, 243.1026, 243.1054, 
    243.1073, 243.1061, 243.1071, 243.106, 243.1055, 243.1112, 243.108, 
    243.1129, 243.1126, 243.1104, 243.1126, 243.0907, 243.0901, 243.0878, 
    243.0896, 243.0864, 243.0882, 243.0892, 243.0931, 243.094, 243.0948, 
    243.0964, 243.0984, 243.1019, 243.1049, 243.1078, 243.1076, 243.1076, 
    243.1082, 243.1067, 243.1085, 243.1088, 243.108, 243.1126, 243.1113, 
    243.1126, 243.1118, 243.0903, 243.0914, 243.0908, 243.0918, 243.0911, 
    243.0945, 243.0955, 243.1003, 243.0983, 243.1014, 243.0987, 243.0992, 
    243.1014, 243.0988, 243.1048, 243.1007, 243.1083, 243.1041, 243.1085, 
    243.1078, 243.1091, 243.1102, 243.1116, 243.1143, 243.1137, 243.1159, 
    243.093, 243.0943, 243.0942, 243.0957, 243.0967, 243.0991, 243.1028, 
    243.1014, 243.104, 243.1045, 243.1006, 243.103, 243.0953, 243.0965, 
    243.0958, 243.093, 243.1017, 243.0972, 243.1055, 243.1031, 243.11, 
    243.1065, 243.1133, 243.1161, 243.1189, 243.122, 243.0951, 243.0942, 
    243.0959, 243.0981, 243.1003, 243.1032, 243.1035, 243.104, 243.1054, 
    243.1066, 243.1042, 243.1069, 243.0967, 243.1021, 243.0938, 243.0962, 
    243.098, 243.0973, 243.1013, 243.1022, 243.1059, 243.104, 243.1154, 
    243.1104, 243.1244, 243.1205, 243.0938, 243.0951, 243.0995, 243.0974, 
    243.1034, 243.1049, 243.1061, 243.1076, 243.1078, 243.1086, 243.1072, 
    243.1086, 243.1032, 243.1056, 243.099, 243.1006, 243.0999, 243.0991, 
    243.1016, 243.1042, 243.1043, 243.1051, 243.1074, 243.1034, 243.1159, 
    243.1081, 243.0965, 243.0989, 243.0993, 243.0983, 243.1047, 243.1024, 
    243.1086, 243.107, 243.1097, 243.1083, 243.1081, 243.1064, 243.1053, 
    243.1025, 243.1003, 243.0985, 243.0989, 243.1008, 243.1044, 243.1077, 
    243.107, 243.1095, 243.103, 243.1057, 243.1046, 243.1074, 243.1013, 
    243.1063, 243.1001, 243.1006, 243.1024, 243.1058, 243.1067, 243.1075, 
    243.107, 243.1045, 243.1041, 243.1023, 243.1018, 243.1005, 243.0994, 
    243.1004, 243.1014, 243.1045, 243.1072, 243.1102, 243.1109, 243.1143, 
    243.1115, 243.116, 243.112, 243.1189, 243.1067, 243.112, 243.1025, 
    243.1035, 243.1053, 243.1097, 243.1074, 243.1101, 243.1041, 243.1009, 
    243.1001, 243.0986, 243.1002, 243.1, 243.1015, 243.101, 243.1046, 
    243.1027, 243.1081, 243.1101, 243.1156, 243.119, 243.1225, 243.124, 
    243.1245, 243.1246 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7644, 270.7623, 270.7627, 270.761, 270.7619, 270.7608, 270.7639, 
    270.7622, 270.7633, 270.7642, 270.7578, 270.7609, 270.7544, 270.7564, 
    270.7513, 270.7547, 270.7506, 270.7513, 270.749, 270.7496, 270.7467, 
    270.7486, 270.7451, 270.7471, 270.7468, 270.7487, 270.7603, 270.7582, 
    270.7604, 270.7601, 270.7602, 270.7619, 270.7628, 270.7645, 270.7642, 
    270.7629, 270.7599, 270.7609, 270.7584, 270.7585, 270.7556, 270.7569, 
    270.7522, 270.7535, 270.7496, 270.7506, 270.7497, 270.7499, 270.7497, 
    270.7511, 270.7505, 270.7517, 270.7567, 270.7552, 270.7596, 270.7622, 
    270.7639, 270.7651, 270.7649, 270.7646, 270.7629, 270.7613, 270.7601, 
    270.7593, 270.7585, 270.7561, 270.7548, 270.7519, 270.7524, 270.7516, 
    270.7507, 270.7493, 270.7495, 270.7489, 270.7516, 270.7498, 270.7527, 
    270.7519, 270.7584, 270.7607, 270.7617, 270.7626, 270.7648, 270.7633, 
    270.7639, 270.7625, 270.7616, 270.762, 270.7592, 270.7603, 270.7547, 
    270.7571, 270.7508, 270.7523, 270.7504, 270.7514, 270.7498, 270.7512, 
    270.7487, 270.7481, 270.7485, 270.747, 270.7513, 270.7497, 270.762, 
    270.7619, 270.7616, 270.7631, 270.7632, 270.7646, 270.7633, 270.7628, 
    270.7615, 270.7607, 270.76, 270.7584, 270.7566, 270.7541, 270.7522, 
    270.751, 270.7517, 270.7511, 270.7518, 270.7521, 270.7483, 270.7505, 
    270.7472, 270.7474, 270.7489, 270.7474, 270.7619, 270.7623, 270.7638, 
    270.7626, 270.7647, 270.7635, 270.7629, 270.7603, 270.7597, 270.7592, 
    270.7582, 270.7568, 270.7545, 270.7525, 270.7506, 270.7508, 270.7507, 
    270.7503, 270.7513, 270.7502, 270.75, 270.7505, 270.7474, 270.7483, 
    270.7474, 270.748, 270.7621, 270.7615, 270.7618, 270.7611, 270.7617, 
    270.7594, 270.7588, 270.7556, 270.7569, 270.7549, 270.7567, 270.7563, 
    270.7548, 270.7566, 270.7527, 270.7553, 270.7503, 270.7531, 270.7501, 
    270.7506, 270.7498, 270.749, 270.748, 270.7463, 270.7467, 270.7452, 
    270.7604, 270.7595, 270.7596, 270.7586, 270.7579, 270.7564, 270.7539, 
    270.7549, 270.7531, 270.7528, 270.7554, 270.7538, 270.7589, 270.7581, 
    270.7586, 270.7603, 270.7547, 270.7576, 270.7522, 270.7538, 270.7491, 
    270.7515, 270.7469, 270.7451, 270.7432, 270.7411, 270.759, 270.7596, 
    270.7585, 270.757, 270.7556, 270.7537, 270.7534, 270.7531, 270.7522, 
    270.7514, 270.753, 270.7512, 270.758, 270.7544, 270.7599, 270.7583, 
    270.7571, 270.7576, 270.7549, 270.7543, 270.7519, 270.7531, 270.7455, 
    270.7489, 270.7395, 270.7421, 270.7598, 270.759, 270.7561, 270.7575, 
    270.7535, 270.7526, 270.7518, 270.7508, 270.7506, 270.7501, 270.751, 
    270.7501, 270.7537, 270.7521, 270.7564, 270.7554, 270.7559, 270.7564, 
    270.7547, 270.753, 270.7529, 270.7524, 270.7509, 270.7535, 270.7452, 
    270.7504, 270.7581, 270.7565, 270.7563, 270.7569, 270.7527, 270.7542, 
    270.7501, 270.7512, 270.7494, 270.7502, 270.7504, 270.7516, 270.7523, 
    270.7541, 270.7556, 270.7568, 270.7565, 270.7552, 270.7529, 270.7506, 
    270.7512, 270.7495, 270.7538, 270.752, 270.7527, 270.7509, 270.7549, 
    270.7516, 270.7557, 270.7554, 270.7542, 270.7519, 270.7513, 270.7508, 
    270.7512, 270.7528, 270.7531, 270.7542, 270.7546, 270.7555, 270.7562, 
    270.7555, 270.7548, 270.7528, 270.751, 270.749, 270.7485, 270.7463, 
    270.7482, 270.7452, 270.7478, 270.7432, 270.7513, 270.7478, 270.7542, 
    270.7534, 270.7523, 270.7494, 270.7509, 270.7491, 270.7531, 270.7552, 
    270.7557, 270.7567, 270.7557, 270.7558, 270.7548, 270.7551, 270.7527, 
    270.754, 270.7504, 270.7491, 270.7454, 270.7431, 270.7408, 270.7397, 
    270.7394, 270.7393 ;

 TREFMXAV_R =
  270.7644, 270.7623, 270.7627, 270.761, 270.7619, 270.7608, 270.7639, 
    270.7622, 270.7633, 270.7642, 270.7578, 270.7609, 270.7544, 270.7564, 
    270.7513, 270.7547, 270.7506, 270.7513, 270.749, 270.7496, 270.7467, 
    270.7486, 270.7451, 270.7471, 270.7468, 270.7487, 270.7603, 270.7582, 
    270.7604, 270.7601, 270.7602, 270.7619, 270.7628, 270.7645, 270.7642, 
    270.7629, 270.7599, 270.7609, 270.7584, 270.7585, 270.7556, 270.7569, 
    270.7522, 270.7535, 270.7496, 270.7506, 270.7497, 270.7499, 270.7497, 
    270.7511, 270.7505, 270.7517, 270.7567, 270.7552, 270.7596, 270.7622, 
    270.7639, 270.7651, 270.7649, 270.7646, 270.7629, 270.7613, 270.7601, 
    270.7593, 270.7585, 270.7561, 270.7548, 270.7519, 270.7524, 270.7516, 
    270.7507, 270.7493, 270.7495, 270.7489, 270.7516, 270.7498, 270.7527, 
    270.7519, 270.7584, 270.7607, 270.7617, 270.7626, 270.7648, 270.7633, 
    270.7639, 270.7625, 270.7616, 270.762, 270.7592, 270.7603, 270.7547, 
    270.7571, 270.7508, 270.7523, 270.7504, 270.7514, 270.7498, 270.7512, 
    270.7487, 270.7481, 270.7485, 270.747, 270.7513, 270.7497, 270.762, 
    270.7619, 270.7616, 270.7631, 270.7632, 270.7646, 270.7633, 270.7628, 
    270.7615, 270.7607, 270.76, 270.7584, 270.7566, 270.7541, 270.7522, 
    270.751, 270.7517, 270.7511, 270.7518, 270.7521, 270.7483, 270.7505, 
    270.7472, 270.7474, 270.7489, 270.7474, 270.7619, 270.7623, 270.7638, 
    270.7626, 270.7647, 270.7635, 270.7629, 270.7603, 270.7597, 270.7592, 
    270.7582, 270.7568, 270.7545, 270.7525, 270.7506, 270.7508, 270.7507, 
    270.7503, 270.7513, 270.7502, 270.75, 270.7505, 270.7474, 270.7483, 
    270.7474, 270.748, 270.7621, 270.7615, 270.7618, 270.7611, 270.7617, 
    270.7594, 270.7588, 270.7556, 270.7569, 270.7549, 270.7567, 270.7563, 
    270.7548, 270.7566, 270.7527, 270.7553, 270.7503, 270.7531, 270.7501, 
    270.7506, 270.7498, 270.749, 270.748, 270.7463, 270.7467, 270.7452, 
    270.7604, 270.7595, 270.7596, 270.7586, 270.7579, 270.7564, 270.7539, 
    270.7549, 270.7531, 270.7528, 270.7554, 270.7538, 270.7589, 270.7581, 
    270.7586, 270.7603, 270.7547, 270.7576, 270.7522, 270.7538, 270.7491, 
    270.7515, 270.7469, 270.7451, 270.7432, 270.7411, 270.759, 270.7596, 
    270.7585, 270.757, 270.7556, 270.7537, 270.7534, 270.7531, 270.7522, 
    270.7514, 270.753, 270.7512, 270.758, 270.7544, 270.7599, 270.7583, 
    270.7571, 270.7576, 270.7549, 270.7543, 270.7519, 270.7531, 270.7455, 
    270.7489, 270.7395, 270.7421, 270.7598, 270.759, 270.7561, 270.7575, 
    270.7535, 270.7526, 270.7518, 270.7508, 270.7506, 270.7501, 270.751, 
    270.7501, 270.7537, 270.7521, 270.7564, 270.7554, 270.7559, 270.7564, 
    270.7547, 270.753, 270.7529, 270.7524, 270.7509, 270.7535, 270.7452, 
    270.7504, 270.7581, 270.7565, 270.7563, 270.7569, 270.7527, 270.7542, 
    270.7501, 270.7512, 270.7494, 270.7502, 270.7504, 270.7516, 270.7523, 
    270.7541, 270.7556, 270.7568, 270.7565, 270.7552, 270.7529, 270.7506, 
    270.7512, 270.7495, 270.7538, 270.752, 270.7527, 270.7509, 270.7549, 
    270.7516, 270.7557, 270.7554, 270.7542, 270.7519, 270.7513, 270.7508, 
    270.7512, 270.7528, 270.7531, 270.7542, 270.7546, 270.7555, 270.7562, 
    270.7555, 270.7548, 270.7528, 270.751, 270.749, 270.7485, 270.7463, 
    270.7482, 270.7452, 270.7478, 270.7432, 270.7513, 270.7478, 270.7542, 
    270.7534, 270.7523, 270.7494, 270.7509, 270.7491, 270.7531, 270.7552, 
    270.7557, 270.7567, 270.7557, 270.7558, 270.7548, 270.7551, 270.7527, 
    270.754, 270.7504, 270.7491, 270.7454, 270.7431, 270.7408, 270.7397, 
    270.7394, 270.7393 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.2032, 255.203, 255.203, 255.2029, 255.203, 255.2029, 255.2031, 255.203, 
    255.2031, 255.2031, 255.2027, 255.2029, 255.2024, 255.2026, 255.2022, 
    255.2025, 255.2021, 255.2022, 255.202, 255.2021, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2019, 255.202, 255.2029, 255.2027, 255.2029, 
    255.2028, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.203, 
    255.2028, 255.2029, 255.2027, 255.2027, 255.2025, 255.2026, 255.2023, 
    255.2024, 255.2021, 255.2021, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2021, 255.2022, 255.2026, 255.2025, 255.2028, 255.203, 255.2031, 
    255.2032, 255.2032, 255.2032, 255.203, 255.2029, 255.2028, 255.2028, 
    255.2027, 255.2026, 255.2025, 255.2022, 255.2023, 255.2022, 255.2021, 
    255.202, 255.2021, 255.202, 255.2022, 255.2021, 255.2023, 255.2022, 
    255.2027, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.2031, 
    255.203, 255.2029, 255.203, 255.2028, 255.2029, 255.2025, 255.2026, 
    255.2021, 255.2023, 255.2021, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.203, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2022, 255.2022, 255.2022, 255.2023, 255.202, 255.2021, 255.2019, 
    255.2019, 255.202, 255.2019, 255.203, 255.203, 255.2031, 255.203, 
    255.2032, 255.2031, 255.203, 255.2029, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 
    255.2022, 255.2021, 255.2021, 255.2021, 255.2019, 255.202, 255.2019, 
    255.2019, 255.203, 255.2029, 255.203, 255.2029, 255.203, 255.2028, 
    255.2027, 255.2025, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 
    255.2026, 255.2023, 255.2025, 255.2021, 255.2023, 255.2021, 255.2021, 
    255.2021, 255.202, 255.202, 255.2018, 255.2018, 255.2017, 255.2029, 
    255.2028, 255.2028, 255.2027, 255.2027, 255.2026, 255.2024, 255.2025, 
    255.2023, 255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2027, 
    255.2029, 255.2024, 255.2027, 255.2023, 255.2024, 255.202, 255.2022, 
    255.2019, 255.2017, 255.2016, 255.2014, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2025, 255.2024, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2027, 255.2024, 255.2028, 255.2027, 255.2026, 
    255.2027, 255.2025, 255.2024, 255.2022, 255.2023, 255.2018, 255.202, 
    255.2013, 255.2015, 255.2028, 255.2028, 255.2025, 255.2027, 255.2024, 
    255.2023, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2026, 255.2025, 255.2025, 255.2026, 255.2025, 
    255.2023, 255.2023, 255.2023, 255.2022, 255.2024, 255.2017, 255.2021, 
    255.2027, 255.2026, 255.2026, 255.2026, 255.2023, 255.2024, 255.2021, 
    255.2022, 255.202, 255.2021, 255.2021, 255.2022, 255.2023, 255.2024, 
    255.2025, 255.2026, 255.2026, 255.2025, 255.2023, 255.2021, 255.2022, 
    255.2021, 255.2024, 255.2022, 255.2023, 255.2022, 255.2025, 255.2022, 
    255.2025, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 255.2022, 
    255.2023, 255.2023, 255.2024, 255.2024, 255.2025, 255.2026, 255.2025, 
    255.2025, 255.2023, 255.2022, 255.202, 255.202, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2016, 255.2022, 255.2019, 255.2024, 255.2023, 
    255.2023, 255.202, 255.2022, 255.202, 255.2023, 255.2025, 255.2025, 
    255.2026, 255.2025, 255.2025, 255.2025, 255.2025, 255.2023, 255.2024, 
    255.2021, 255.202, 255.2018, 255.2016, 255.2014, 255.2013, 255.2013, 
    255.2013 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  255.2032, 255.203, 255.203, 255.2029, 255.203, 255.2029, 255.2031, 255.203, 
    255.2031, 255.2031, 255.2027, 255.2029, 255.2024, 255.2026, 255.2022, 
    255.2025, 255.2021, 255.2022, 255.202, 255.2021, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2019, 255.202, 255.2029, 255.2027, 255.2029, 
    255.2028, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.203, 
    255.2028, 255.2029, 255.2027, 255.2027, 255.2025, 255.2026, 255.2023, 
    255.2024, 255.2021, 255.2021, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2021, 255.2022, 255.2026, 255.2025, 255.2028, 255.203, 255.2031, 
    255.2032, 255.2032, 255.2032, 255.203, 255.2029, 255.2028, 255.2028, 
    255.2027, 255.2026, 255.2025, 255.2022, 255.2023, 255.2022, 255.2021, 
    255.202, 255.2021, 255.202, 255.2022, 255.2021, 255.2023, 255.2022, 
    255.2027, 255.2029, 255.203, 255.203, 255.2032, 255.2031, 255.2031, 
    255.203, 255.2029, 255.203, 255.2028, 255.2029, 255.2025, 255.2026, 
    255.2021, 255.2023, 255.2021, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.203, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2022, 255.2022, 255.2022, 255.2023, 255.202, 255.2021, 255.2019, 
    255.2019, 255.202, 255.2019, 255.203, 255.203, 255.2031, 255.203, 
    255.2032, 255.2031, 255.203, 255.2029, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2023, 255.2021, 255.2021, 255.2021, 255.2021, 
    255.2022, 255.2021, 255.2021, 255.2021, 255.2019, 255.202, 255.2019, 
    255.2019, 255.203, 255.2029, 255.203, 255.2029, 255.203, 255.2028, 
    255.2027, 255.2025, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 
    255.2026, 255.2023, 255.2025, 255.2021, 255.2023, 255.2021, 255.2021, 
    255.2021, 255.202, 255.202, 255.2018, 255.2018, 255.2017, 255.2029, 
    255.2028, 255.2028, 255.2027, 255.2027, 255.2026, 255.2024, 255.2025, 
    255.2023, 255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2027, 
    255.2029, 255.2024, 255.2027, 255.2023, 255.2024, 255.202, 255.2022, 
    255.2019, 255.2017, 255.2016, 255.2014, 255.2028, 255.2028, 255.2027, 
    255.2026, 255.2025, 255.2024, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2027, 255.2024, 255.2028, 255.2027, 255.2026, 
    255.2027, 255.2025, 255.2024, 255.2022, 255.2023, 255.2018, 255.202, 
    255.2013, 255.2015, 255.2028, 255.2028, 255.2025, 255.2027, 255.2024, 
    255.2023, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2026, 255.2025, 255.2025, 255.2026, 255.2025, 
    255.2023, 255.2023, 255.2023, 255.2022, 255.2024, 255.2017, 255.2021, 
    255.2027, 255.2026, 255.2026, 255.2026, 255.2023, 255.2024, 255.2021, 
    255.2022, 255.202, 255.2021, 255.2021, 255.2022, 255.2023, 255.2024, 
    255.2025, 255.2026, 255.2026, 255.2025, 255.2023, 255.2021, 255.2022, 
    255.2021, 255.2024, 255.2022, 255.2023, 255.2022, 255.2025, 255.2022, 
    255.2025, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 255.2022, 
    255.2023, 255.2023, 255.2024, 255.2024, 255.2025, 255.2026, 255.2025, 
    255.2025, 255.2023, 255.2022, 255.202, 255.202, 255.2018, 255.202, 
    255.2017, 255.2019, 255.2016, 255.2022, 255.2019, 255.2024, 255.2023, 
    255.2023, 255.202, 255.2022, 255.202, 255.2023, 255.2025, 255.2025, 
    255.2026, 255.2025, 255.2025, 255.2025, 255.2025, 255.2023, 255.2024, 
    255.2021, 255.202, 255.2018, 255.2016, 255.2014, 255.2013, 255.2013, 
    255.2013 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6895, 253.6914, 253.6911, 253.6926, 253.6917, 253.6927, 253.6899, 
    253.6915, 253.6905, 253.6897, 253.6955, 253.6926, 253.6985, 253.6967, 
    253.7013, 253.6982, 253.702, 253.7013, 253.7034, 253.7028, 253.7055, 
    253.7037, 253.707, 253.7051, 253.7054, 253.7037, 253.6933, 253.6951, 
    253.6931, 253.6934, 253.6933, 253.6918, 253.6909, 253.6894, 253.6897, 
    253.6908, 253.6935, 253.6926, 253.6949, 253.6949, 253.6974, 253.6963, 
    253.7005, 253.6993, 253.7029, 253.702, 253.7028, 253.7026, 253.7028, 
    253.7015, 253.7021, 253.7009, 253.6965, 253.6978, 253.6939, 253.6915, 
    253.69, 253.6889, 253.689, 253.6893, 253.6908, 253.6923, 253.6934, 
    253.6942, 253.6949, 253.697, 253.6982, 253.7008, 253.7003, 253.7011, 
    253.7019, 253.7031, 253.7029, 253.7035, 253.7011, 253.7027, 253.7001, 
    253.7008, 253.6949, 253.6929, 253.6919, 253.6911, 253.6891, 253.6905, 
    253.69, 253.6913, 253.6921, 253.6917, 253.6942, 253.6932, 253.6982, 
    253.6961, 253.7018, 253.7004, 253.7021, 253.7013, 253.7027, 253.7014, 
    253.7037, 253.7042, 253.7039, 253.7052, 253.7013, 253.7028, 253.6917, 
    253.6917, 253.692, 253.6907, 253.6906, 253.6894, 253.6905, 253.6909, 
    253.6921, 253.6928, 253.6935, 253.695, 253.6966, 253.6989, 253.7005, 
    253.7016, 253.7009, 253.7015, 253.7009, 253.7006, 253.704, 253.7021, 
    253.705, 253.7048, 253.7035, 253.7049, 253.6918, 253.6914, 253.6901, 
    253.6911, 253.6892, 253.6903, 253.6909, 253.6932, 253.6937, 253.6942, 
    253.6951, 253.6963, 253.6984, 253.7002, 253.7019, 253.7018, 253.7018, 
    253.7022, 253.7013, 253.7024, 253.7025, 253.7021, 253.7048, 253.704, 
    253.7048, 253.7043, 253.6915, 253.6922, 253.6918, 253.6925, 253.692, 
    253.694, 253.6946, 253.6974, 253.6963, 253.6981, 253.6965, 253.6968, 
    253.6981, 253.6966, 253.7001, 253.6977, 253.7022, 253.6998, 253.7024, 
    253.7019, 253.7027, 253.7034, 253.7043, 253.7058, 253.7055, 253.7068, 
    253.6931, 253.6939, 253.6939, 253.6947, 253.6954, 253.6967, 253.6989, 
    253.6981, 253.6997, 253.7, 253.6976, 253.699, 253.6945, 253.6952, 
    253.6948, 253.6932, 253.6983, 253.6956, 253.7005, 253.6991, 253.7033, 
    253.7012, 253.7053, 253.707, 253.7087, 253.7105, 253.6944, 253.6938, 
    253.6948, 253.6962, 253.6975, 253.6992, 253.6994, 253.6997, 253.7005, 
    253.7012, 253.6998, 253.7014, 253.6953, 253.6985, 253.6936, 253.6951, 
    253.6961, 253.6957, 253.698, 253.6986, 253.7008, 253.6997, 253.7065, 
    253.7035, 253.712, 253.7096, 253.6936, 253.6944, 253.697, 253.6958, 
    253.6993, 253.7002, 253.7009, 253.7018, 253.7019, 253.7025, 253.7016, 
    253.7024, 253.6992, 253.7006, 253.6967, 253.6976, 253.6972, 253.6967, 
    253.6982, 253.6998, 253.6999, 253.7003, 253.7017, 253.6993, 253.7068, 
    253.7021, 253.6952, 253.6966, 253.6969, 253.6963, 253.7001, 253.6987, 
    253.7024, 253.7014, 253.7031, 253.7023, 253.7021, 253.7011, 253.7004, 
    253.6988, 253.6974, 253.6964, 253.6966, 253.6978, 253.6999, 253.7019, 
    253.7015, 253.703, 253.6991, 253.7007, 253.7, 253.7017, 253.6981, 
    253.701, 253.6973, 253.6977, 253.6987, 253.7008, 253.7013, 253.7018, 
    253.7015, 253.7, 253.6997, 253.6987, 253.6984, 253.6976, 253.6969, 
    253.6975, 253.6981, 253.7, 253.7016, 253.7034, 253.7038, 253.7058, 
    253.7041, 253.7069, 253.7045, 253.7087, 253.7013, 253.7045, 253.6988, 
    253.6994, 253.7005, 253.7031, 253.7017, 253.7033, 253.6997, 253.6978, 
    253.6974, 253.6964, 253.6974, 253.6973, 253.6982, 253.6979, 253.7, 
    253.6989, 253.7021, 253.7033, 253.7067, 253.7087, 253.7109, 253.7118, 
    253.7121, 253.7122,
  255.2211, 255.2229, 255.2226, 255.224, 255.2232, 255.2241, 255.2215, 
    255.223, 255.222, 255.2213, 255.2267, 255.224, 255.2295, 255.2278, 
    255.2322, 255.2293, 255.2328, 255.2321, 255.2341, 255.2336, 255.2361, 
    255.2344, 255.2374, 255.2357, 255.2359, 255.2343, 255.2246, 255.2263, 
    255.2245, 255.2247, 255.2246, 255.2232, 255.2225, 255.221, 255.2213, 
    255.2224, 255.2249, 255.224, 255.2262, 255.2261, 255.2285, 255.2274, 
    255.2314, 255.2303, 255.2336, 255.2327, 255.2335, 255.2333, 255.2335, 
    255.2323, 255.2328, 255.2318, 255.2276, 255.2288, 255.2252, 255.223, 
    255.2216, 255.2206, 255.2207, 255.221, 255.2224, 255.2237, 255.2248, 
    255.2254, 255.2261, 255.2281, 255.2292, 255.2316, 255.2312, 255.2319, 
    255.2327, 255.2338, 255.2337, 255.2342, 255.2319, 255.2334, 255.231, 
    255.2316, 255.2262, 255.2243, 255.2234, 255.2226, 255.2208, 255.2221, 
    255.2216, 255.2228, 255.2235, 255.2232, 255.2255, 255.2246, 255.2292, 
    255.2272, 255.2326, 255.2313, 255.2329, 255.2321, 255.2334, 255.2322, 
    255.2344, 255.2348, 255.2345, 255.2358, 255.2321, 255.2335, 255.2231, 
    255.2232, 255.2235, 255.2222, 255.2222, 255.221, 255.222, 255.2225, 
    255.2236, 255.2242, 255.2248, 255.2262, 255.2277, 255.2298, 255.2314, 
    255.2324, 255.2318, 255.2323, 255.2317, 255.2314, 255.2346, 255.2328, 
    255.2356, 255.2354, 255.2342, 255.2355, 255.2233, 255.2229, 255.2217, 
    255.2226, 255.2209, 255.2219, 255.2224, 255.2246, 255.2251, 255.2255, 
    255.2264, 255.2275, 255.2294, 255.2311, 255.2327, 255.2326, 255.2326, 
    255.233, 255.2321, 255.2331, 255.2333, 255.2328, 255.2354, 255.2347, 
    255.2354, 255.235, 255.223, 255.2236, 255.2233, 255.2239, 255.2234, 
    255.2253, 255.2259, 255.2285, 255.2274, 255.2292, 255.2276, 255.2279, 
    255.2292, 255.2277, 255.231, 255.2287, 255.233, 255.2307, 255.2331, 
    255.2327, 255.2334, 255.2341, 255.2349, 255.2364, 255.236, 255.2373, 
    255.2245, 255.2252, 255.2252, 255.226, 255.2266, 255.2279, 255.2299, 
    255.2291, 255.2306, 255.2309, 255.2287, 255.23, 255.2257, 255.2264, 
    255.226, 255.2245, 255.2293, 255.2268, 255.2314, 255.2301, 255.234, 
    255.232, 255.2358, 255.2374, 255.239, 255.2408, 255.2257, 255.2251, 
    255.2261, 255.2273, 255.2285, 255.2301, 255.2303, 255.2306, 255.2314, 
    255.232, 255.2307, 255.2322, 255.2265, 255.2295, 255.2249, 255.2263, 
    255.2273, 255.2269, 255.2291, 255.2296, 255.2317, 255.2306, 255.237, 
    255.2342, 255.2422, 255.2399, 255.225, 255.2257, 255.2281, 255.2269, 
    255.2303, 255.2311, 255.2318, 255.2326, 255.2327, 255.2332, 255.2324, 
    255.2332, 255.2301, 255.2315, 255.2278, 255.2287, 255.2283, 255.2279, 
    255.2292, 255.2307, 255.2308, 255.2312, 255.2325, 255.2303, 255.2373, 
    255.2329, 255.2264, 255.2277, 255.228, 255.2274, 255.231, 255.2297, 
    255.2332, 255.2323, 255.2338, 255.233, 255.2329, 255.2319, 255.2313, 
    255.2298, 255.2285, 255.2275, 255.2278, 255.2288, 255.2308, 255.2327, 
    255.2323, 255.2337, 255.23, 255.2315, 255.2309, 255.2325, 255.2291, 
    255.2319, 255.2284, 255.2287, 255.2297, 255.2316, 255.2321, 255.2325, 
    255.2323, 255.2309, 255.2306, 255.2297, 255.2294, 255.2286, 255.228, 
    255.2286, 255.2292, 255.2309, 255.2324, 255.2341, 255.2345, 255.2364, 
    255.2348, 255.2374, 255.2351, 255.239, 255.2321, 255.2351, 255.2297, 
    255.2303, 255.2313, 255.2338, 255.2325, 255.234, 255.2306, 255.2289, 
    255.2284, 255.2276, 255.2285, 255.2284, 255.2292, 255.2289, 255.2309, 
    255.2299, 255.2329, 255.234, 255.2372, 255.2391, 255.2411, 255.242, 
    255.2422, 255.2424,
  257.2871, 257.2885, 257.2882, 257.2894, 257.2888, 257.2895, 257.2874, 
    257.2885, 257.2878, 257.2872, 257.2916, 257.2894, 257.2939, 257.2925, 
    257.296, 257.2936, 257.2965, 257.296, 257.2976, 257.2971, 257.2992, 
    257.2978, 257.3003, 257.2989, 257.2991, 257.2978, 257.2899, 257.2913, 
    257.2898, 257.29, 257.2899, 257.2888, 257.2882, 257.287, 257.2872, 
    257.2881, 257.2901, 257.2894, 257.2911, 257.2911, 257.293, 257.2921, 
    257.2954, 257.2945, 257.2971, 257.2965, 257.2971, 257.2969, 257.2971, 
    257.2961, 257.2965, 257.2957, 257.2923, 257.2933, 257.2903, 257.2886, 
    257.2874, 257.2866, 257.2867, 257.287, 257.2881, 257.2892, 257.29, 
    257.2906, 257.2911, 257.2927, 257.2936, 257.2956, 257.2952, 257.2958, 
    257.2964, 257.2974, 257.2972, 257.2976, 257.2958, 257.297, 257.295, 
    257.2956, 257.2912, 257.2896, 257.2889, 257.2883, 257.2868, 257.2878, 
    257.2874, 257.2884, 257.289, 257.2887, 257.2906, 257.2898, 257.2936, 
    257.292, 257.2963, 257.2953, 257.2966, 257.2959, 257.2971, 257.2961, 
    257.2978, 257.2982, 257.2979, 257.299, 257.296, 257.2971, 257.2887, 
    257.2888, 257.289, 257.288, 257.2879, 257.287, 257.2878, 257.2881, 
    257.289, 257.2896, 257.2901, 257.2912, 257.2924, 257.2941, 257.2953, 
    257.2962, 257.2957, 257.2961, 257.2956, 257.2954, 257.298, 257.2965, 
    257.2988, 257.2987, 257.2976, 257.2987, 257.2888, 257.2885, 257.2875, 
    257.2883, 257.2869, 257.2877, 257.2881, 257.2898, 257.2902, 257.2906, 
    257.2913, 257.2922, 257.2938, 257.2952, 257.2964, 257.2964, 257.2964, 
    257.2967, 257.296, 257.2968, 257.2969, 257.2966, 257.2987, 257.2981, 
    257.2987, 257.2983, 257.2886, 257.2891, 257.2888, 257.2893, 257.2889, 
    257.2904, 257.2909, 257.293, 257.2922, 257.2935, 257.2923, 257.2925, 
    257.2936, 257.2924, 257.2951, 257.2932, 257.2967, 257.2948, 257.2968, 
    257.2964, 257.297, 257.2975, 257.2982, 257.2994, 257.2992, 257.3002, 
    257.2898, 257.2904, 257.2903, 257.291, 257.2914, 257.2925, 257.2942, 
    257.2935, 257.2947, 257.2949, 257.2932, 257.2943, 257.2908, 257.2913, 
    257.291, 257.2898, 257.2937, 257.2917, 257.2954, 257.2943, 257.2975, 
    257.2959, 257.299, 257.3003, 257.3016, 257.3031, 257.2907, 257.2903, 
    257.2911, 257.2921, 257.2931, 257.2944, 257.2945, 257.2947, 257.2954, 
    257.2959, 257.2948, 257.2961, 257.2914, 257.2939, 257.2901, 257.2912, 
    257.292, 257.2917, 257.2935, 257.2939, 257.2956, 257.2947, 257.3, 
    257.2976, 257.3043, 257.3024, 257.2902, 257.2907, 257.2927, 257.2917, 
    257.2945, 257.2951, 257.2957, 257.2964, 257.2964, 257.2968, 257.2962, 
    257.2968, 257.2944, 257.2955, 257.2925, 257.2932, 257.2929, 257.2925, 
    257.2936, 257.2948, 257.2949, 257.2952, 257.2963, 257.2945, 257.3002, 
    257.2966, 257.2914, 257.2924, 257.2926, 257.2922, 257.295, 257.294, 
    257.2968, 257.2961, 257.2973, 257.2967, 257.2966, 257.2958, 257.2953, 
    257.294, 257.293, 257.2922, 257.2924, 257.2933, 257.2949, 257.2964, 
    257.2961, 257.2972, 257.2943, 257.2955, 257.295, 257.2963, 257.2935, 
    257.2958, 257.2929, 257.2932, 257.294, 257.2956, 257.2959, 257.2963, 
    257.2961, 257.295, 257.2948, 257.294, 257.2937, 257.2932, 257.2926, 
    257.2931, 257.2935, 257.295, 257.2962, 257.2975, 257.2979, 257.2994, 
    257.2982, 257.3003, 257.2984, 257.3016, 257.296, 257.2984, 257.294, 
    257.2945, 257.2953, 257.2973, 257.2963, 257.2975, 257.2948, 257.2933, 
    257.293, 257.2923, 257.293, 257.2929, 257.2936, 257.2934, 257.295, 
    257.2941, 257.2966, 257.2975, 257.3001, 257.3017, 257.3033, 257.3041, 
    257.3043, 257.3044,
  259.794, 259.7949, 259.7947, 259.7953, 259.795, 259.7954, 259.7942, 
    259.7949, 259.7944, 259.7941, 259.7966, 259.7954, 259.798, 259.7972, 
    259.7993, 259.7979, 259.7996, 259.7993, 259.8003, 259.8, 259.8012, 
    259.8004, 259.8019, 259.801, 259.8011, 259.8004, 259.7957, 259.7965, 
    259.7956, 259.7957, 259.7957, 259.795, 259.7946, 259.794, 259.7941, 
    259.7946, 259.7958, 259.7954, 259.7964, 259.7964, 259.7975, 259.797, 
    259.7989, 259.7984, 259.8, 259.7996, 259.8, 259.7998, 259.8, 259.7993, 
    259.7996, 259.7991, 259.7971, 259.7977, 259.7959, 259.7949, 259.7942, 
    259.7938, 259.7938, 259.7939, 259.7946, 259.7952, 259.7957, 259.7961, 
    259.7964, 259.7973, 259.7979, 259.799, 259.7988, 259.7992, 259.7995, 
    259.8001, 259.8, 259.8003, 259.7992, 259.7999, 259.7987, 259.799, 
    259.7964, 259.7955, 259.795, 259.7947, 259.7939, 259.7945, 259.7942, 
    259.7948, 259.7951, 259.795, 259.7961, 259.7956, 259.7979, 259.7969, 
    259.7995, 259.7989, 259.7997, 259.7993, 259.7999, 259.7993, 259.8004, 
    259.8006, 259.8004, 259.8011, 259.7993, 259.8, 259.795, 259.795, 
    259.7951, 259.7945, 259.7945, 259.794, 259.7944, 259.7946, 259.7952, 
    259.7955, 259.7957, 259.7964, 259.7971, 259.7982, 259.7989, 259.7994, 
    259.7991, 259.7994, 259.7991, 259.7989, 259.8005, 259.7996, 259.801, 
    259.8009, 259.8003, 259.8009, 259.795, 259.7948, 259.7943, 259.7947, 
    259.7939, 259.7943, 259.7946, 259.7956, 259.7959, 259.7961, 259.7965, 
    259.797, 259.7979, 259.7988, 259.7996, 259.7995, 259.7995, 259.7997, 
    259.7993, 259.7997, 259.7998, 259.7996, 259.8009, 259.8005, 259.8009, 
    259.8007, 259.7949, 259.7952, 259.795, 259.7953, 259.7951, 259.796, 
    259.7962, 259.7975, 259.797, 259.7978, 259.7971, 259.7972, 259.7978, 
    259.7971, 259.7987, 259.7976, 259.7997, 259.7986, 259.7998, 259.7996, 
    259.7999, 259.8002, 259.8006, 259.8014, 259.8012, 259.8018, 259.7956, 
    259.7959, 259.7959, 259.7963, 259.7966, 259.7972, 259.7982, 259.7978, 
    259.7985, 259.7986, 259.7976, 259.7982, 259.7962, 259.7965, 259.7963, 
    259.7956, 259.7979, 259.7967, 259.7989, 259.7982, 259.8002, 259.7992, 
    259.8011, 259.8019, 259.8027, 259.8036, 259.7961, 259.7959, 259.7964, 
    259.7969, 259.7975, 259.7983, 259.7984, 259.7985, 259.7989, 259.7992, 
    259.7986, 259.7993, 259.7966, 259.798, 259.7958, 259.7964, 259.7969, 
    259.7967, 259.7978, 259.798, 259.799, 259.7985, 259.8017, 259.8003, 
    259.8043, 259.8032, 259.7958, 259.7961, 259.7973, 259.7968, 259.7984, 
    259.7988, 259.7991, 259.7995, 259.7995, 259.7998, 259.7994, 259.7998, 
    259.7983, 259.799, 259.7972, 259.7976, 259.7974, 259.7972, 259.7979, 
    259.7986, 259.7986, 259.7988, 259.7994, 259.7984, 259.8018, 259.7997, 
    259.7965, 259.7971, 259.7972, 259.797, 259.7987, 259.7981, 259.7998, 
    259.7993, 259.8001, 259.7997, 259.7997, 259.7992, 259.7989, 259.7981, 
    259.7975, 259.797, 259.7971, 259.7977, 259.7986, 259.7995, 259.7993, 
    259.8, 259.7982, 259.799, 259.7987, 259.7994, 259.7978, 259.7992, 
    259.7975, 259.7976, 259.7981, 259.799, 259.7993, 259.7995, 259.7993, 
    259.7986, 259.7986, 259.7981, 259.7979, 259.7976, 259.7973, 259.7975, 
    259.7978, 259.7986, 259.7994, 259.8002, 259.8004, 259.8014, 259.8006, 
    259.8019, 259.8008, 259.8027, 259.7993, 259.8008, 259.7981, 259.7984, 
    259.7989, 259.8001, 259.7994, 259.8002, 259.7985, 259.7977, 259.7975, 
    259.7971, 259.7975, 259.7975, 259.7979, 259.7977, 259.7987, 259.7982, 
    259.7997, 259.8002, 259.8018, 259.8027, 259.8038, 259.8042, 259.8044, 
    259.8044,
  262.0097, 262.0099, 262.0099, 262.0101, 262.01, 262.0101, 262.0098, 
    262.0099, 262.0098, 262.0097, 262.0104, 262.0101, 262.0108, 262.0106, 
    262.0111, 262.0107, 262.0112, 262.0111, 262.0114, 262.0113, 262.0117, 
    262.0114, 262.0119, 262.0116, 262.0117, 262.0114, 262.0101, 262.0103, 
    262.0101, 262.0102, 262.0102, 262.01, 262.0099, 262.0097, 262.0097, 
    262.0099, 262.0102, 262.0101, 262.0103, 262.0103, 262.0107, 262.0105, 
    262.011, 262.0109, 262.0113, 262.0112, 262.0113, 262.0113, 262.0113, 
    262.0111, 262.0112, 262.0111, 262.0105, 262.0107, 262.0102, 262.0099, 
    262.0098, 262.0096, 262.0097, 262.0097, 262.0099, 262.01, 262.0102, 
    262.0103, 262.0103, 262.0106, 262.0107, 262.011, 262.011, 262.0111, 
    262.0112, 262.0114, 262.0114, 262.0114, 262.0111, 262.0113, 262.011, 
    262.011, 262.0103, 262.0101, 262.01, 262.0099, 262.0097, 262.0098, 
    262.0098, 262.0099, 262.01, 262.01, 262.0103, 262.0101, 262.0107, 
    262.0105, 262.0112, 262.011, 262.0112, 262.0111, 262.0113, 262.0111, 
    262.0114, 262.0115, 262.0115, 262.0117, 262.0111, 262.0113, 262.01, 
    262.01, 262.01, 262.0099, 262.0099, 262.0097, 262.0098, 262.0099, 262.01, 
    262.0101, 262.0102, 262.0103, 262.0105, 262.0108, 262.011, 262.0112, 
    262.0111, 262.0112, 262.0111, 262.011, 262.0115, 262.0112, 262.0116, 
    262.0116, 262.0114, 262.0116, 262.01, 262.0099, 262.0098, 262.0099, 
    262.0097, 262.0098, 262.0099, 262.0101, 262.0102, 262.0103, 262.0104, 
    262.0105, 262.0108, 262.011, 262.0112, 262.0112, 262.0112, 262.0113, 
    262.0111, 262.0113, 262.0113, 262.0112, 262.0116, 262.0115, 262.0116, 
    262.0115, 262.0099, 262.01, 262.01, 262.01, 262.01, 262.0102, 262.0103, 
    262.0107, 262.0105, 262.0107, 262.0105, 262.0106, 262.0107, 262.0105, 
    262.011, 262.0107, 262.0113, 262.0109, 262.0113, 262.0112, 262.0113, 
    262.0114, 262.0115, 262.0117, 262.0117, 262.0119, 262.0101, 262.0102, 
    262.0102, 262.0103, 262.0104, 262.0106, 262.0108, 262.0107, 262.0109, 
    262.011, 262.0107, 262.0108, 262.0103, 262.0104, 262.0103, 262.0101, 
    262.0107, 262.0104, 262.011, 262.0108, 262.0114, 262.0111, 262.0117, 
    262.0119, 262.0121, 262.0124, 262.0103, 262.0102, 262.0103, 262.0105, 
    262.0107, 262.0109, 262.0109, 262.0109, 262.011, 262.0111, 262.0109, 
    262.0111, 262.0104, 262.0108, 262.0102, 262.0103, 262.0105, 262.0104, 
    262.0107, 262.0108, 262.0111, 262.0109, 262.0118, 262.0114, 262.0126, 
    262.0123, 262.0102, 262.0103, 262.0106, 262.0104, 262.0109, 262.011, 
    262.0111, 262.0112, 262.0112, 262.0113, 262.0112, 262.0113, 262.0109, 
    262.011, 262.0106, 262.0107, 262.0106, 262.0106, 262.0107, 262.0109, 
    262.011, 262.011, 262.0112, 262.0109, 262.0119, 262.0112, 262.0104, 
    262.0105, 262.0106, 262.0105, 262.011, 262.0108, 262.0113, 262.0111, 
    262.0114, 262.0113, 262.0112, 262.0111, 262.011, 262.0108, 262.0107, 
    262.0105, 262.0105, 262.0107, 262.011, 262.0112, 262.0111, 262.0114, 
    262.0108, 262.011, 262.011, 262.0112, 262.0107, 262.0111, 262.0106, 
    262.0107, 262.0108, 262.011, 262.0111, 262.0112, 262.0111, 262.011, 
    262.0109, 262.0108, 262.0107, 262.0107, 262.0106, 262.0107, 262.0107, 
    262.011, 262.0112, 262.0114, 262.0115, 262.0117, 262.0115, 262.0119, 
    262.0115, 262.0121, 262.0111, 262.0115, 262.0108, 262.0109, 262.011, 
    262.0114, 262.0112, 262.0114, 262.0109, 262.0107, 262.0106, 262.0105, 
    262.0106, 262.0106, 262.0107, 262.0107, 262.011, 262.0108, 262.0112, 
    262.0114, 262.0118, 262.0121, 262.0125, 262.0126, 262.0126, 262.0126,
  262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985,
  263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.2737, 263.2855, 263.2832, 263.2927, 263.2874, 263.2936, 263.2761, 
    263.2859, 263.2797, 263.2748, 263.3111, 263.2931, 263.3296, 263.3183, 
    263.3466, 263.3278, 263.3504, 263.3461, 263.3591, 263.3554, 263.3719, 
    263.3608, 263.3806, 263.3693, 263.371, 263.3604, 263.2968, 263.3088, 
    263.2961, 263.2978, 263.297, 263.2875, 263.2828, 263.2728, 263.2746, 
    263.282, 263.2986, 263.2929, 263.3071, 263.3068, 263.3225, 263.3154, 
    263.3416, 263.3342, 263.3555, 263.3502, 263.3553, 263.3537, 263.3553, 
    263.3474, 263.3508, 263.3438, 263.3168, 263.3248, 263.3008, 263.2862, 
    263.2765, 263.2697, 263.2706, 263.2725, 263.282, 263.2909, 263.2977, 
    263.3023, 263.3068, 263.3202, 263.3273, 263.343, 263.3402, 263.345, 
    263.3496, 263.3573, 263.356, 263.3594, 263.3449, 263.3546, 263.3386, 
    263.343, 263.3079, 263.2944, 263.2887, 263.2836, 263.2714, 263.2798, 
    263.2765, 263.2845, 263.2895, 263.287, 263.3024, 263.2964, 263.3277, 
    263.3143, 263.3491, 263.3408, 263.3511, 263.3458, 263.3548, 263.3467, 
    263.3607, 263.3637, 263.3617, 263.3697, 263.3463, 263.3553, 263.287, 
    263.2874, 263.2892, 263.2809, 263.2804, 263.2727, 263.2795, 263.2824, 
    263.2898, 263.2941, 263.2983, 263.3073, 263.3174, 263.3314, 263.3413, 
    263.348, 263.3439, 263.3475, 263.3435, 263.3416, 263.3626, 263.3508, 
    263.3685, 263.3676, 263.3595, 263.3676, 263.2876, 263.2853, 263.2772, 
    263.2835, 263.2719, 263.2784, 263.2821, 263.2965, 263.2997, 263.3026, 
    263.3084, 263.3158, 263.3286, 263.3397, 263.3499, 263.3492, 263.3494, 
    263.3517, 263.346, 263.3526, 263.3537, 263.3508, 263.3674, 263.3627, 
    263.3675, 263.3644, 263.2861, 263.29, 263.2879, 263.2919, 263.289, 
    263.3015, 263.3053, 263.3228, 263.3156, 263.327, 263.3168, 263.3186, 
    263.3273, 263.3174, 263.3391, 263.3244, 263.3517, 263.337, 263.3527, 
    263.3498, 263.3545, 263.3587, 263.364, 263.3737, 263.3715, 263.3796, 
    263.2959, 263.301, 263.3005, 263.3058, 263.3098, 263.3183, 263.3318, 
    263.3268, 263.3361, 263.3379, 263.3238, 263.3325, 263.3044, 263.3089, 
    263.3062, 263.2963, 263.3279, 263.3117, 263.3415, 263.3328, 263.3581, 
    263.3455, 263.3702, 263.3807, 263.3907, 263.4022, 263.3037, 263.3003, 
    263.3065, 263.315, 263.3229, 263.3333, 263.3344, 263.3364, 263.3414, 
    263.3456, 263.3369, 263.3467, 263.31, 263.3293, 263.299, 263.3081, 
    263.3145, 263.3117, 263.3262, 263.3296, 263.3432, 263.3362, 263.3781, 
    263.3596, 263.411, 263.3967, 263.2991, 263.3037, 263.3199, 263.3122, 
    263.334, 263.3394, 263.3437, 263.3492, 263.3498, 263.3531, 263.3477, 
    263.3529, 263.3334, 263.3421, 263.3181, 263.3239, 263.3213, 263.3183, 
    263.3274, 263.3371, 263.3373, 263.3404, 263.3491, 263.3341, 263.3805, 
    263.3518, 263.3088, 263.3177, 263.3191, 263.3156, 263.3388, 263.3304, 
    263.353, 263.3469, 263.3569, 263.352, 263.3512, 263.3448, 263.3409, 
    263.3308, 263.3226, 263.3161, 263.3176, 263.3248, 263.3377, 263.3499, 
    263.3472, 263.3562, 263.3325, 263.3424, 263.3386, 263.3486, 263.3266, 
    263.3452, 263.3218, 263.3239, 263.3303, 263.343, 263.3459, 263.3489, 
    263.3471, 263.338, 263.3365, 263.3301, 263.3283, 263.3235, 263.3194, 
    263.3231, 263.327, 263.338, 263.348, 263.3588, 263.3615, 263.374, 
    263.3637, 263.3806, 263.3662, 263.3912, 263.3464, 263.3658, 263.3306, 
    263.3344, 263.3412, 263.357, 263.3485, 263.3585, 263.3365, 263.325, 
    263.3221, 263.3165, 263.3222, 263.3217, 263.3271, 263.3254, 263.3384, 
    263.3314, 263.3512, 263.3584, 263.3788, 263.3912, 263.4039, 263.4094, 
    263.4111, 263.4118 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9096, 253.9104, 253.9103, 253.911, 253.9106, 253.911, 253.9098, 
    253.9105, 253.91, 253.9097, 253.9123, 253.911, 253.9137, 253.9128, 
    253.9149, 253.9135, 253.9152, 253.9149, 253.9158, 253.9155, 253.9167, 
    253.9159, 253.9174, 253.9165, 253.9167, 253.9159, 253.9113, 253.9121, 
    253.9112, 253.9113, 253.9113, 253.9106, 253.9102, 253.9095, 253.9097, 
    253.9102, 253.9114, 253.911, 253.912, 253.912, 253.9131, 253.9126, 
    253.9145, 253.914, 253.9156, 253.9152, 253.9155, 253.9154, 253.9155, 
    253.915, 253.9152, 253.9147, 253.9127, 253.9133, 253.9116, 253.9105, 
    253.9098, 253.9093, 253.9094, 253.9095, 253.9102, 253.9109, 253.9113, 
    253.9117, 253.912, 253.9129, 253.9135, 253.9146, 253.9144, 253.9148, 
    253.9151, 253.9157, 253.9156, 253.9158, 253.9148, 253.9155, 253.9143, 
    253.9146, 253.912, 253.9111, 253.9107, 253.9103, 253.9094, 253.91, 
    253.9098, 253.9104, 253.9108, 253.9106, 253.9117, 253.9113, 253.9135, 
    253.9125, 253.9151, 253.9145, 253.9152, 253.9148, 253.9155, 253.9149, 
    253.9159, 253.9162, 253.916, 253.9166, 253.9149, 253.9155, 253.9106, 
    253.9106, 253.9107, 253.9101, 253.9101, 253.9095, 253.91, 253.9102, 
    253.9108, 253.9111, 253.9114, 253.912, 253.9128, 253.9138, 253.9145, 
    253.915, 253.9147, 253.915, 253.9147, 253.9145, 253.9161, 253.9152, 
    253.9165, 253.9164, 253.9158, 253.9164, 253.9106, 253.9104, 253.9099, 
    253.9103, 253.9095, 253.9099, 253.9102, 253.9113, 253.9115, 253.9117, 
    253.9121, 253.9127, 253.9136, 253.9144, 253.9151, 253.9151, 253.9151, 
    253.9153, 253.9149, 253.9153, 253.9154, 253.9152, 253.9164, 253.9161, 
    253.9164, 253.9162, 253.9105, 253.9108, 253.9106, 253.9109, 253.9107, 
    253.9116, 253.9119, 253.9131, 253.9126, 253.9135, 253.9127, 253.9129, 
    253.9135, 253.9128, 253.9143, 253.9133, 253.9153, 253.9142, 253.9153, 
    253.9151, 253.9155, 253.9158, 253.9162, 253.9169, 253.9167, 253.9173, 
    253.9112, 253.9116, 253.9115, 253.9119, 253.9122, 253.9128, 253.9138, 
    253.9135, 253.9141, 253.9143, 253.9132, 253.9139, 253.9118, 253.9121, 
    253.912, 253.9112, 253.9135, 253.9124, 253.9145, 253.9139, 253.9157, 
    253.9148, 253.9166, 253.9174, 253.9181, 253.919, 253.9118, 253.9115, 
    253.912, 253.9126, 253.9132, 253.9139, 253.914, 253.9142, 253.9145, 
    253.9148, 253.9142, 253.9149, 253.9122, 253.9136, 253.9114, 253.9121, 
    253.9126, 253.9124, 253.9134, 253.9137, 253.9146, 253.9141, 253.9172, 
    253.9158, 253.9196, 253.9186, 253.9115, 253.9118, 253.9129, 253.9124, 
    253.914, 253.9144, 253.9147, 253.9151, 253.9151, 253.9154, 253.915, 
    253.9154, 253.9139, 253.9146, 253.9128, 253.9133, 253.9131, 253.9128, 
    253.9135, 253.9142, 253.9142, 253.9144, 253.915, 253.914, 253.9173, 
    253.9152, 253.9122, 253.9128, 253.9129, 253.9126, 253.9143, 253.9137, 
    253.9154, 253.9149, 253.9157, 253.9153, 253.9152, 253.9148, 253.9145, 
    253.9137, 253.9131, 253.9127, 253.9128, 253.9133, 253.9142, 253.9151, 
    253.9149, 253.9156, 253.9139, 253.9146, 253.9143, 253.915, 253.9134, 
    253.9148, 253.9131, 253.9133, 253.9137, 253.9146, 253.9149, 253.9151, 
    253.9149, 253.9143, 253.9142, 253.9137, 253.9136, 253.9132, 253.9129, 
    253.9132, 253.9135, 253.9143, 253.915, 253.9158, 253.916, 253.9169, 
    253.9161, 253.9173, 253.9163, 253.9181, 253.9149, 253.9163, 253.9137, 
    253.914, 253.9145, 253.9156, 253.915, 253.9158, 253.9142, 253.9133, 
    253.9131, 253.9127, 253.9131, 253.9131, 253.9135, 253.9134, 253.9143, 
    253.9138, 253.9152, 253.9158, 253.9173, 253.9182, 253.9191, 253.9195, 
    253.9196, 253.9197 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1456412, 0.1456404, 0.1456405, 0.1456398, 0.1456402, 0.1456398, 0.145641, 
    0.1456403, 0.1456408, 0.1456411, 0.1456386, 0.1456398, 0.1456374, 
    0.1456381, 0.1456363, 0.1456375, 0.1456361, 0.1456363, 0.1456356, 
    0.1456358, 0.145635, 0.1456355, 0.1456345, 0.1456351, 0.145635, 
    0.1456355, 0.1456396, 0.1456387, 0.1456396, 0.1456395, 0.1456395, 
    0.1456402, 0.1456406, 0.1456413, 0.1456411, 0.1456406, 0.1456394, 
    0.1456398, 0.1456388, 0.1456389, 0.1456378, 0.1456383, 0.1456366, 
    0.1456371, 0.1456358, 0.1456361, 0.1456358, 0.1456359, 0.1456358, 
    0.1456363, 0.1456361, 0.1456365, 0.1456382, 0.1456377, 0.1456393, 
    0.1456403, 0.145641, 0.1456415, 0.1456414, 0.1456413, 0.1456406, 0.14564, 
    0.1456395, 0.1456392, 0.1456389, 0.145638, 0.1456375, 0.1456365, 
    0.1456367, 0.1456364, 0.1456361, 0.1456357, 0.1456358, 0.1456356, 
    0.1456364, 0.1456359, 0.1456368, 0.1456365, 0.1456388, 0.1456397, 
    0.1456401, 0.1456405, 0.1456414, 0.1456408, 0.145641, 0.1456404, 
    0.1456401, 0.1456402, 0.1456392, 0.1456396, 0.1456375, 0.1456384, 
    0.1456362, 0.1456367, 0.1456361, 0.1456364, 0.1456359, 0.1456363, 
    0.1456355, 0.1456354, 0.1456355, 0.1456351, 0.1456363, 0.1456358, 
    0.1456402, 0.1456402, 0.1456401, 0.1456407, 0.1456407, 0.1456413, 
    0.1456408, 0.1456406, 0.14564, 0.1456397, 0.1456394, 0.1456388, 
    0.1456382, 0.1456373, 0.1456366, 0.1456362, 0.1456365, 0.1456363, 
    0.1456365, 0.1456366, 0.1456354, 0.1456361, 0.1456351, 0.1456352, 
    0.1456356, 0.1456352, 0.1456402, 0.1456404, 0.145641, 0.1456405, 
    0.1456414, 0.1456409, 0.1456406, 0.1456396, 0.1456393, 0.1456392, 
    0.1456388, 0.1456383, 0.1456374, 0.1456367, 0.1456361, 0.1456362, 
    0.1456362, 0.145636, 0.1456363, 0.145636, 0.1456359, 0.1456361, 
    0.1456352, 0.1456354, 0.1456352, 0.1456353, 0.1456403, 0.14564, 
    0.1456402, 0.1456399, 0.1456401, 0.1456392, 0.145639, 0.1456378, 
    0.1456383, 0.1456375, 0.1456382, 0.1456381, 0.1456375, 0.1456382, 
    0.1456368, 0.1456377, 0.145636, 0.1456369, 0.145636, 0.1456361, 
    0.1456359, 0.1456356, 0.1456354, 0.1456349, 0.145635, 0.1456346, 
    0.1456396, 0.1456393, 0.1456393, 0.1456389, 0.1456387, 0.1456381, 
    0.1456372, 0.1456376, 0.145637, 0.1456369, 0.1456378, 0.1456372, 
    0.145639, 0.1456387, 0.1456389, 0.1456396, 0.1456375, 0.1456385, 
    0.1456366, 0.1456372, 0.1456357, 0.1456364, 0.145635, 0.1456345, 
    0.1456341, 0.1456336, 0.1456391, 0.1456393, 0.1456389, 0.1456383, 
    0.1456378, 0.1456371, 0.1456371, 0.145637, 0.1456366, 0.1456364, 
    0.1456369, 0.1456363, 0.1456387, 0.1456374, 0.1456394, 0.1456388, 
    0.1456383, 0.1456385, 0.1456376, 0.1456374, 0.1456365, 0.145637, 
    0.1456347, 0.1456356, 0.1456333, 0.1456338, 0.1456394, 0.1456391, 
    0.145638, 0.1456385, 0.1456371, 0.1456368, 0.1456365, 0.1456362, 
    0.1456361, 0.1456359, 0.1456362, 0.145636, 0.1456371, 0.1456366, 
    0.1456381, 0.1456377, 0.1456379, 0.1456381, 0.1456375, 0.1456369, 
    0.1456369, 0.1456367, 0.1456362, 0.1456371, 0.1456345, 0.145636, 
    0.1456387, 0.1456381, 0.145638, 0.1456383, 0.1456368, 0.1456373, 
    0.1456359, 0.1456363, 0.1456357, 0.145636, 0.1456361, 0.1456364, 
    0.1456366, 0.1456373, 0.1456378, 0.1456382, 0.1456382, 0.1456377, 
    0.1456369, 0.1456361, 0.1456363, 0.1456358, 0.1456372, 0.1456366, 
    0.1456368, 0.1456362, 0.1456376, 0.1456364, 0.1456379, 0.1456377, 
    0.1456373, 0.1456365, 0.1456363, 0.1456362, 0.1456363, 0.1456369, 
    0.1456369, 0.1456373, 0.1456375, 0.1456378, 0.145638, 0.1456378, 
    0.1456375, 0.1456369, 0.1456362, 0.1456356, 0.1456355, 0.1456349, 
    0.1456354, 0.1456345, 0.1456352, 0.1456341, 0.1456363, 0.1456353, 
    0.1456373, 0.1456371, 0.1456366, 0.1456357, 0.1456362, 0.1456356, 
    0.1456369, 0.1456377, 0.1456379, 0.1456382, 0.1456379, 0.1456379, 
    0.1456375, 0.1456376, 0.1456368, 0.1456373, 0.1456361, 0.1456357, 
    0.1456346, 0.1456341, 0.1456336, 0.1456334, 0.1456333, 0.1456333,
  0.1512734, 0.1512782, 0.1512772, 0.151281, 0.151279, 0.1512814, 0.1512744, 
    0.1512783, 0.1512758, 0.1512739, 0.1512883, 0.1512812, 0.151296, 
    0.1512914, 0.1513031, 0.1512952, 0.1513047, 0.1513029, 0.1513084, 
    0.1513069, 0.1513138, 0.1513092, 0.1513175, 0.1513127, 0.1513134, 
    0.151309, 0.1512827, 0.1512874, 0.1512824, 0.1512831, 0.1512828, 
    0.151279, 0.151277, 0.1512731, 0.1512738, 0.1512767, 0.1512834, 
    0.1512812, 0.1512869, 0.1512868, 0.1512931, 0.1512903, 0.151301, 
    0.151298, 0.1513069, 0.1513047, 0.1513068, 0.1513062, 0.1513068, 
    0.1513035, 0.1513049, 0.151302, 0.1512908, 0.1512941, 0.1512843, 
    0.1512783, 0.1512746, 0.1512718, 0.1512722, 0.151273, 0.1512767, 
    0.1512804, 0.1512831, 0.1512849, 0.1512868, 0.1512921, 0.1512951, 
    0.1513016, 0.1513005, 0.1513025, 0.1513044, 0.1513077, 0.1513072, 
    0.1513086, 0.1513025, 0.1513065, 0.1512999, 0.1513017, 0.151287, 
    0.1512818, 0.1512793, 0.1512774, 0.1512725, 0.1512759, 0.1512746, 
    0.1512778, 0.1512798, 0.1512788, 0.151285, 0.1512826, 0.1512952, 
    0.1512898, 0.1513042, 0.1513007, 0.151305, 0.1513029, 0.1513066, 
    0.1513032, 0.1513091, 0.1513104, 0.1513095, 0.1513129, 0.151303, 
    0.1513068, 0.1512788, 0.1512789, 0.1512797, 0.1512763, 0.1512761, 
    0.1512731, 0.1512758, 0.1512769, 0.1512799, 0.1512817, 0.1512833, 
    0.151287, 0.151291, 0.1512968, 0.151301, 0.1513038, 0.1513021, 0.1513036, 
    0.1513019, 0.1513011, 0.1513099, 0.1513049, 0.1513124, 0.151312, 
    0.1513086, 0.1513121, 0.151279, 0.1512781, 0.1512748, 0.1512774, 
    0.1512728, 0.1512753, 0.1512768, 0.1512826, 0.1512839, 0.1512851, 
    0.1512874, 0.1512904, 0.1512957, 0.1513003, 0.1513046, 0.1513043, 
    0.1513044, 0.1513053, 0.1513029, 0.1513057, 0.1513061, 0.1513049, 
    0.1513119, 0.1513099, 0.151312, 0.1513107, 0.1512784, 0.15128, 0.1512791, 
    0.1512807, 0.1512796, 0.1512846, 0.1512861, 0.1512932, 0.1512903, 
    0.151295, 0.1512908, 0.1512915, 0.151295, 0.1512911, 0.1513, 0.1512938, 
    0.1513053, 0.1512991, 0.1513057, 0.1513045, 0.1513065, 0.1513083, 
    0.1513105, 0.1513146, 0.1513136, 0.1513171, 0.1512824, 0.1512844, 
    0.1512842, 0.1512864, 0.151288, 0.1512915, 0.151297, 0.1512949, 
    0.1512988, 0.1512996, 0.1512937, 0.1512973, 0.1512858, 0.1512876, 
    0.1512865, 0.1512825, 0.1512953, 0.1512887, 0.151301, 0.1512974, 
    0.151308, 0.1513027, 0.1513131, 0.1513175, 0.1513219, 0.1513268, 
    0.1512855, 0.1512841, 0.1512867, 0.15129, 0.1512933, 0.1512976, 
    0.1512981, 0.1512989, 0.151301, 0.1513028, 0.1512991, 0.1513032, 
    0.1512879, 0.1512959, 0.1512836, 0.1512872, 0.1512899, 0.1512888, 
    0.1512947, 0.1512961, 0.1513017, 0.1512989, 0.1513164, 0.1513086, 
    0.1513307, 0.1513244, 0.1512837, 0.1512855, 0.1512921, 0.151289, 
    0.151298, 0.1513002, 0.151302, 0.1513042, 0.1513045, 0.1513059, 
    0.1513037, 0.1513058, 0.1512976, 0.1513013, 0.1512914, 0.1512938, 
    0.1512927, 0.1512915, 0.1512952, 0.1512991, 0.1512993, 0.1513005, 
    0.1513039, 0.151298, 0.1513172, 0.1513051, 0.1512876, 0.1512911, 
    0.1512917, 0.1512904, 0.1512999, 0.1512964, 0.1513059, 0.1513033, 
    0.1513075, 0.1513054, 0.1513051, 0.1513024, 0.1513008, 0.1512966, 
    0.1512932, 0.1512906, 0.1512912, 0.1512941, 0.1512994, 0.1513045, 
    0.1513034, 0.1513072, 0.1512973, 0.1513014, 0.1512998, 0.151304, 
    0.1512949, 0.1513024, 0.1512929, 0.1512938, 0.1512964, 0.1513016, 
    0.1513029, 0.1513041, 0.1513034, 0.1512996, 0.151299, 0.1512963, 
    0.1512956, 0.1512936, 0.1512919, 0.1512934, 0.151295, 0.1512996, 
    0.1513037, 0.1513083, 0.1513094, 0.1513146, 0.1513103, 0.1513173, 
    0.1513111, 0.1513219, 0.1513029, 0.1513111, 0.1512965, 0.1512981, 
    0.1513009, 0.1513075, 0.151304, 0.1513081, 0.151299, 0.1512941, 0.151293, 
    0.1512907, 0.1512931, 0.1512929, 0.1512951, 0.1512944, 0.1512998, 
    0.1512969, 0.1513051, 0.1513081, 0.1513167, 0.151322, 0.1513276, 0.15133, 
    0.1513307, 0.1513311,
  0.1611242, 0.1611302, 0.161129, 0.1611339, 0.1611312, 0.1611344, 0.1611254, 
    0.1611304, 0.1611273, 0.1611248, 0.1611432, 0.1611341, 0.161153, 
    0.1611471, 0.1611622, 0.1611521, 0.1611642, 0.161162, 0.161169, 0.161167, 
    0.1611759, 0.16117, 0.1611807, 0.1611745, 0.1611754, 0.1611697, 0.161136, 
    0.161142, 0.1611356, 0.1611365, 0.1611361, 0.1611312, 0.1611287, 
    0.1611238, 0.1611247, 0.1611284, 0.1611369, 0.161134, 0.1611414, 
    0.1611412, 0.1611494, 0.1611457, 0.1611595, 0.1611556, 0.1611671, 
    0.1611642, 0.1611669, 0.1611661, 0.1611669, 0.1611627, 0.1611645, 
    0.1611608, 0.1611464, 0.1611505, 0.161138, 0.1611304, 0.1611256, 
    0.1611222, 0.1611227, 0.1611236, 0.1611284, 0.161133, 0.1611365, 
    0.1611389, 0.1611412, 0.161148, 0.1611518, 0.1611603, 0.1611588, 
    0.1611613, 0.1611639, 0.161168, 0.1611674, 0.1611692, 0.1611613, 
    0.1611665, 0.161158, 0.1611603, 0.1611415, 0.1611348, 0.1611317, 
    0.1611293, 0.161123, 0.1611273, 0.1611256, 0.1611297, 0.1611323, 
    0.161131, 0.1611389, 0.1611358, 0.161152, 0.161145, 0.1611636, 0.1611591, 
    0.1611647, 0.1611619, 0.1611667, 0.1611623, 0.1611699, 0.1611715, 
    0.1611704, 0.1611748, 0.1611621, 0.1611669, 0.161131, 0.1611312, 
    0.1611322, 0.1611278, 0.1611276, 0.1611237, 0.1611272, 0.1611287, 
    0.1611325, 0.1611347, 0.1611368, 0.1611415, 0.1611466, 0.161154, 
    0.1611594, 0.161163, 0.1611608, 0.1611628, 0.1611606, 0.1611596, 
    0.1611709, 0.1611645, 0.1611741, 0.1611736, 0.1611692, 0.1611737, 
    0.1611313, 0.1611302, 0.161126, 0.1611293, 0.1611233, 0.1611266, 
    0.1611284, 0.1611358, 0.1611376, 0.161139, 0.161142, 0.1611459, 
    0.1611526, 0.1611585, 0.161164, 0.1611636, 0.1611638, 0.161165, 0.161162, 
    0.1611655, 0.161166, 0.1611645, 0.1611735, 0.161171, 0.1611736, 
    0.1611719, 0.1611305, 0.1611325, 0.1611315, 0.1611335, 0.161132, 
    0.1611384, 0.1611403, 0.1611494, 0.1611458, 0.1611517, 0.1611464, 
    0.1611473, 0.1611518, 0.1611467, 0.1611581, 0.1611502, 0.161165, 
    0.161157, 0.1611655, 0.161164, 0.1611665, 0.1611688, 0.1611717, 
    0.1611769, 0.1611757, 0.1611802, 0.1611356, 0.1611381, 0.161138, 
    0.1611407, 0.1611427, 0.1611472, 0.1611543, 0.1611517, 0.1611566, 
    0.1611576, 0.1611501, 0.1611546, 0.1611399, 0.1611422, 0.1611409, 
    0.1611357, 0.1611522, 0.1611437, 0.1611595, 0.1611549, 0.1611685, 
    0.1611616, 0.1611751, 0.1611807, 0.1611864, 0.1611926, 0.1611396, 
    0.1611378, 0.1611411, 0.1611454, 0.1611496, 0.1611551, 0.1611557, 
    0.1611568, 0.1611595, 0.1611617, 0.161157, 0.1611623, 0.1611426, 
    0.161153, 0.1611371, 0.1611418, 0.1611452, 0.1611437, 0.1611514, 
    0.1611532, 0.1611604, 0.1611567, 0.1611792, 0.1611692, 0.1611977, 
    0.1611896, 0.1611372, 0.1611396, 0.161148, 0.161144, 0.1611555, 
    0.1611584, 0.1611607, 0.1611636, 0.161164, 0.1611657, 0.1611629, 
    0.1611657, 0.1611551, 0.1611598, 0.1611471, 0.1611501, 0.1611488, 
    0.1611472, 0.161152, 0.1611571, 0.1611573, 0.1611589, 0.1611633, 
    0.1611556, 0.1611804, 0.1611648, 0.1611423, 0.1611468, 0.1611476, 
    0.1611458, 0.1611581, 0.1611536, 0.1611657, 0.1611625, 0.1611678, 
    0.1611651, 0.1611647, 0.1611613, 0.1611592, 0.1611538, 0.1611494, 
    0.1611461, 0.1611468, 0.1611506, 0.1611574, 0.161164, 0.1611625, 
    0.1611674, 0.1611547, 0.1611599, 0.1611579, 0.1611633, 0.1611516, 
    0.1611613, 0.1611491, 0.1611501, 0.1611535, 0.1611602, 0.1611619, 
    0.1611635, 0.1611625, 0.1611576, 0.1611568, 0.1611535, 0.1611525, 
    0.1611499, 0.1611478, 0.1611497, 0.1611517, 0.1611577, 0.1611629, 
    0.1611688, 0.1611703, 0.1611769, 0.1611714, 0.1611804, 0.1611725, 
    0.1611864, 0.161162, 0.1611725, 0.1611537, 0.1611557, 0.1611593, 
    0.1611678, 0.1611633, 0.1611686, 0.1611568, 0.1611506, 0.1611492, 
    0.1611462, 0.1611492, 0.161149, 0.1611519, 0.161151, 0.1611578, 
    0.1611542, 0.1611647, 0.1611686, 0.1611797, 0.1611865, 0.1611937, 
    0.1611968, 0.1611978, 0.1611982,
  0.175334, 0.1753385, 0.1753376, 0.1753412, 0.1753393, 0.1753416, 0.1753349, 
    0.1753386, 0.1753363, 0.1753344, 0.1753483, 0.1753414, 0.1753558, 
    0.1753513, 0.1753628, 0.1753551, 0.1753644, 0.1753627, 0.1753681, 
    0.1753666, 0.1753735, 0.1753689, 0.1753772, 0.1753724, 0.1753732, 
    0.1753687, 0.1753429, 0.1753474, 0.1753426, 0.1753432, 0.1753429, 
    0.1753393, 0.1753374, 0.1753337, 0.1753344, 0.1753371, 0.1753435, 
    0.1753414, 0.1753469, 0.1753468, 0.175353, 0.1753502, 0.1753608, 
    0.1753578, 0.1753667, 0.1753644, 0.1753665, 0.1753659, 0.1753665, 
    0.1753632, 0.1753646, 0.1753618, 0.1753507, 0.1753539, 0.1753444, 
    0.1753386, 0.1753351, 0.1753325, 0.1753328, 0.1753335, 0.1753371, 
    0.1753406, 0.1753432, 0.175345, 0.1753468, 0.1753519, 0.1753549, 
    0.1753614, 0.1753603, 0.1753622, 0.1753642, 0.1753674, 0.1753669, 
    0.1753683, 0.1753622, 0.1753662, 0.1753596, 0.1753614, 0.175347, 
    0.175342, 0.1753396, 0.1753378, 0.1753331, 0.1753363, 0.175335, 
    0.1753381, 0.1753401, 0.1753391, 0.1753451, 0.1753427, 0.175355, 
    0.1753497, 0.1753639, 0.1753605, 0.1753648, 0.1753626, 0.1753663, 
    0.175363, 0.1753688, 0.1753701, 0.1753692, 0.1753726, 0.1753628, 
    0.1753665, 0.1753391, 0.1753392, 0.17534, 0.1753367, 0.1753365, 
    0.1753336, 0.1753362, 0.1753373, 0.1753402, 0.1753418, 0.1753434, 
    0.175347, 0.1753509, 0.1753566, 0.1753607, 0.1753635, 0.1753618, 
    0.1753633, 0.1753616, 0.1753608, 0.1753696, 0.1753646, 0.1753721, 
    0.1753717, 0.1753683, 0.1753718, 0.1753393, 0.1753384, 0.1753353, 
    0.1753378, 0.1753333, 0.1753358, 0.1753372, 0.1753427, 0.175344, 
    0.1753451, 0.1753474, 0.1753503, 0.1753555, 0.17536, 0.1753643, 0.175364, 
    0.1753641, 0.175365, 0.1753627, 0.1753654, 0.1753658, 0.1753647, 
    0.1753717, 0.1753697, 0.1753717, 0.1753704, 0.1753387, 0.1753403, 
    0.1753394, 0.175341, 0.1753399, 0.1753447, 0.1753461, 0.1753531, 
    0.1753503, 0.1753548, 0.1753507, 0.1753514, 0.1753548, 0.175351, 
    0.1753597, 0.1753537, 0.175365, 0.1753588, 0.1753654, 0.1753643, 
    0.1753662, 0.175368, 0.1753702, 0.1753743, 0.1753734, 0.1753769, 
    0.1753425, 0.1753445, 0.1753443, 0.1753464, 0.175348, 0.1753514, 
    0.1753568, 0.1753547, 0.1753586, 0.1753593, 0.1753536, 0.175357, 
    0.1753458, 0.1753476, 0.1753466, 0.1753426, 0.1753552, 0.1753487, 
    0.1753608, 0.1753572, 0.1753677, 0.1753624, 0.1753729, 0.1753773, 
    0.1753817, 0.1753867, 0.1753456, 0.1753442, 0.1753467, 0.17535, 
    0.1753532, 0.1753574, 0.1753579, 0.1753587, 0.1753608, 0.1753625, 
    0.1753589, 0.175363, 0.1753479, 0.1753557, 0.1753437, 0.1753472, 
    0.1753498, 0.1753487, 0.1753545, 0.1753559, 0.1753615, 0.1753586, 
    0.1753761, 0.1753683, 0.1753907, 0.1753843, 0.1753438, 0.1753456, 
    0.1753519, 0.1753489, 0.1753577, 0.1753599, 0.1753617, 0.175364, 
    0.1753643, 0.1753656, 0.1753634, 0.1753655, 0.1753574, 0.175361, 
    0.1753513, 0.1753536, 0.1753525, 0.1753514, 0.175355, 0.1753589, 
    0.1753591, 0.1753603, 0.1753637, 0.1753578, 0.175377, 0.1753649, 
    0.1753476, 0.175351, 0.1753516, 0.1753503, 0.1753597, 0.1753562, 
    0.1753656, 0.1753631, 0.1753672, 0.1753651, 0.1753648, 0.1753622, 
    0.1753605, 0.1753564, 0.1753531, 0.1753505, 0.1753511, 0.1753539, 
    0.1753592, 0.1753643, 0.1753631, 0.1753669, 0.1753571, 0.1753611, 
    0.1753595, 0.1753637, 0.1753547, 0.1753621, 0.1753528, 0.1753536, 
    0.1753562, 0.1753614, 0.1753626, 0.1753639, 0.1753631, 0.1753593, 
    0.1753587, 0.1753561, 0.1753554, 0.1753534, 0.1753518, 0.1753533, 
    0.1753548, 0.1753594, 0.1753635, 0.175368, 0.1753691, 0.1753743, 0.17537, 
    0.1753771, 0.1753709, 0.1753817, 0.1753627, 0.1753709, 0.1753563, 
    0.1753579, 0.1753606, 0.1753672, 0.1753637, 0.1753678, 0.1753587, 
    0.175354, 0.1753529, 0.1753506, 0.1753529, 0.1753527, 0.1753549, 
    0.1753542, 0.1753595, 0.1753567, 0.1753648, 0.1753678, 0.1753765, 
    0.1753819, 0.1753875, 0.17539, 0.1753908, 0.1753911,
  0.1899463, 0.1899477, 0.1899474, 0.1899485, 0.1899479, 0.1899487, 
    0.1899466, 0.1899477, 0.189947, 0.1899465, 0.1899508, 0.1899486, 
    0.1899533, 0.1899518, 0.1899556, 0.189953, 0.1899562, 0.1899556, 
    0.1899575, 0.1899569, 0.1899593, 0.1899577, 0.1899607, 0.1899589, 
    0.1899592, 0.1899576, 0.1899491, 0.1899505, 0.189949, 0.1899492, 
    0.1899491, 0.1899479, 0.1899474, 0.1899462, 0.1899464, 0.1899473, 
    0.1899493, 0.1899486, 0.1899504, 0.1899503, 0.1899523, 0.1899514, 
    0.1899549, 0.1899539, 0.1899569, 0.1899561, 0.1899569, 0.1899567, 
    0.1899569, 0.1899558, 0.1899562, 0.1899552, 0.1899516, 0.1899526, 
    0.1899495, 0.1899477, 0.1899467, 0.1899459, 0.189946, 0.1899462, 
    0.1899473, 0.1899484, 0.1899492, 0.1899498, 0.1899503, 0.189952, 
    0.1899529, 0.1899551, 0.1899547, 0.1899554, 0.1899561, 0.1899572, 
    0.189957, 0.1899575, 0.1899554, 0.1899568, 0.1899545, 0.1899551, 
    0.1899504, 0.1899488, 0.189948, 0.1899475, 0.1899461, 0.189947, 
    0.1899466, 0.1899476, 0.1899482, 0.1899479, 0.1899498, 0.189949, 
    0.189953, 0.1899513, 0.189956, 0.1899548, 0.1899563, 0.1899555, 
    0.1899568, 0.1899557, 0.1899577, 0.1899581, 0.1899578, 0.189959, 
    0.1899556, 0.1899569, 0.1899479, 0.1899479, 0.1899482, 0.1899471, 
    0.1899471, 0.1899462, 0.189947, 0.1899473, 0.1899482, 0.1899487, 
    0.1899492, 0.1899504, 0.1899516, 0.1899535, 0.1899549, 0.1899558, 
    0.1899553, 0.1899558, 0.1899552, 0.1899549, 0.1899579, 0.1899562, 
    0.1899588, 0.1899587, 0.1899575, 0.1899587, 0.189948, 0.1899477, 
    0.1899467, 0.1899475, 0.1899461, 0.1899469, 0.1899473, 0.189949, 
    0.1899494, 0.1899498, 0.1899505, 0.1899514, 0.1899531, 0.1899547, 
    0.1899561, 0.189956, 0.189956, 0.1899564, 0.1899556, 0.1899565, 
    0.1899567, 0.1899562, 0.1899587, 0.189958, 0.1899587, 0.1899582, 
    0.1899478, 0.1899482, 0.189948, 0.1899485, 0.1899481, 0.1899496, 
    0.1899501, 0.1899523, 0.1899514, 0.1899529, 0.1899516, 0.1899518, 
    0.1899529, 0.1899517, 0.1899546, 0.1899525, 0.1899564, 0.1899543, 
    0.1899565, 0.1899561, 0.1899568, 0.1899574, 0.1899582, 0.1899596, 
    0.1899593, 0.1899605, 0.189949, 0.1899496, 0.1899495, 0.1899502, 
    0.1899507, 0.1899518, 0.1899536, 0.1899529, 0.1899542, 0.1899544, 
    0.1899525, 0.1899537, 0.18995, 0.1899506, 0.1899502, 0.189949, 0.189953, 
    0.1899509, 0.1899549, 0.1899537, 0.1899573, 0.1899555, 0.1899591, 
    0.1899607, 0.1899623, 0.1899641, 0.1899499, 0.1899495, 0.1899503, 
    0.1899513, 0.1899524, 0.1899538, 0.1899539, 0.1899542, 0.1899549, 
    0.1899555, 0.1899543, 0.1899557, 0.1899506, 0.1899532, 0.1899493, 
    0.1899505, 0.1899513, 0.1899509, 0.1899528, 0.1899533, 0.1899551, 
    0.1899542, 0.1899603, 0.1899575, 0.1899656, 0.1899632, 0.1899493, 
    0.1899499, 0.189952, 0.189951, 0.1899539, 0.1899546, 0.1899552, 0.189956, 
    0.1899561, 0.1899566, 0.1899558, 0.1899565, 0.1899538, 0.189955, 
    0.1899518, 0.1899525, 0.1899522, 0.1899518, 0.189953, 0.1899543, 
    0.1899543, 0.1899548, 0.1899559, 0.1899539, 0.1899606, 0.1899563, 
    0.1899506, 0.1899517, 0.1899519, 0.1899514, 0.1899545, 0.1899534, 
    0.1899566, 0.1899557, 0.1899571, 0.1899564, 0.1899563, 0.1899554, 
    0.1899548, 0.1899534, 0.1899523, 0.1899515, 0.1899517, 0.1899526, 
    0.1899544, 0.1899561, 0.1899557, 0.189957, 0.1899537, 0.189955, 
    0.1899545, 0.1899559, 0.1899529, 0.1899554, 0.1899523, 0.1899525, 
    0.1899534, 0.1899551, 0.1899555, 0.189956, 0.1899557, 0.1899544, 
    0.1899542, 0.1899534, 0.1899531, 0.1899525, 0.1899519, 0.1899524, 
    0.1899529, 0.1899544, 0.1899558, 0.1899574, 0.1899578, 0.1899596, 
    0.1899581, 0.1899606, 0.1899584, 0.1899623, 0.1899556, 0.1899584, 
    0.1899534, 0.1899539, 0.1899549, 0.1899571, 0.1899559, 0.1899573, 
    0.1899542, 0.1899526, 0.1899523, 0.1899516, 0.1899523, 0.1899522, 
    0.189953, 0.1899527, 0.1899545, 0.1899535, 0.1899563, 0.1899573, 
    0.1899604, 0.1899623, 0.1899644, 0.1899653, 0.1899656, 0.1899657,
  0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.197319, 0.197319, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.197319, 0.1973189, 0.197319, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 
    0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.197319, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.197319, 0.1973191, 0.1973192, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 0.1973193, 
    0.1973191, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 
    0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.197319, 0.1973189, 0.197319, 0.1973189, 
    0.1973191, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 
    0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973191, 0.1973192, 
    0.1973193, 0.1973193, 0.1973193,
  0.1984799, 0.1984798, 0.1984799, 0.1984798, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984797, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 
    0.1984799, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984798, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984796, 
    0.1984796, 0.1984796,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.611716, 5.611768, 5.611758, 5.6118, 5.611777, 5.611804, 5.611727, 
    5.61177, 5.611742, 5.611721, 5.611879, 5.611802, 5.611963, 5.611914, 
    5.612042, 5.611955, 5.61206, 5.612041, 5.612102, 5.612084, 5.612159, 
    5.61211, 5.6122, 5.612148, 5.612156, 5.612108, 5.611819, 5.611869, 
    5.611815, 5.611823, 5.61182, 5.611777, 5.611755, 5.611712, 5.611721, 
    5.611753, 5.611826, 5.611802, 5.611865, 5.611864, 5.611932, 5.611901, 
    5.612019, 5.611985, 5.612085, 5.61206, 5.612083, 5.612077, 5.612084, 
    5.612047, 5.612062, 5.61203, 5.611907, 5.611942, 5.611836, 5.61177, 
    5.611729, 5.611698, 5.611702, 5.611711, 5.611753, 5.611793, 5.611823, 
    5.611844, 5.611863, 5.61192, 5.611953, 5.612025, 5.612012, 5.612035, 
    5.612057, 5.612093, 5.612087, 5.612103, 5.612035, 5.61208, 5.612005, 
    5.612026, 5.611865, 5.611808, 5.611781, 5.61176, 5.611706, 5.611743, 
    5.611728, 5.611764, 5.611786, 5.611776, 5.611844, 5.611817, 5.611955, 
    5.611896, 5.612055, 5.612015, 5.612064, 5.61204, 5.612081, 5.612044, 
    5.612109, 5.612123, 5.612113, 5.612151, 5.612041, 5.612083, 5.611775, 
    5.611777, 5.611785, 5.611748, 5.611745, 5.611712, 5.611742, 5.611755, 
    5.611788, 5.611807, 5.611825, 5.611866, 5.611909, 5.611972, 5.612018, 
    5.61205, 5.612031, 5.612048, 5.612029, 5.61202, 5.612117, 5.612062, 
    5.612145, 5.612141, 5.612103, 5.612141, 5.611778, 5.611768, 5.611732, 
    5.61176, 5.611708, 5.611737, 5.611753, 5.611817, 5.611832, 5.611845, 
    5.61187, 5.611903, 5.611959, 5.61201, 5.612059, 5.612055, 5.612056, 
    5.612067, 5.612041, 5.612071, 5.612076, 5.612063, 5.61214, 5.612118, 
    5.612141, 5.612126, 5.611772, 5.611789, 5.611779, 5.611797, 5.611784, 
    5.611839, 5.611856, 5.611933, 5.611902, 5.611952, 5.611907, 5.611915, 
    5.611952, 5.61191, 5.612006, 5.611939, 5.612067, 5.611996, 5.612072, 
    5.612059, 5.612081, 5.6121, 5.612124, 5.612168, 5.612158, 5.612196, 
    5.611815, 5.611837, 5.611835, 5.611859, 5.611876, 5.611914, 5.611974, 
    5.611952, 5.611994, 5.612002, 5.611939, 5.611977, 5.611852, 5.611872, 
    5.611861, 5.611816, 5.611956, 5.611884, 5.612019, 5.611979, 5.612097, 
    5.612037, 5.612153, 5.6122, 5.612247, 5.612298, 5.61185, 5.611835, 
    5.611862, 5.611899, 5.611935, 5.611981, 5.611986, 5.611995, 5.612019, 
    5.612039, 5.611997, 5.612044, 5.611875, 5.611963, 5.611828, 5.611868, 
    5.611897, 5.611885, 5.611949, 5.611965, 5.612026, 5.611994, 5.612187, 
    5.612103, 5.612339, 5.612273, 5.611829, 5.61185, 5.611921, 5.611887, 
    5.611985, 5.612008, 5.61203, 5.612055, 5.612058, 5.612073, 5.612049, 
    5.612073, 5.611981, 5.612021, 5.611914, 5.611939, 5.611928, 5.611914, 
    5.611955, 5.611997, 5.611999, 5.612013, 5.612051, 5.611985, 5.612196, 
    5.612064, 5.611872, 5.61191, 5.611917, 5.611902, 5.612006, 5.611968, 
    5.612073, 5.612045, 5.612092, 5.612068, 5.612065, 5.612035, 5.612016, 
    5.611969, 5.611933, 5.611905, 5.611911, 5.611943, 5.612, 5.612058, 
    5.612045, 5.612088, 5.611978, 5.612022, 5.612004, 5.612052, 5.611951, 
    5.612033, 5.61193, 5.611939, 5.611968, 5.612025, 5.61204, 5.612054, 
    5.612046, 5.612001, 5.611995, 5.611967, 5.611959, 5.611938, 5.611919, 
    5.611936, 5.611952, 5.612002, 5.612049, 5.6121, 5.612113, 5.612168, 
    5.612121, 5.612196, 5.61213, 5.612246, 5.61204, 5.61213, 5.611969, 
    5.611986, 5.612017, 5.612091, 5.612052, 5.612098, 5.611995, 5.611943, 
    5.611931, 5.611906, 5.611932, 5.61193, 5.611954, 5.611946, 5.612004, 
    5.611973, 5.612064, 5.612097, 5.612192, 5.612248, 5.612308, 5.612333, 
    5.61234, 5.612344 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  5.913039e-15, 5.911907e-15, 5.912122e-15, 5.911222e-15, 5.911713e-15, 
    5.91113e-15, 5.9128e-15, 5.911871e-15, 5.912458e-15, 5.912924e-15, 
    5.909506e-15, 5.911179e-15, 5.907683e-15, 5.908762e-15, 5.906028e-15, 
    5.907863e-15, 5.905655e-15, 5.906059e-15, 5.904791e-15, 5.905153e-15, 
    5.903578e-15, 5.904624e-15, 5.90273e-15, 5.903816e-15, 5.903654e-15, 
    5.904662e-15, 5.910821e-15, 5.90972e-15, 5.910892e-15, 5.910734e-15, 
    5.9108e-15, 5.91171e-15, 5.912184e-15, 5.913111e-15, 5.912938e-15, 
    5.91225e-15, 5.910662e-15, 5.911186e-15, 5.909824e-15, 5.909854e-15, 
    5.908355e-15, 5.909031e-15, 5.9065e-15, 5.907214e-15, 5.905137e-15, 
    5.905662e-15, 5.905166e-15, 5.905313e-15, 5.905163e-15, 5.905932e-15, 
    5.905604e-15, 5.906273e-15, 5.908909e-15, 5.90814e-15, 5.910446e-15, 
    5.911869e-15, 5.912763e-15, 5.913414e-15, 5.913323e-15, 5.913151e-15, 
    5.912246e-15, 5.911378e-15, 5.910723e-15, 5.910289e-15, 5.909859e-15, 
    5.908613e-15, 5.907908e-15, 5.906366e-15, 5.906626e-15, 5.906172e-15, 
    5.905713e-15, 5.904968e-15, 5.905088e-15, 5.904764e-15, 5.906171e-15, 
    5.905242e-15, 5.906779e-15, 5.90636e-15, 5.909814e-15, 5.911041e-15, 
    5.911626e-15, 5.912083e-15, 5.913253e-15, 5.912449e-15, 5.912768e-15, 
    5.911995e-15, 5.911515e-15, 5.911749e-15, 5.910277e-15, 5.910852e-15, 
    5.907866e-15, 5.90915e-15, 5.905767e-15, 5.906571e-15, 5.905571e-15, 
    5.906077e-15, 5.905216e-15, 5.905991e-15, 5.904637e-15, 5.904351e-15, 
    5.904549e-15, 5.903768e-15, 5.906036e-15, 5.905172e-15, 5.911759e-15, 
    5.911721e-15, 5.911537e-15, 5.91235e-15, 5.912395e-15, 5.913119e-15, 
    5.912468e-15, 5.912197e-15, 5.911481e-15, 5.911071e-15, 5.910677e-15, 
    5.909811e-15, 5.908856e-15, 5.907503e-15, 5.90652e-15, 5.905866e-15, 
    5.906262e-15, 5.905913e-15, 5.906306e-15, 5.906487e-15, 5.904463e-15, 
    5.905605e-15, 5.90388e-15, 5.903973e-15, 5.904759e-15, 5.903962e-15, 
    5.911694e-15, 5.911913e-15, 5.912701e-15, 5.912084e-15, 5.913197e-15, 
    5.912583e-15, 5.912235e-15, 5.910856e-15, 5.910535e-15, 5.910261e-15, 
    5.909704e-15, 5.908997e-15, 5.907763e-15, 5.90668e-15, 5.905684e-15, 
    5.905755e-15, 5.90573e-15, 5.905515e-15, 5.906058e-15, 5.905426e-15, 
    5.905327e-15, 5.905596e-15, 5.903986e-15, 5.904444e-15, 5.903975e-15, 
    5.904272e-15, 5.91184e-15, 5.911467e-15, 5.91167e-15, 5.911292e-15, 
    5.911564e-15, 5.910378e-15, 5.910023e-15, 5.908344e-15, 5.909015e-15, 
    5.907928e-15, 5.908899e-15, 5.908731e-15, 5.907923e-15, 5.908842e-15, 
    5.906755e-15, 5.908195e-15, 5.905507e-15, 5.906972e-15, 5.905417e-15, 
    5.905688e-15, 5.905232e-15, 5.904832e-15, 5.904316e-15, 5.903387e-15, 
    5.903599e-15, 5.902811e-15, 5.910904e-15, 5.910427e-15, 5.910456e-15, 
    5.909948e-15, 5.909576e-15, 5.908752e-15, 5.907449e-15, 5.907934e-15, 
    5.907029e-15, 5.906852e-15, 5.90822e-15, 5.907392e-15, 5.910098e-15, 
    5.909674e-15, 5.909917e-15, 5.910874e-15, 5.907841e-15, 5.909404e-15, 
    5.906506e-15, 5.907349e-15, 5.904891e-15, 5.906125e-15, 5.903719e-15, 
    5.902728e-15, 5.901736e-15, 5.90065e-15, 5.910153e-15, 5.910478e-15, 
    5.909884e-15, 5.909087e-15, 5.90831e-15, 5.907301e-15, 5.90719e-15, 
    5.907004e-15, 5.906508e-15, 5.906098e-15, 5.906959e-15, 5.905994e-15, 
    5.909603e-15, 5.907699e-15, 5.910613e-15, 5.909753e-15, 5.909128e-15, 
    5.909388e-15, 5.907986e-15, 5.907661e-15, 5.906345e-15, 5.907018e-15, 
    5.902984e-15, 5.904767e-15, 5.89978e-15, 5.901178e-15, 5.910595e-15, 
    5.910147e-15, 5.908612e-15, 5.90934e-15, 5.907226e-15, 5.906712e-15, 
    5.906282e-15, 5.905757e-15, 5.90569e-15, 5.905378e-15, 5.905892e-15, 
    5.905393e-15, 5.907298e-15, 5.906443e-15, 5.908771e-15, 5.908212e-15, 
    5.908465e-15, 5.908752e-15, 5.907867e-15, 5.906949e-15, 5.906908e-15, 
    5.906616e-15, 5.905837e-15, 5.907216e-15, 5.902795e-15, 5.905558e-15, 
    5.909661e-15, 5.908831e-15, 5.908685e-15, 5.909012e-15, 5.906765e-15, 
    5.90758e-15, 5.905382e-15, 5.905971e-15, 5.905001e-15, 5.905484e-15, 
    5.905557e-15, 5.906173e-15, 5.906564e-15, 5.907547e-15, 5.908342e-15, 
    5.908962e-15, 5.908816e-15, 5.908135e-15, 5.906888e-15, 5.905694e-15, 
    5.905958e-15, 5.905075e-15, 5.907379e-15, 5.906423e-15, 5.9068e-15, 
    5.905814e-15, 5.907951e-15, 5.906196e-15, 5.908409e-15, 5.90821e-15, 
    5.907597e-15, 5.906373e-15, 5.90607e-15, 5.905786e-15, 5.905957e-15, 
    5.906852e-15, 5.906989e-15, 5.907606e-15, 5.907788e-15, 5.908252e-15, 
    5.908646e-15, 5.908291e-15, 5.907923e-15, 5.906843e-15, 5.905882e-15, 
    5.90483e-15, 5.904564e-15, 5.903392e-15, 5.904376e-15, 5.902783e-15, 
    5.904181e-15, 5.901741e-15, 5.906062e-15, 5.90418e-15, 5.907561e-15, 
    5.907191e-15, 5.906543e-15, 5.905018e-15, 5.905818e-15, 5.904872e-15, 
    5.906993e-15, 5.908122e-15, 5.908388e-15, 5.908928e-15, 5.908375e-15, 
    5.908419e-15, 5.907892e-15, 5.90806e-15, 5.906807e-15, 5.907479e-15, 
    5.905564e-15, 5.904874e-15, 5.902901e-15, 5.901709e-15, 5.900464e-15, 
    5.899926e-15, 5.899761e-15, 5.899693e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  7.136423, 7.162951, 7.15779, 7.179227, 7.167332, 7.181376, 7.141799, 
    7.164002, 7.149824, 7.138813, 7.220966, 7.180186, 7.263556, 7.237401, 
    7.303249, 7.259477, 7.312101, 7.301992, 7.332471, 7.32373, 7.362805, 
    7.336509, 7.383138, 7.356524, 7.360679, 7.335641, 7.188386, 7.215877, 
    7.186758, 7.190673, 7.188918, 7.167575, 7.156833, 7.134405, 7.138474, 
    7.154952, 7.192434, 7.179698, 7.211846, 7.211119, 7.247035, 7.230824, 
    7.2914, 7.274148, 7.324095, 7.311508, 7.323502, 7.319864, 7.323549, 
    7.305096, 7.312997, 7.296778, 7.233856, 7.252303, 7.197389, 7.164516, 
    7.14277, 7.127365, 7.129541, 7.133689, 7.155048, 7.175185, 7.190559, 
    7.200856, 7.211015, 7.241811, 7.258172, 7.294888, 7.288259, 7.299497, 
    7.310256, 7.328338, 7.325361, 7.333334, 7.299206, 7.321871, 7.284483, 
    7.294693, 7.213749, 7.183134, 7.170127, 7.158781, 7.131214, 7.15024, 
    7.142734, 7.160608, 7.171979, 7.166355, 7.201138, 7.187598, 7.259142, 
    7.228258, 7.309001, 7.28962, 7.313653, 7.301383, 7.322415, 7.303485, 
    7.336306, 7.343464, 7.338571, 7.357391, 7.302436, 7.323499, 7.166196, 
    7.167113, 7.171389, 7.152606, 7.151459, 7.134292, 7.149569, 7.15608, 
    7.172642, 7.182447, 7.19178, 7.212336, 7.235343, 7.267618, 7.290874, 
    7.306494, 7.296916, 7.305371, 7.295918, 7.291492, 7.340779, 7.313069, 
    7.354682, 7.352376, 7.333523, 7.352635, 7.167757, 7.16248, 7.144175, 
    7.158497, 7.132424, 7.147006, 7.155399, 7.187874, 7.195032, 7.201665, 
    7.214788, 7.231653, 7.26131, 7.287192, 7.310884, 7.309146, 7.309758, 
    7.315055, 7.301935, 7.317211, 7.319775, 7.313069, 7.352067, 7.340909, 
    7.352326, 7.345061, 7.164196, 7.173079, 7.168278, 7.177308, 7.170943, 
    7.199273, 7.207784, 7.247724, 7.231319, 7.257449, 7.233972, 7.238126, 
    7.258291, 7.235241, 7.285758, 7.25147, 7.315261, 7.280907, 7.317418, 
    7.310781, 7.321774, 7.331627, 7.344043, 7.366986, 7.36167, 7.380894, 
    7.186343, 7.197893, 7.196881, 7.208986, 7.217949, 7.237411, 7.268704, 
    7.256926, 7.278565, 7.282912, 7.250045, 7.270208, 7.205636, 7.216032, 
    7.209844, 7.18725, 7.259631, 7.22241, 7.291258, 7.271014, 7.330221, 
    7.300724, 7.358743, 7.383641, 7.407158, 7.434684, 7.204209, 7.196353, 
    7.210429, 7.229929, 7.248076, 7.272246, 7.274726, 7.279259, 7.291019, 
    7.300916, 7.280688, 7.303399, 7.218434, 7.262871, 7.193379, 7.214242, 
    7.228781, 7.222406, 7.255582, 7.263416, 7.295313, 7.278815, 7.377485, 
    7.333702, 7.455713, 7.421457, 7.193608, 7.204184, 7.24108, 7.223507, 
    7.273865, 7.286296, 7.29642, 7.309367, 7.31077, 7.318451, 7.305866, 
    7.317956, 7.272298, 7.292675, 7.236862, 7.250414, 7.244179, 7.237341, 
    7.258461, 7.281004, 7.281496, 7.288733, 7.309144, 7.27407, 7.383134, 
    7.315614, 7.21573, 7.23615, 7.239081, 7.231161, 7.285049, 7.265489, 
    7.318265, 7.303975, 7.327403, 7.315753, 7.31404, 7.299103, 7.289813, 
    7.266383, 7.247362, 7.232311, 7.235809, 7.25235, 7.282387, 7.310893, 
    7.30464, 7.325621, 7.270205, 7.293397, 7.284424, 7.307842, 7.256611, 
    7.300193, 7.245499, 7.250284, 7.2651, 7.294967, 7.3016, 7.308671, 
    7.304309, 7.283153, 7.279695, 7.264742, 7.260613, 7.249243, 7.239835, 
    7.248428, 7.257459, 7.283165, 7.306383, 7.331766, 7.337992, 7.367734, 
    7.343504, 7.38351, 7.349469, 7.408483, 7.302738, 7.348486, 7.265779, 
    7.274658, 7.290726, 7.327703, 7.307732, 7.331097, 7.27956, 7.252917, 
    7.246047, 7.233223, 7.24634, 7.245273, 7.257839, 7.253799, 7.284019, 
    7.267776, 7.313994, 7.330914, 7.378874, 7.408389, 7.43854, 7.451876, 
    7.455939, 7.457638 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002557226, 0.0002556717, 0.0002556814, 0.0002556408, 0.0002556629, 
    0.0002556367, 0.0002557119, 0.00025567, 0.0002556965, 0.0002557175, 
    0.0002555634, 0.0002556389, 0.0002554815, 0.0002555301, 0.000255407, 
    0.0002554896, 0.0002553902, 0.0002554085, 0.0002553514, 0.0002553677, 
    0.0002552966, 0.0002553438, 0.0002552583, 0.0002553074, 0.0002553, 
    0.0002553455, 0.0002556228, 0.0002555731, 0.000255626, 0.0002556188, 
    0.0002556219, 0.0002556628, 0.0002556841, 0.0002557259, 0.0002557182, 
    0.0002556871, 0.0002556156, 0.0002556393, 0.0002555779, 0.0002555793, 
    0.0002555118, 0.0002555422, 0.0002554283, 0.0002554605, 0.000255367, 
    0.0002553906, 0.0002553682, 0.0002553749, 0.0002553681, 0.0002554027, 
    0.0002553879, 0.0002554181, 0.0002555367, 0.0002555021, 0.0002556059, 
    0.0002556699, 0.0002557102, 0.0002557395, 0.0002557354, 0.0002557277, 
    0.0002556869, 0.0002556479, 0.0002556184, 0.0002555989, 0.0002555795, 
    0.0002555233, 0.0002554916, 0.0002554223, 0.000255434, 0.0002554135, 
    0.0002553929, 0.0002553593, 0.0002553647, 0.0002553501, 0.0002554135, 
    0.0002553716, 0.0002554409, 0.000255422, 0.0002555773, 0.0002556327, 
    0.000255659, 0.0002556796, 0.0002557323, 0.0002556961, 0.0002557104, 
    0.0002556756, 0.000255654, 0.0002556646, 0.0002555983, 0.0002556242, 
    0.0002554898, 0.0002555476, 0.0002553953, 0.0002554315, 0.0002553865, 
    0.0002554093, 0.0002553705, 0.0002554054, 0.0002553444, 0.0002553315, 
    0.0002553404, 0.0002553052, 0.0002554075, 0.0002553685, 0.000255665, 
    0.0002556633, 0.000255655, 0.0002556916, 0.0002556937, 0.0002557263, 
    0.000255697, 0.0002556847, 0.0002556525, 0.0002556341, 0.0002556163, 
    0.0002555773, 0.0002555343, 0.0002554734, 0.0002554292, 0.0002553998, 
    0.0002554176, 0.0002554019, 0.0002554196, 0.0002554278, 0.0002553365, 
    0.000255388, 0.0002553103, 0.0002553145, 0.0002553499, 0.000255314, 
    0.0002556621, 0.000255672, 0.0002557074, 0.0002556797, 0.0002557298, 
    0.0002557021, 0.0002556864, 0.0002556243, 0.0002556099, 0.0002555976, 
    0.0002555725, 0.0002555407, 0.0002554852, 0.0002554364, 0.0002553916, 
    0.0002553948, 0.0002553937, 0.000255384, 0.0002554084, 0.0002553799, 
    0.0002553755, 0.0002553877, 0.000255315, 0.0002553357, 0.0002553145, 
    0.000255328, 0.0002556687, 0.0002556519, 0.000255661, 0.000255644, 
    0.0002556562, 0.0002556028, 0.0002555868, 0.0002555113, 0.0002555415, 
    0.0002554925, 0.0002555363, 0.0002555287, 0.0002554923, 0.0002555337, 
    0.0002554397, 0.0002555046, 0.0002553836, 0.0002554495, 0.0002553796, 
    0.0002553918, 0.0002553712, 0.0002553532, 0.00025533, 0.000255288, 
    0.0002552976, 0.000255262, 0.0002556266, 0.0002556051, 0.0002556064, 
    0.0002555835, 0.0002555667, 0.0002555297, 0.000255471, 0.0002554929, 
    0.0002554521, 0.0002554441, 0.0002555057, 0.0002554684, 0.0002555902, 
    0.0002555711, 0.0002555821, 0.0002556252, 0.0002554886, 0.000255559, 
    0.0002554286, 0.0002554665, 0.0002553558, 0.0002554114, 0.000255303, 
    0.0002552582, 0.0002552135, 0.0002551643, 0.0002555927, 0.0002556074, 
    0.0002555806, 0.0002555447, 0.0002555098, 0.0002554643, 0.0002554593, 
    0.000255451, 0.0002554287, 0.0002554103, 0.0002554489, 0.0002554056, 
    0.0002555679, 0.0002554822, 0.0002556134, 0.0002555746, 0.0002555466, 
    0.0002555583, 0.0002554952, 0.0002554806, 0.0002554213, 0.0002554516, 
    0.0002552698, 0.0002553502, 0.000255125, 0.0002551882, 0.0002556127, 
    0.0002555925, 0.0002555233, 0.0002555561, 0.000255461, 0.0002554379, 
    0.0002554186, 0.0002553949, 0.0002553919, 0.0002553778, 0.000255401, 
    0.0002553785, 0.0002554642, 0.0002554258, 0.0002555306, 0.0002555054, 
    0.0002555167, 0.0002555297, 0.0002554899, 0.0002554485, 0.0002554466, 
    0.0002554336, 0.0002553983, 0.0002554606, 0.0002552611, 0.0002553858, 
    0.0002555706, 0.0002555331, 0.0002555267, 0.0002555414, 0.0002554402, 
    0.0002554769, 0.000255378, 0.0002554045, 0.0002553608, 0.0002553826, 
    0.0002553859, 0.0002554136, 0.0002554312, 0.0002554754, 0.0002555112, 
    0.0002555391, 0.0002555326, 0.0002555019, 0.0002554457, 0.000255392, 
    0.0002554039, 0.0002553641, 0.0002554679, 0.0002554248, 0.0002554418, 
    0.0002553974, 0.0002554937, 0.0002554145, 0.0002555142, 0.0002555053, 
    0.0002554777, 0.0002554225, 0.000255409, 0.0002553962, 0.0002554039, 
    0.0002554441, 0.0002554503, 0.0002554781, 0.0002554863, 0.0002555072, 
    0.0002555249, 0.0002555089, 0.0002554923, 0.0002554437, 0.0002554005, 
    0.0002553531, 0.0002553411, 0.0002552881, 0.0002553325, 0.0002552606, 
    0.0002553237, 0.0002552136, 0.0002554086, 0.0002553237, 0.0002554761, 
    0.0002554594, 0.0002554303, 0.0002553615, 0.0002553976, 0.0002553549, 
    0.0002554505, 0.0002555013, 0.0002555133, 0.0002555376, 0.0002555127, 
    0.0002555147, 0.000255491, 0.0002554985, 0.0002554421, 0.0002554724, 
    0.0002553862, 0.000255355, 0.0002552661, 0.0002552122, 0.000255156, 
    0.0002551317, 0.0002551242, 0.0002551211 ;

 W_SCALAR =
  0.6254858, 0.6271458, 0.6268232, 0.628161, 0.6274189, 0.6282948, 0.6258224, 
    0.6272117, 0.6263249, 0.6256352, 0.6307536, 0.6282206, 0.6333788, 
    0.6317673, 0.6358114, 0.6331283, 0.6363517, 0.6357339, 0.637592, 
    0.6370599, 0.6394339, 0.6378374, 0.6406623, 0.6390527, 0.6393047, 
    0.6377848, 0.6287306, 0.6304386, 0.6286293, 0.6288731, 0.6287637, 
    0.6274344, 0.6267641, 0.6253587, 0.6256139, 0.626646, 0.6289826, 
    0.6281898, 0.6301867, 0.6301416, 0.6323614, 0.631361, 0.6350861, 
    0.6340284, 0.6370822, 0.6363149, 0.6370462, 0.6368244, 0.637049, 
    0.6359236, 0.6364059, 0.635415, 0.6315484, 0.6326861, 0.6292902, 
    0.6272444, 0.6258834, 0.6249169, 0.6250536, 0.6253141, 0.6266521, 
    0.6279086, 0.6288654, 0.6295052, 0.6301351, 0.6320406, 0.6330476, 
    0.6352999, 0.6348936, 0.6355817, 0.6362385, 0.6373407, 0.6371593, 
    0.6376447, 0.6355634, 0.6369471, 0.6346622, 0.6352875, 0.630307, 
    0.6284037, 0.6275944, 0.6268852, 0.6251587, 0.6263512, 0.6258813, 
    0.626999, 0.6277088, 0.6273578, 0.6295226, 0.6286814, 0.6331073, 
    0.6312028, 0.6361619, 0.634977, 0.6364458, 0.6356965, 0.6369801, 
    0.6358249, 0.6378253, 0.6382605, 0.6379631, 0.6391048, 0.6357608, 
    0.6370462, 0.6273479, 0.6274052, 0.6276719, 0.6264992, 0.6264275, 
    0.6253517, 0.6263089, 0.6267164, 0.6277499, 0.628361, 0.6289415, 
    0.6302172, 0.6316405, 0.633628, 0.6350538, 0.6360087, 0.6354232, 
    0.6359402, 0.6353623, 0.6350914, 0.6380975, 0.6364105, 0.6389407, 
    0.6388008, 0.6376563, 0.6388165, 0.6274454, 0.6271158, 0.6259713, 
    0.6268671, 0.6252345, 0.6261487, 0.6266741, 0.6286991, 0.6291435, 
    0.6295556, 0.630369, 0.6314122, 0.6332403, 0.6348286, 0.6362767, 
    0.6361706, 0.636208, 0.6365314, 0.6357303, 0.6366628, 0.6368193, 
    0.6364102, 0.638782, 0.6381049, 0.6387978, 0.6383569, 0.627223, 
    0.6277773, 0.6274778, 0.628041, 0.6276444, 0.6294076, 0.6299358, 
    0.6324044, 0.6313917, 0.6330029, 0.6315554, 0.631812, 0.6330557, 
    0.6316336, 0.6347412, 0.6326354, 0.6365439, 0.6344444, 0.6366754, 
    0.6362705, 0.6369407, 0.6375408, 0.6382952, 0.6396862, 0.6393642, 
    0.6405264, 0.6286033, 0.6293216, 0.6292583, 0.6300095, 0.6305649, 
    0.6317676, 0.6336944, 0.6329702, 0.6342993, 0.6345661, 0.6325465, 
    0.633787, 0.629802, 0.6304468, 0.6300629, 0.6286601, 0.6331373, 
    0.6308416, 0.6350774, 0.6338362, 0.6374553, 0.6356568, 0.639187, 
    0.6406932, 0.6421086, 0.6437612, 0.6297134, 0.6292255, 0.6300988, 
    0.6313064, 0.6324254, 0.6339119, 0.6340638, 0.6343421, 0.6350625, 
    0.6356679, 0.6344302, 0.6358196, 0.6305966, 0.6333363, 0.6290411, 
    0.6303361, 0.6312352, 0.6308407, 0.6328873, 0.6333693, 0.6353258, 
    0.6343147, 0.6403218, 0.6376677, 0.6450174, 0.6429682, 0.629055, 
    0.6297116, 0.6319945, 0.6309088, 0.634011, 0.6347735, 0.6353929, 
    0.6361845, 0.6362698, 0.6367385, 0.6359704, 0.6367081, 0.6339151, 
    0.635164, 0.6317336, 0.6325694, 0.632185, 0.6317632, 0.6330645, 
    0.6344497, 0.6344791, 0.634923, 0.6361732, 0.6340235, 0.6406643, 
    0.6365677, 0.6304272, 0.6316907, 0.6318708, 0.6313816, 0.6346971, 
    0.6334968, 0.636727, 0.6358548, 0.6372836, 0.6365739, 0.6364694, 
    0.6355571, 0.6349888, 0.6335519, 0.6323815, 0.6314526, 0.6316686, 
    0.6326888, 0.6345344, 0.6362776, 0.635896, 0.6371751, 0.6337863, 
    0.6352085, 0.6346591, 0.6360911, 0.632951, 0.6356261, 0.6322663, 
    0.6325612, 0.633473, 0.635305, 0.6357097, 0.636142, 0.6358752, 0.6345811, 
    0.6343689, 0.6334507, 0.6331972, 0.632497, 0.6319171, 0.632447, 
    0.6330033, 0.6345816, 0.6360024, 0.6375494, 0.6379277, 0.6397327, 
    0.6382638, 0.6406871, 0.6386275, 0.6421903, 0.6357806, 0.6385665, 
    0.6335143, 0.6340595, 0.6350453, 0.6373029, 0.6360844, 0.6375092, 
    0.6343606, 0.6327241, 0.6323001, 0.6315091, 0.6323182, 0.6322524, 
    0.6330262, 0.6327776, 0.634634, 0.6336371, 0.6364668, 0.6374979, 
    0.6404048, 0.6421834, 0.6439909, 0.6447881, 0.6450306, 0.645132,
  0.5466921, 0.5487348, 0.5483378, 0.5499842, 0.549071, 0.5501489, 0.5471063, 
    0.5488159, 0.5477247, 0.546876, 0.5531755, 0.5500576, 0.5564078, 
    0.5544235, 0.5594037, 0.5560993, 0.5600693, 0.5593082, 0.5615971, 
    0.5609417, 0.5638664, 0.5618995, 0.5653803, 0.5633968, 0.5637074, 
    0.5618346, 0.5506853, 0.5527877, 0.5505607, 0.5508606, 0.550726, 0.54909, 
    0.5482651, 0.5465358, 0.5468498, 0.5481198, 0.5509955, 0.5500197, 
    0.5524776, 0.5524221, 0.5551549, 0.5539232, 0.5585103, 0.5572077, 
    0.5609691, 0.5600239, 0.5609247, 0.5606515, 0.5609282, 0.5595419, 
    0.560136, 0.5589155, 0.554154, 0.5555547, 0.5513741, 0.5488562, 
    0.5471814, 0.5459922, 0.5461604, 0.546481, 0.5481272, 0.5496736, 
    0.5508513, 0.5516387, 0.5524141, 0.5547601, 0.556, 0.5587737, 0.5582733, 
    0.5591208, 0.5599298, 0.5612875, 0.5610641, 0.5616621, 0.5590983, 
    0.5608027, 0.5579882, 0.5587584, 0.5526257, 0.550283, 0.549287, 
    0.5484142, 0.5462897, 0.5477571, 0.5471787, 0.5485542, 0.5494277, 
    0.5489957, 0.5516602, 0.5506248, 0.5560735, 0.5537285, 0.5598355, 
    0.558376, 0.5601851, 0.5592622, 0.5608433, 0.5594203, 0.5618845, 
    0.5624207, 0.5620543, 0.5634611, 0.5593414, 0.5609248, 0.5489836, 
    0.5490541, 0.5493823, 0.5479392, 0.5478508, 0.5465272, 0.547705, 
    0.5482064, 0.5494783, 0.5502304, 0.550945, 0.5525152, 0.5542674, 
    0.5567147, 0.5584706, 0.5596468, 0.5589256, 0.5595623, 0.5588506, 
    0.5585169, 0.5622199, 0.5601416, 0.5632588, 0.5630865, 0.5616763, 
    0.5631058, 0.5491036, 0.548698, 0.5472896, 0.5483919, 0.546383, 
    0.5475078, 0.5481544, 0.5506466, 0.5511935, 0.5517008, 0.5527021, 
    0.5539863, 0.5562372, 0.5581932, 0.5599768, 0.5598462, 0.5598922, 
    0.5602905, 0.5593038, 0.5604525, 0.5606452, 0.5601413, 0.5630633, 
    0.562229, 0.5630828, 0.5625396, 0.5488299, 0.5495121, 0.5491435, 
    0.5498366, 0.5493484, 0.5515186, 0.5521688, 0.555208, 0.5539611, 
    0.5559449, 0.5541627, 0.5544786, 0.5560099, 0.5542589, 0.5580856, 
    0.5554924, 0.560306, 0.55772, 0.560468, 0.5599691, 0.5607948, 0.5615341, 
    0.5624635, 0.5641775, 0.5637807, 0.5652128, 0.5505286, 0.5514128, 
    0.5513348, 0.5522596, 0.5529432, 0.5544239, 0.5567964, 0.5559046, 
    0.5575414, 0.5578699, 0.5553829, 0.5569104, 0.5520042, 0.5527979, 
    0.5523252, 0.5505985, 0.5561103, 0.5532838, 0.5584996, 0.556971, 
    0.5614287, 0.5592133, 0.5635623, 0.5654185, 0.5671629, 0.5692, 0.551895, 
    0.5512944, 0.5523694, 0.553856, 0.5552338, 0.5570642, 0.5572513, 
    0.5575941, 0.5584813, 0.559227, 0.5577025, 0.5594139, 0.5529822, 
    0.5563554, 0.5510675, 0.5526615, 0.5537683, 0.5532828, 0.5558026, 
    0.556396, 0.5588056, 0.5575603, 0.5649607, 0.5616904, 0.5707489, 
    0.5682224, 0.5510846, 0.5518928, 0.5547032, 0.5533665, 0.5571863, 
    0.5581254, 0.5588883, 0.5598632, 0.5599684, 0.5605457, 0.5595995, 
    0.5605083, 0.5570682, 0.5586063, 0.554382, 0.5554112, 0.5549378, 
    0.5544184, 0.5560208, 0.5577266, 0.5577627, 0.5583094, 0.5598494, 
    0.5572017, 0.5653827, 0.5603353, 0.5527738, 0.5543292, 0.5545509, 
    0.5539487, 0.5580313, 0.5565531, 0.5605316, 0.5594572, 0.5612172, 
    0.5603428, 0.5602142, 0.5590904, 0.5583905, 0.5566209, 0.5551798, 
    0.554036, 0.554302, 0.5555581, 0.5578308, 0.5599779, 0.5595079, 
    0.5610835, 0.5569096, 0.5586611, 0.5579844, 0.5597483, 0.5558809, 
    0.5591754, 0.5550379, 0.555401, 0.5565237, 0.55878, 0.5592784, 0.5598109, 
    0.5594823, 0.5578884, 0.5576271, 0.5564964, 0.5561842, 0.555322, 
    0.5546079, 0.5552604, 0.5559454, 0.557889, 0.5596389, 0.5615447, 
    0.5620106, 0.5642347, 0.5624248, 0.5654109, 0.5628729, 0.5672635, 
    0.5593658, 0.5627978, 0.5565747, 0.5572461, 0.5584601, 0.5612409, 
    0.5597399, 0.5614951, 0.5576168, 0.5556016, 0.5550796, 0.5541056, 
    0.5551018, 0.5550208, 0.5559736, 0.5556675, 0.5579535, 0.5567259, 
    0.560211, 0.5614812, 0.5650629, 0.5672551, 0.5694832, 0.5704661, 
    0.5707651, 0.5708901,
  0.514178, 0.5164279, 0.5159906, 0.5178043, 0.5167983, 0.5179858, 0.5146342, 
    0.5165172, 0.5153152, 0.5143805, 0.5213212, 0.5178852, 0.5248849, 
    0.522697, 0.5281896, 0.5245447, 0.5289239, 0.5280843, 0.5306099, 
    0.5298866, 0.533115, 0.5309437, 0.5347865, 0.5325965, 0.5329393, 
    0.5308721, 0.5185768, 0.5208938, 0.5184395, 0.51877, 0.5186217, 
    0.5168191, 0.5159105, 0.5140058, 0.5143517, 0.5157505, 0.5189186, 
    0.5178434, 0.520552, 0.5204908, 0.5235035, 0.5221456, 0.527204, 
    0.5257671, 0.5299168, 0.5288739, 0.5298679, 0.5295665, 0.5298718, 
    0.528342, 0.5289976, 0.527651, 0.5224, 0.5239443, 0.5193359, 0.5165616, 
    0.5147169, 0.5134073, 0.5135924, 0.5139455, 0.5157586, 0.5174621, 
    0.5187597, 0.5196274, 0.5204821, 0.5230681, 0.5244353, 0.5274945, 
    0.5269425, 0.5278774, 0.5287701, 0.5302683, 0.5300217, 0.5306817, 
    0.5278527, 0.5297332, 0.526628, 0.5274777, 0.5207152, 0.5181335, 
    0.5170361, 0.5160747, 0.5137348, 0.5153509, 0.5147139, 0.5162289, 
    0.5171912, 0.5167153, 0.5196511, 0.5185102, 0.5245163, 0.5219308, 
    0.528666, 0.5270558, 0.5290517, 0.5280334, 0.5297781, 0.528208, 
    0.5309271, 0.531519, 0.5311146, 0.5326674, 0.5281209, 0.5298679, 
    0.516702, 0.5167796, 0.5171412, 0.5155516, 0.5154542, 0.5139964, 
    0.5152935, 0.5158458, 0.517247, 0.5180755, 0.518863, 0.5205934, 0.522525, 
    0.5252234, 0.5271602, 0.5284578, 0.5276622, 0.5283646, 0.5275794, 
    0.5272112, 0.5312973, 0.5290037, 0.5324441, 0.5322538, 0.5306973, 
    0.5322753, 0.5168341, 0.5163874, 0.514836, 0.5160502, 0.5138376, 
    0.5150764, 0.5157886, 0.5185342, 0.5191368, 0.5196959, 0.5207994, 
    0.5222151, 0.5246968, 0.5268542, 0.5288219, 0.5286778, 0.5287285, 
    0.5291681, 0.5280794, 0.5293468, 0.5295594, 0.5290034, 0.5322284, 
    0.5313074, 0.5322498, 0.5316502, 0.5165326, 0.5172842, 0.5168781, 
    0.5176417, 0.5171039, 0.5194951, 0.5202116, 0.523562, 0.5221872, 
    0.5243745, 0.5224094, 0.5227578, 0.5244462, 0.5225156, 0.5267354, 
    0.5238755, 0.5291851, 0.5263322, 0.5293638, 0.5288135, 0.5297246, 
    0.5305404, 0.5315663, 0.5334583, 0.5330203, 0.5346016, 0.5184042, 
    0.5193785, 0.5192925, 0.5203117, 0.5210652, 0.5226974, 0.5253136, 
    0.52433, 0.5261352, 0.5264975, 0.5237548, 0.5254393, 0.5200302, 0.520905, 
    0.520384, 0.5184811, 0.5245569, 0.5214406, 0.5271922, 0.525506, 
    0.5304241, 0.5279796, 0.5327791, 0.5348286, 0.5367553, 0.5390058, 
    0.5199099, 0.5192481, 0.5204328, 0.5220714, 0.5235904, 0.525609, 
    0.5258153, 0.5261933, 0.527172, 0.5279946, 0.5263129, 0.5282007, 
    0.5211082, 0.5248272, 0.518998, 0.5207548, 0.5219747, 0.5214395, 
    0.5242175, 0.524872, 0.5275297, 0.5261561, 0.5343231, 0.5307129, 
    0.5407174, 0.5379257, 0.5190168, 0.5199075, 0.5230054, 0.5215318, 
    0.5257435, 0.5267794, 0.5276209, 0.5286966, 0.5288126, 0.5294496, 
    0.5284056, 0.5294083, 0.5256132, 0.5273098, 0.5226513, 0.523786, 
    0.523264, 0.5226914, 0.5244582, 0.5263395, 0.5263794, 0.5269824, 
    0.5286813, 0.5257606, 0.5347891, 0.5292174, 0.5208784, 0.522593, 
    0.5228375, 0.5221736, 0.5266755, 0.5250452, 0.5294341, 0.5282486, 
    0.5301906, 0.5292258, 0.5290838, 0.527844, 0.5270718, 0.52512, 0.5235308, 
    0.5222698, 0.5225631, 0.5239481, 0.5264544, 0.5288232, 0.5283045, 
    0.5300431, 0.5254384, 0.5273703, 0.5266239, 0.5285698, 0.524304, 
    0.5279378, 0.5233744, 0.5237748, 0.5250128, 0.5275015, 0.5280514, 
    0.5286389, 0.5282763, 0.526518, 0.5262297, 0.5249827, 0.5246384, 
    0.5236876, 0.5229003, 0.5236197, 0.5243751, 0.5265186, 0.5284491, 
    0.530552, 0.5310664, 0.5335215, 0.5315234, 0.5348202, 0.5320181, 
    0.5368664, 0.5281478, 0.5319352, 0.5250691, 0.5258095, 0.5271487, 
    0.5302169, 0.5285606, 0.5304974, 0.5262184, 0.5239959, 0.5234203, 
    0.5223466, 0.5234449, 0.5233555, 0.5244061, 0.5240686, 0.5265898, 
    0.5252358, 0.5290803, 0.530482, 0.534436, 0.5368571, 0.5393187, 
    0.5404049, 0.5407354, 0.5408735,
  0.507082, 0.5094725, 0.5090078, 0.5109357, 0.5098662, 0.5111286, 0.5075666, 
    0.5095676, 0.5082902, 0.507297, 0.5146761, 0.5110217, 0.5184693, 
    0.5161401, 0.5219896, 0.5181071, 0.5227721, 0.5218773, 0.5245695, 
    0.5237983, 0.5272413, 0.5249254, 0.529025, 0.5266882, 0.5270539, 
    0.5248491, 0.511757, 0.5142213, 0.511611, 0.5119625, 0.5118047, 
    0.5098884, 0.5089227, 0.5068991, 0.5072665, 0.5087526, 0.5121205, 
    0.5109772, 0.5138577, 0.5137927, 0.5169985, 0.5155532, 0.5209394, 
    0.5194088, 0.5238305, 0.5227188, 0.5237784, 0.5234571, 0.5237826, 
    0.522152, 0.5228506, 0.5214157, 0.515824, 0.5174678, 0.5125642, 
    0.5096147, 0.5076544, 0.5062633, 0.50646, 0.5068349, 0.5087613, 
    0.5105719, 0.5119515, 0.5128742, 0.5137833, 0.516535, 0.5179905, 
    0.5212489, 0.5206608, 0.5216569, 0.5226082, 0.5242053, 0.5239424, 
    0.524646, 0.5216305, 0.5236348, 0.5203258, 0.521231, 0.5140313, 
    0.5112857, 0.5101191, 0.5090972, 0.5066112, 0.5083281, 0.5076513, 
    0.5092611, 0.5102839, 0.509778, 0.5128995, 0.5116861, 0.5180768, 
    0.5153247, 0.5224972, 0.5207815, 0.5229084, 0.5218231, 0.5236827, 
    0.5220091, 0.5249078, 0.5255389, 0.5251076, 0.5267639, 0.5219163, 
    0.5237784, 0.5097639, 0.5098464, 0.5102307, 0.5085413, 0.5084379, 
    0.506889, 0.5082671, 0.508854, 0.5103431, 0.511224, 0.5120613, 0.5139018, 
    0.515957, 0.5188297, 0.5208927, 0.5222753, 0.5214275, 0.522176, 
    0.5213393, 0.520947, 0.5253025, 0.5228572, 0.5265257, 0.5263227, 
    0.5246627, 0.5263456, 0.5099043, 0.5094295, 0.507781, 0.5090712, 
    0.5067204, 0.5080364, 0.5087931, 0.5117117, 0.5123526, 0.5129471, 
    0.5141209, 0.5156272, 0.518269, 0.5205667, 0.5226635, 0.5225099, 
    0.5225639, 0.5230324, 0.5218721, 0.5232229, 0.5234496, 0.5228568, 
    0.5262955, 0.5253133, 0.5263184, 0.5256788, 0.5095838, 0.5103827, 
    0.5099511, 0.5107628, 0.510191, 0.5127335, 0.5134957, 0.5170608, 
    0.5155976, 0.5179259, 0.5158341, 0.5162048, 0.5180022, 0.515947, 
    0.5204402, 0.5173946, 0.5230506, 0.5200107, 0.523241, 0.5226544, 
    0.5236256, 0.5244954, 0.5255893, 0.5276076, 0.5271403, 0.5288277, 
    0.5115735, 0.5126095, 0.5125181, 0.5136021, 0.5144036, 0.5161406, 
    0.5189258, 0.5178785, 0.5198008, 0.5201868, 0.5172661, 0.5190596, 
    0.5133026, 0.5142332, 0.513679, 0.5116553, 0.5181201, 0.5148031, 
    0.5209268, 0.5191307, 0.5243714, 0.5217658, 0.526883, 0.52907, 0.5311269, 
    0.5335307, 0.5131747, 0.5124708, 0.5137309, 0.5154743, 0.5170911, 
    0.5192403, 0.5194601, 0.5198627, 0.5209053, 0.5217817, 0.5199901, 
    0.5220014, 0.5144494, 0.5184078, 0.5122048, 0.5140734, 0.5153715, 
    0.5148019, 0.5177587, 0.5184555, 0.5212864, 0.519823, 0.5285304, 
    0.5246793, 0.53536, 0.5323769, 0.5122249, 0.5131721, 0.5164683, 
    0.5149002, 0.5193837, 0.520487, 0.5213836, 0.5225298, 0.5226535, 
    0.5233325, 0.5222198, 0.5232885, 0.5192449, 0.5210521, 0.5160915, 
    0.5172992, 0.5167436, 0.5161342, 0.5180149, 0.5200184, 0.5200609, 
    0.5207033, 0.5225136, 0.5194018, 0.5290278, 0.523085, 0.514205, 
    0.5160294, 0.5162897, 0.515583, 0.5203764, 0.5186399, 0.523316, 
    0.5220524, 0.5241225, 0.5230939, 0.5229426, 0.5216213, 0.5207986, 
    0.5187196, 0.5170276, 0.5156855, 0.5159976, 0.5174718, 0.5201409, 
    0.5226648, 0.522112, 0.5239652, 0.5190587, 0.5211166, 0.5203214, 
    0.5223947, 0.5178507, 0.5217212, 0.5168612, 0.5172874, 0.5186055, 
    0.5212563, 0.5218423, 0.5224684, 0.522082, 0.5202085, 0.5199015, 
    0.5185734, 0.5182068, 0.5171946, 0.5163565, 0.5171223, 0.5179264, 
    0.5202093, 0.5222661, 0.5245078, 0.5250562, 0.5276751, 0.5255436, 
    0.529061, 0.5260713, 0.5312456, 0.521945, 0.5259828, 0.5186654, 
    0.5194539, 0.5208804, 0.5241504, 0.5223849, 0.5244495, 0.5198894, 
    0.5175228, 0.51691, 0.5157672, 0.5169361, 0.5168411, 0.5179595, 
    0.5176001, 0.520285, 0.5188429, 0.5229389, 0.5244331, 0.528651, 
    0.5312356, 0.5338652, 0.5350259, 0.5353791, 0.5355268,
  0.5310288, 0.5334982, 0.5330179, 0.5350106, 0.533905, 0.5352101, 0.5315292, 
    0.5335963, 0.5322765, 0.5312509, 0.5388809, 0.5350995, 0.5428115, 
    0.5403972, 0.5464646, 0.5424359, 0.5472774, 0.546348, 0.5491452, 
    0.5483436, 0.5519241, 0.5495152, 0.5537811, 0.5513485, 0.5517291, 
    0.5494357, 0.5358599, 0.53841, 0.535709, 0.5360725, 0.5359093, 0.5339279, 
    0.53293, 0.5308399, 0.5312192, 0.5327542, 0.5362359, 0.5350536, 
    0.5380336, 0.5379663, 0.5412867, 0.5397893, 0.5453742, 0.543786, 
    0.548377, 0.547222, 0.5483229, 0.547989, 0.5483272, 0.5466332, 0.5473589, 
    0.5458686, 0.5400698, 0.5417732, 0.536695, 0.533645, 0.5316199, 
    0.5301836, 0.5303866, 0.5307737, 0.5327632, 0.5346345, 0.5360612, 
    0.5370158, 0.5379566, 0.5408065, 0.5423151, 0.5456956, 0.5450851, 
    0.5461192, 0.5471071, 0.5487666, 0.5484933, 0.5492246, 0.5460917, 
    0.5481737, 0.5447374, 0.545677, 0.5382133, 0.5353725, 0.5341663, 
    0.5331103, 0.5305427, 0.5323157, 0.5316167, 0.5332797, 0.5343368, 
    0.5338139, 0.5370419, 0.5357866, 0.5424045, 0.5395526, 0.5469918, 
    0.5452104, 0.547419, 0.5462918, 0.5482234, 0.5464849, 0.5494968, 
    0.5501531, 0.5497046, 0.5514272, 0.5463886, 0.5483229, 0.5337992, 
    0.5338845, 0.5342818, 0.5325359, 0.5324291, 0.5308296, 0.5322527, 
    0.532859, 0.534398, 0.5353088, 0.5361747, 0.5380793, 0.5402075, 
    0.5431852, 0.5453258, 0.5467613, 0.545881, 0.5466582, 0.5457894, 
    0.5453822, 0.5499072, 0.5473658, 0.5511795, 0.5509683, 0.5492421, 
    0.5509921, 0.5339444, 0.5334537, 0.5317506, 0.5330834, 0.5306554, 
    0.5320144, 0.5327961, 0.5358131, 0.536476, 0.5370911, 0.5383061, 
    0.5398659, 0.5426038, 0.5449874, 0.5471645, 0.5470049, 0.5470611, 
    0.5475478, 0.5463426, 0.5477456, 0.5479812, 0.5473654, 0.55094, 
    0.5499184, 0.5509638, 0.5502986, 0.5336131, 0.5344389, 0.5339927, 
    0.5348319, 0.5342407, 0.5368702, 0.5376589, 0.5413513, 0.5398353, 
    0.542248, 0.5400802, 0.5404643, 0.5423271, 0.5401973, 0.5448561, 
    0.5416973, 0.5475667, 0.5444103, 0.5477645, 0.5471551, 0.5481641, 
    0.5490681, 0.5502055, 0.5523053, 0.551819, 0.5535756, 0.5356702, 
    0.5367419, 0.5366473, 0.537769, 0.5385988, 0.5403978, 0.5432849, 
    0.5421989, 0.5441927, 0.5445932, 0.5415641, 0.5434238, 0.5374591, 
    0.5384223, 0.5378487, 0.5357548, 0.5424494, 0.5390124, 0.5453612, 
    0.5434975, 0.5489392, 0.5462322, 0.5515513, 0.5538279, 0.555971, 
    0.5584781, 0.5373267, 0.5365984, 0.5379024, 0.5397075, 0.5413827, 
    0.5436112, 0.5438392, 0.5442569, 0.5453388, 0.5462488, 0.5443891, 
    0.546477, 0.5386461, 0.5427478, 0.5363232, 0.5382569, 0.539601, 
    0.5390112, 0.5420747, 0.5427972, 0.5457345, 0.5442157, 0.553266, 
    0.5492593, 0.5603875, 0.5572744, 0.536344, 0.5373241, 0.5407374, 
    0.5391129, 0.5437599, 0.5449046, 0.5458354, 0.5470257, 0.5471541, 
    0.5478596, 0.5467037, 0.5478138, 0.5436159, 0.5454913, 0.5403469, 
    0.5415984, 0.5410226, 0.5403911, 0.5423404, 0.5444184, 0.5444626, 
    0.5451292, 0.5470088, 0.5437787, 0.553784, 0.5476024, 0.5383931, 
    0.5402825, 0.5405522, 0.5398202, 0.5447899, 0.5429885, 0.5478423, 
    0.5465299, 0.5486805, 0.5476117, 0.5474545, 0.5460821, 0.5452281, 
    0.5430712, 0.5413169, 0.5399263, 0.5402496, 0.5417773, 0.5445455, 
    0.5471659, 0.5465918, 0.548517, 0.5434228, 0.5455582, 0.5447328, 
    0.5468853, 0.5421701, 0.5461859, 0.5411444, 0.5415861, 0.5429527, 
    0.5457033, 0.5463117, 0.5469618, 0.5465606, 0.5446157, 0.5442971, 
    0.5429195, 0.5425393, 0.54149, 0.5406215, 0.541415, 0.5422486, 0.5446165, 
    0.5467517, 0.549081, 0.5496511, 0.5523756, 0.550158, 0.5538185, 
    0.5507067, 0.5560948, 0.5464183, 0.5506147, 0.5430148, 0.5438328, 
    0.545313, 0.5487095, 0.5468752, 0.5490204, 0.5442846, 0.5418302, 
    0.541195, 0.5400109, 0.5412221, 0.5411236, 0.5422829, 0.5419103, 
    0.5446951, 0.5431989, 0.5474506, 0.5490034, 0.5533916, 0.5560843, 
    0.558827, 0.5600387, 0.5604075, 0.5605617,
  0.535215, 0.5380583, 0.537505, 0.5398022, 0.5385273, 0.5400323, 0.5357908, 
    0.5381714, 0.5366511, 0.5354705, 0.5442734, 0.5399048, 0.5488272, 
    0.5460286, 0.5530714, 0.5483914, 0.5540173, 0.5529358, 0.5561932, 
    0.555259, 0.5594366, 0.5566247, 0.5616078, 0.5587642, 0.5592087, 
    0.5565321, 0.5407823, 0.5437287, 0.5406081, 0.5410277, 0.5408393, 
    0.5385537, 0.5374036, 0.5349978, 0.5354341, 0.5372012, 0.5412164, 
    0.5398518, 0.5432935, 0.5432156, 0.5470591, 0.5453246, 0.5518034, 
    0.5499582, 0.555298, 0.5539528, 0.5552348, 0.5548459, 0.5552399, 
    0.5532677, 0.5541123, 0.5523782, 0.5456493, 0.5476229, 0.5417466, 
    0.5382276, 0.5358952, 0.5342429, 0.5344764, 0.5349216, 0.5372116, 
    0.5393683, 0.5410146, 0.5421172, 0.5432045, 0.5465026, 0.5482513, 
    0.552177, 0.5514672, 0.5526696, 0.5538191, 0.5557519, 0.5554335, 
    0.5562859, 0.5526377, 0.5550611, 0.5510632, 0.5521553, 0.5435013, 
    0.5402197, 0.5388285, 0.5376113, 0.5346559, 0.5366962, 0.5358915, 
    0.5378065, 0.539025, 0.5384222, 0.5421473, 0.5406978, 0.548355, 
    0.5450506, 0.5536849, 0.5516129, 0.5541821, 0.5528703, 0.555119, 
    0.553095, 0.5566033, 0.5573688, 0.5568456, 0.5588562, 0.5529829, 
    0.555235, 0.5384053, 0.5385036, 0.5389616, 0.5369498, 0.5368267, 
    0.5349858, 0.5366237, 0.5373218, 0.5390956, 0.5401462, 0.5411457, 
    0.5433463, 0.5458089, 0.5492609, 0.5517471, 0.5534167, 0.5523925, 
    0.5532967, 0.5522861, 0.5518126, 0.5570819, 0.5541202, 0.5585667, 
    0.5583202, 0.5563062, 0.558348, 0.5385727, 0.538007, 0.5360457, 
    0.5375804, 0.5347855, 0.5363493, 0.5372494, 0.5407283, 0.5414937, 
    0.5422042, 0.5436085, 0.5454133, 0.5485862, 0.5513538, 0.5538859, 
    0.5537002, 0.5537656, 0.5543321, 0.5529295, 0.5545625, 0.5548369, 
    0.5541198, 0.5582872, 0.557095, 0.558315, 0.5575385, 0.5381908, 
    0.5391428, 0.5386283, 0.539596, 0.5389143, 0.5419489, 0.5428603, 
    0.5471339, 0.5453779, 0.5481735, 0.5456614, 0.5461062, 0.5482653, 
    0.545797, 0.5512012, 0.5475349, 0.5543541, 0.5506833, 0.5545846, 
    0.553875, 0.55505, 0.5561034, 0.55743, 0.559882, 0.5593137, 0.5613673, 
    0.5405633, 0.5418007, 0.5416915, 0.5429876, 0.5439471, 0.5460292, 
    0.5493765, 0.5481166, 0.5504305, 0.5508956, 0.5473805, 0.5495377, 
    0.5426294, 0.543743, 0.5430797, 0.540661, 0.5484071, 0.5444255, 
    0.5517883, 0.5496233, 0.5559531, 0.552801, 0.559001, 0.5616626, 
    0.5641724, 0.5671141, 0.5424764, 0.541635, 0.5431418, 0.54523, 0.5471703, 
    0.5497553, 0.5500199, 0.550505, 0.5517622, 0.5528204, 0.5506586, 
    0.5530857, 0.5440018, 0.5487532, 0.5413172, 0.5435517, 0.5451067, 
    0.5444241, 0.5479726, 0.5488106, 0.5522222, 0.5504572, 0.5610052, 
    0.5563263, 0.5693585, 0.5657009, 0.5413412, 0.5424734, 0.5464225, 
    0.5445418, 0.5499279, 0.5512576, 0.5523396, 0.5537243, 0.5538738, 
    0.5546952, 0.5533496, 0.554642, 0.5497608, 0.5519395, 0.5459703, 
    0.5474204, 0.546753, 0.5460215, 0.5482807, 0.5506927, 0.5507439, 
    0.5515185, 0.5537046, 0.5499498, 0.5616112, 0.5543957, 0.5437092, 
    0.5458958, 0.546208, 0.5453604, 0.5511243, 0.5490325, 0.5546752, 
    0.5531473, 0.5556517, 0.5544065, 0.5542235, 0.5526266, 0.5516335, 
    0.5491284, 0.547094, 0.5454832, 0.5458576, 0.5476277, 0.5508403, 
    0.5538875, 0.5532194, 0.5554611, 0.5495365, 0.5520173, 0.5510579, 
    0.553561, 0.5480832, 0.5527471, 0.5468942, 0.5474061, 0.548991, 0.552186, 
    0.5528935, 0.5536501, 0.5531831, 0.5509219, 0.5505518, 0.5489524, 
    0.5485114, 0.5472946, 0.5462883, 0.5472078, 0.5481742, 0.5509228, 
    0.5534055, 0.5561185, 0.5567833, 0.5599641, 0.5573745, 0.5616516, 
    0.5580149, 0.5643175, 0.5530175, 0.5579075, 0.5490631, 0.5500126, 
    0.5517322, 0.5556855, 0.5535492, 0.5560478, 0.5505372, 0.547689, 
    0.5469528, 0.5455812, 0.5469842, 0.54687, 0.548214, 0.5477819, 0.5510141, 
    0.5492768, 0.554219, 0.5560279, 0.561152, 0.5643053, 0.567524, 0.5689483, 
    0.5693821, 0.5695636,
  0.5840928, 0.5875039, 0.586839, 0.5896026, 0.5880677, 0.5898799, 0.5847825, 
    0.5876399, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057424, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041865, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048915, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.58908, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046446, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052099, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834237, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924328, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.603953, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912229, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041979, 0.6106832, 0.6070316, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065955, 0.6072922, 0.6055682, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106994, 0.6122084, 0.6112477, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.592193, 0.593295, 0.598482, 0.5963469, 
    0.5997487, 0.5966913, 0.5972319, 0.5998606, 0.596856, 0.6034486, 
    0.5989705, 0.6073194, 0.6028146, 0.607603, 0.6067299, 0.6081761, 
    0.6094749, 0.6111134, 0.614151, 0.6134459, 0.6159967, 0.59052, 0.5920138, 
    0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 0.5996793, 
    0.6025052, 0.6030745, 0.5987824, 0.6014137, 0.5930157, 0.5943638, 
    0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 0.6015183, 
    0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 0.6231793, 
    0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 0.6016796, 
    0.6020032, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 0.5946774, 
    0.6004559, 0.5914299, 0.5941321, 0.5960177, 0.5951895, 0.5995038, 
    0.6005259, 0.6047001, 0.6025379, 0.6155463, 0.60975, 0.6260031, 
    0.6214069, 0.5914588, 0.592827, 0.5976165, 0.5953323, 0.6018906, 
    0.6035177, 0.604844, 0.6065448, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980185, 
    0.5971288, 0.5998793, 0.6028261, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073706, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039783, 0.6009138, 0.5984336, 0.5964749, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014124, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007462, 0.6046556, 0.6055239, 0.6064534, 
    0.6058796, 0.6031066, 0.6026536, 0.600699, 0.6001608, 0.5986778, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103142, 0.6142529, 0.6110448, 0.6163503, 0.6118369, 0.6196756, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040993, 0.6089594, 
    0.6063294, 0.6094063, 0.6026358, 0.5991582, 0.5982617, 0.5965938, 
    0.5982998, 0.5981609, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260328, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026052, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01193812, 0.01193812, 0.01193812, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01193812, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 0.01193812, 
    0.01893771, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 0.01193812, 
    0.01193812, 0.01193812 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.348378e-11, 3.363205e-11, 3.360314e-11, 3.372281e-11, 3.365637e-11, 
    3.373469e-11, 3.351366e-11, 3.36377e-11, 3.355845e-11, 3.349683e-11, 
    3.395502e-11, 3.372788e-11, 3.419126e-11, 3.40461e-11, 3.44108e-11, 
    3.416857e-11, 3.445965e-11, 3.440371e-11, 3.457194e-11, 3.452368e-11, 
    3.4739e-11, 3.459411e-11, 3.485067e-11, 3.470432e-11, 3.472717e-11, 
    3.458916e-11, 3.37738e-11, 3.392697e-11, 3.376467e-11, 3.37865e-11, 
    3.377667e-11, 3.36576e-11, 3.359765e-11, 3.347214e-11, 3.349487e-11, 
    3.358702e-11, 3.379607e-11, 3.372501e-11, 3.390399e-11, 3.389996e-11, 
    3.409942e-11, 3.400943e-11, 3.434511e-11, 3.424958e-11, 3.452565e-11, 
    3.445612e-11, 3.452232e-11, 3.450218e-11, 3.452248e-11, 3.44206e-11, 
    3.446417e-11, 3.437455e-11, 3.402669e-11, 3.412902e-11, 3.382384e-11, 
    3.364057e-11, 3.351895e-11, 3.343275e-11, 3.344486e-11, 3.34681e-11, 
    3.358749e-11, 3.369982e-11, 3.37855e-11, 3.384279e-11, 3.389928e-11, 
    3.407051e-11, 3.416116e-11, 3.436435e-11, 3.432764e-11, 3.438976e-11, 
    3.444917e-11, 3.454892e-11, 3.453248e-11, 3.457641e-11, 3.438794e-11, 
    3.451315e-11, 3.430645e-11, 3.436294e-11, 3.391499e-11, 3.374432e-11, 
    3.367184e-11, 3.360839e-11, 3.345421e-11, 3.356064e-11, 3.351863e-11, 
    3.361843e-11, 3.36819e-11, 3.365044e-11, 3.384432e-11, 3.376886e-11, 
    3.416648e-11, 3.399508e-11, 3.444228e-11, 3.433509e-11, 3.446787e-11, 
    3.440009e-11, 3.451618e-11, 3.441163e-11, 3.459271e-11, 3.463219e-11, 
    3.460514e-11, 3.470879e-11, 3.440563e-11, 3.452197e-11, 3.364976e-11, 
    3.365489e-11, 3.367871e-11, 3.357381e-11, 3.356738e-11, 3.347131e-11, 
    3.35567e-11, 3.35931e-11, 3.368549e-11, 3.374013e-11, 3.37921e-11, 
    3.390653e-11, 3.403437e-11, 3.421331e-11, 3.434199e-11, 3.442828e-11, 
    3.437532e-11, 3.442201e-11, 3.436974e-11, 3.43452e-11, 3.46173e-11, 
    3.446444e-11, 3.469378e-11, 3.468109e-11, 3.457719e-11, 3.468242e-11, 
    3.365842e-11, 3.36289e-11, 3.352663e-11, 3.36066e-11, 3.346079e-11, 
    3.354237e-11, 3.358925e-11, 3.377039e-11, 3.381018e-11, 3.384714e-11, 
    3.39201e-11, 3.401377e-11, 3.417832e-11, 3.432156e-11, 3.445249e-11, 
    3.444283e-11, 3.44462e-11, 3.447541e-11, 3.440291e-11, 3.448724e-11, 
    3.450136e-11, 3.446433e-11, 3.467929e-11, 3.461784e-11, 3.468068e-11, 
    3.464061e-11, 3.363844e-11, 3.368798e-11, 3.366113e-11, 3.371153e-11, 
    3.367595e-11, 3.383389e-11, 3.388123e-11, 3.410307e-11, 3.401193e-11, 
    3.415695e-11, 3.402658e-11, 3.404967e-11, 3.416157e-11, 3.403353e-11, 
    3.431357e-11, 3.41236e-11, 3.44765e-11, 3.428663e-11, 3.448834e-11, 
    3.445164e-11, 3.451228e-11, 3.456666e-11, 3.4635e-11, 3.476134e-11, 
    3.4732e-11, 3.48377e-11, 3.376189e-11, 3.382621e-11, 3.382052e-11, 
    3.388786e-11, 3.393767e-11, 3.404579e-11, 3.421929e-11, 3.415396e-11, 
    3.427378e-11, 3.429786e-11, 3.411569e-11, 3.422748e-11, 3.386895e-11, 
    3.392676e-11, 3.389229e-11, 3.376644e-11, 3.416871e-11, 3.396208e-11, 
    3.434371e-11, 3.423161e-11, 3.45588e-11, 3.439598e-11, 3.471587e-11, 
    3.485283e-11, 3.498178e-11, 3.513258e-11, 3.386131e-11, 3.38175e-11, 
    3.389581e-11, 3.400427e-11, 3.410489e-11, 3.423886e-11, 3.425253e-11, 
    3.427759e-11, 3.434258e-11, 3.439731e-11, 3.428544e-11, 3.441094e-11, 
    3.394014e-11, 3.418665e-11, 3.380052e-11, 3.391669e-11, 3.399739e-11, 
    3.396196e-11, 3.414605e-11, 3.418943e-11, 3.436596e-11, 3.427467e-11, 
    3.481892e-11, 3.457789e-11, 3.524745e-11, 3.506008e-11, 3.380218e-11, 
    3.386101e-11, 3.406607e-11, 3.396846e-11, 3.424771e-11, 3.431655e-11, 
    3.437243e-11, 3.444401e-11, 3.445166e-11, 3.44941e-11, 3.44245e-11, 
    3.449128e-11, 3.423878e-11, 3.435153e-11, 3.404224e-11, 3.41174e-11, 
    3.408278e-11, 3.404477e-11, 3.416189e-11, 3.428682e-11, 3.428944e-11, 
    3.432945e-11, 3.44424e-11, 3.42482e-11, 3.484992e-11, 3.447799e-11, 
    3.392521e-11, 3.403868e-11, 3.405486e-11, 3.401087e-11, 3.430954e-11, 
    3.420124e-11, 3.449306e-11, 3.441407e-11, 3.454338e-11, 3.44791e-11, 
    3.446956e-11, 3.438704e-11, 3.43356e-11, 3.420593e-11, 3.410041e-11, 
    3.401685e-11, 3.40362e-11, 3.412802e-11, 3.429436e-11, 3.445194e-11, 
    3.441736e-11, 3.453311e-11, 3.422673e-11, 3.435512e-11, 3.430542e-11, 
    3.443486e-11, 3.415208e-11, 3.439347e-11, 3.409039e-11, 3.411689e-11, 
    3.419899e-11, 3.436435e-11, 3.440088e-11, 3.443998e-11, 3.441578e-11, 
    3.429884e-11, 3.427965e-11, 3.419677e-11, 3.417387e-11, 3.41108e-11, 
    3.405853e-11, 3.410622e-11, 3.415625e-11, 3.429862e-11, 3.442696e-11, 
    3.4567e-11, 3.460129e-11, 3.47651e-11, 3.463168e-11, 3.485182e-11, 
    3.466458e-11, 3.498874e-11, 3.440737e-11, 3.465979e-11, 3.420274e-11, 
    3.425186e-11, 3.434081e-11, 3.454503e-11, 3.443467e-11, 3.456369e-11, 
    3.427887e-11, 3.413124e-11, 3.409304e-11, 3.402188e-11, 3.40946e-11, 
    3.408869e-11, 3.415833e-11, 3.413588e-11, 3.430325e-11, 3.421331e-11, 
    3.446887e-11, 3.456226e-11, 3.482622e-11, 3.49882e-11, 3.515327e-11, 
    3.522614e-11, 3.524833e-11, 3.525757e-11,
  1.906728e-11, 1.921124e-11, 1.918322e-11, 1.929956e-11, 1.923499e-11, 
    1.931122e-11, 1.909643e-11, 1.921696e-11, 1.913999e-11, 1.908022e-11, 
    1.952606e-11, 1.930476e-11, 1.975694e-11, 1.961508e-11, 1.997214e-11, 
    1.973483e-11, 2.002011e-11, 1.996528e-11, 2.013048e-11, 2.008311e-11, 
    2.029492e-11, 2.015236e-11, 2.040504e-11, 2.026085e-11, 2.028338e-11, 
    2.014766e-11, 1.934922e-11, 1.949846e-11, 1.934039e-11, 1.936165e-11, 
    1.935211e-11, 1.923632e-11, 1.917807e-11, 1.905629e-11, 1.907838e-11, 
    1.916783e-11, 1.937121e-11, 1.930208e-11, 1.947647e-11, 1.947252e-11, 
    1.966732e-11, 1.95794e-11, 1.990786e-11, 1.981431e-11, 2.008508e-11, 
    2.001686e-11, 2.008187e-11, 2.006215e-11, 2.008213e-11, 1.998211e-11, 
    2.002494e-11, 1.993701e-11, 1.959586e-11, 1.96959e-11, 1.939807e-11, 
    1.921978e-11, 1.910171e-11, 1.901809e-11, 1.90299e-11, 1.905243e-11, 
    1.916836e-11, 1.92776e-11, 1.9361e-11, 1.941686e-11, 1.947196e-11, 
    1.963907e-11, 1.972774e-11, 1.992679e-11, 1.989082e-11, 1.995177e-11, 
    2.001008e-11, 2.010809e-11, 2.009195e-11, 2.013517e-11, 1.995017e-11, 
    2.007305e-11, 1.987034e-11, 1.992571e-11, 1.948693e-11, 1.932072e-11, 
    1.925022e-11, 1.91886e-11, 1.903899e-11, 1.914226e-11, 1.910152e-11, 
    1.91985e-11, 1.926021e-11, 1.922968e-11, 1.941839e-11, 1.934494e-11, 
    1.9733e-11, 1.956551e-11, 2.000327e-11, 1.98982e-11, 2.002849e-11, 
    1.996197e-11, 2.007599e-11, 1.997336e-11, 2.015127e-11, 2.019008e-11, 
    2.016355e-11, 2.026552e-11, 1.996768e-11, 2.008187e-11, 1.922882e-11, 
    1.92338e-11, 1.9257e-11, 1.91551e-11, 1.914888e-11, 1.905569e-11, 
    1.91386e-11, 1.917395e-11, 1.926379e-11, 1.9317e-11, 1.936763e-11, 
    1.947914e-11, 1.960393e-11, 1.977894e-11, 1.9905e-11, 1.998968e-11, 
    1.993774e-11, 1.998359e-11, 1.993234e-11, 1.990834e-11, 2.017553e-11, 
    2.002534e-11, 2.025084e-11, 2.023834e-11, 2.01362e-11, 2.023975e-11, 
    1.92373e-11, 1.920866e-11, 1.910933e-11, 1.918705e-11, 1.904555e-11, 
    1.91247e-11, 1.917027e-11, 1.934647e-11, 1.938527e-11, 1.942126e-11, 
    1.949243e-11, 1.95839e-11, 1.974473e-11, 1.988505e-11, 2.001347e-11, 
    2.000405e-11, 2.000737e-11, 2.003609e-11, 1.996497e-11, 2.004778e-11, 
    2.006168e-11, 2.002532e-11, 2.023667e-11, 2.017621e-11, 2.023808e-11, 
    2.01987e-11, 1.921796e-11, 1.926617e-11, 1.924012e-11, 1.928913e-11, 
    1.925459e-11, 1.940831e-11, 1.945449e-11, 1.967109e-11, 1.95821e-11, 
    1.972381e-11, 1.959648e-11, 1.961901e-11, 1.972843e-11, 1.960335e-11, 
    1.987731e-11, 1.969142e-11, 2.003721e-11, 1.985103e-11, 2.004889e-11, 
    2.001291e-11, 2.00725e-11, 2.012592e-11, 2.019319e-11, 2.031753e-11, 
    2.028872e-11, 2.039286e-11, 1.933813e-11, 1.940081e-11, 1.939529e-11, 
    1.946096e-11, 1.950958e-11, 1.961512e-11, 1.978481e-11, 1.972094e-11, 
    1.983826e-11, 1.986184e-11, 1.968362e-11, 1.979297e-11, 1.944281e-11, 
    1.949922e-11, 1.946563e-11, 1.934307e-11, 1.973564e-11, 1.953381e-11, 
    1.990709e-11, 1.979732e-11, 2.01183e-11, 1.995843e-11, 2.027286e-11, 
    2.04078e-11, 2.05351e-11, 2.06842e-11, 1.943505e-11, 1.939243e-11, 
    1.946878e-11, 1.957459e-11, 1.967296e-11, 1.980401e-11, 1.981744e-11, 
    1.984203e-11, 1.990578e-11, 1.995944e-11, 1.98498e-11, 1.997289e-11, 
    1.951231e-11, 1.97532e-11, 1.937632e-11, 1.948952e-11, 1.956835e-11, 
    1.953376e-11, 1.971364e-11, 1.975612e-11, 1.992909e-11, 1.983961e-11, 
    2.037446e-11, 2.01372e-11, 2.079799e-11, 2.061257e-11, 1.937754e-11, 
    1.943491e-11, 1.963505e-11, 1.953973e-11, 1.981277e-11, 1.988019e-11, 
    1.993505e-11, 2.000527e-11, 2.001286e-11, 2.00545e-11, 1.998627e-11, 
    2.005181e-11, 1.980429e-11, 1.991476e-11, 1.961213e-11, 1.968564e-11, 
    1.965181e-11, 1.961473e-11, 1.972926e-11, 1.985153e-11, 1.985415e-11, 
    1.989341e-11, 2.000419e-11, 1.981388e-11, 2.040515e-11, 2.003925e-11, 
    1.949754e-11, 1.960833e-11, 1.962418e-11, 1.958122e-11, 1.987343e-11, 
    1.976737e-11, 2.005349e-11, 1.997602e-11, 2.010301e-11, 2.003987e-11, 
    2.003058e-11, 1.99496e-11, 1.989925e-11, 1.977223e-11, 1.966909e-11, 
    1.958745e-11, 1.960642e-11, 1.969614e-11, 1.985902e-11, 2.001354e-11, 
    1.997965e-11, 2.009335e-11, 1.979293e-11, 1.99187e-11, 1.987006e-11, 
    1.999699e-11, 1.971924e-11, 1.995565e-11, 1.965897e-11, 1.968492e-11, 
    1.976527e-11, 1.992724e-11, 1.996314e-11, 2.00015e-11, 1.997783e-11, 
    1.986316e-11, 1.98444e-11, 1.976331e-11, 1.974094e-11, 1.967927e-11, 
    1.962826e-11, 1.967486e-11, 1.972385e-11, 1.986321e-11, 1.99891e-11, 
    2.012668e-11, 2.01604e-11, 2.032166e-11, 2.019034e-11, 2.040719e-11, 
    2.022277e-11, 2.054239e-11, 1.996939e-11, 2.021736e-11, 1.976893e-11, 
    1.981707e-11, 1.990423e-11, 2.01047e-11, 1.999639e-11, 2.012308e-11, 
    1.984366e-11, 1.969924e-11, 1.966194e-11, 1.959241e-11, 1.966353e-11, 
    1.965774e-11, 1.972588e-11, 1.970397e-11, 1.986784e-11, 1.977976e-11, 
    2.003035e-11, 2.012208e-11, 2.038193e-11, 2.054181e-11, 2.070501e-11, 
    2.07772e-11, 2.079919e-11, 2.080839e-11,
  1.783518e-11, 1.799284e-11, 1.796215e-11, 1.808964e-11, 1.801887e-11, 
    1.810242e-11, 1.78671e-11, 1.799911e-11, 1.791479e-11, 1.784936e-11, 
    1.833814e-11, 1.809534e-11, 1.85918e-11, 1.84359e-11, 1.882859e-11, 
    1.85675e-11, 1.888142e-11, 1.882105e-11, 1.900303e-11, 1.895082e-11, 
    1.918437e-11, 1.902715e-11, 1.930591e-11, 1.914678e-11, 1.917163e-11, 
    1.902197e-11, 1.814409e-11, 1.830783e-11, 1.813441e-11, 1.815772e-11, 
    1.814726e-11, 1.802033e-11, 1.795651e-11, 1.782316e-11, 1.784734e-11, 
    1.794529e-11, 1.81682e-11, 1.809241e-11, 1.828369e-11, 1.827937e-11, 
    1.849329e-11, 1.839671e-11, 1.875783e-11, 1.86549e-11, 1.8953e-11, 
    1.887784e-11, 1.894947e-11, 1.892774e-11, 1.894975e-11, 1.883957e-11, 
    1.888674e-11, 1.878992e-11, 1.841478e-11, 1.85247e-11, 1.819767e-11, 
    1.800221e-11, 1.787288e-11, 1.778135e-11, 1.779428e-11, 1.781893e-11, 
    1.794587e-11, 1.806556e-11, 1.815701e-11, 1.821828e-11, 1.827874e-11, 
    1.846225e-11, 1.85597e-11, 1.877867e-11, 1.873908e-11, 1.880617e-11, 
    1.887037e-11, 1.897836e-11, 1.896056e-11, 1.90082e-11, 1.880441e-11, 
    1.893975e-11, 1.871654e-11, 1.877748e-11, 1.829518e-11, 1.811284e-11, 
    1.803556e-11, 1.796805e-11, 1.780422e-11, 1.791729e-11, 1.787268e-11, 
    1.797888e-11, 1.80465e-11, 1.801305e-11, 1.821996e-11, 1.81394e-11, 
    1.856549e-11, 1.838145e-11, 1.886288e-11, 1.87472e-11, 1.889065e-11, 
    1.88174e-11, 1.894298e-11, 1.882994e-11, 1.902594e-11, 1.906873e-11, 
    1.903949e-11, 1.915194e-11, 1.882368e-11, 1.894946e-11, 1.801211e-11, 
    1.801756e-11, 1.804299e-11, 1.793135e-11, 1.792453e-11, 1.78225e-11, 
    1.791327e-11, 1.795199e-11, 1.805043e-11, 1.810876e-11, 1.816429e-11, 
    1.828662e-11, 1.842365e-11, 1.861599e-11, 1.875469e-11, 1.884791e-11, 
    1.879073e-11, 1.88412e-11, 1.878478e-11, 1.875836e-11, 1.905269e-11, 
    1.888718e-11, 1.913575e-11, 1.912196e-11, 1.900933e-11, 1.912351e-11, 
    1.80214e-11, 1.799001e-11, 1.788123e-11, 1.796634e-11, 1.78114e-11, 
    1.789806e-11, 1.794796e-11, 1.814108e-11, 1.818363e-11, 1.822311e-11, 
    1.830121e-11, 1.840165e-11, 1.857838e-11, 1.873274e-11, 1.887411e-11, 
    1.886374e-11, 1.886739e-11, 1.889903e-11, 1.88207e-11, 1.89119e-11, 
    1.892722e-11, 1.888717e-11, 1.912011e-11, 1.905344e-11, 1.912166e-11, 
    1.907824e-11, 1.800021e-11, 1.805304e-11, 1.802449e-11, 1.80782e-11, 
    1.804035e-11, 1.820891e-11, 1.825957e-11, 1.849744e-11, 1.839967e-11, 
    1.855538e-11, 1.841546e-11, 1.844022e-11, 1.856046e-11, 1.842301e-11, 
    1.872421e-11, 1.851978e-11, 1.890026e-11, 1.86953e-11, 1.891313e-11, 
    1.88735e-11, 1.893914e-11, 1.8998e-11, 1.907217e-11, 1.920932e-11, 
    1.917753e-11, 1.929246e-11, 1.813193e-11, 1.820068e-11, 1.819462e-11, 
    1.826668e-11, 1.832004e-11, 1.843594e-11, 1.862245e-11, 1.855222e-11, 
    1.868124e-11, 1.870718e-11, 1.851121e-11, 1.863143e-11, 1.824675e-11, 
    1.830867e-11, 1.827179e-11, 1.813734e-11, 1.856839e-11, 1.834664e-11, 
    1.875699e-11, 1.863621e-11, 1.89896e-11, 1.88135e-11, 1.916003e-11, 
    1.930896e-11, 1.944957e-11, 1.961441e-11, 1.823825e-11, 1.819148e-11, 
    1.827525e-11, 1.839142e-11, 1.849949e-11, 1.864357e-11, 1.865834e-11, 
    1.868539e-11, 1.875554e-11, 1.881461e-11, 1.869395e-11, 1.882943e-11, 
    1.832304e-11, 1.858769e-11, 1.817381e-11, 1.829802e-11, 1.838457e-11, 
    1.834658e-11, 1.85442e-11, 1.859091e-11, 1.87812e-11, 1.868273e-11, 
    1.927216e-11, 1.901044e-11, 1.974031e-11, 1.95352e-11, 1.817515e-11, 
    1.823809e-11, 1.845783e-11, 1.835314e-11, 1.865321e-11, 1.872738e-11, 
    1.878777e-11, 1.886508e-11, 1.887343e-11, 1.891931e-11, 1.884416e-11, 
    1.891634e-11, 1.864388e-11, 1.876543e-11, 1.843266e-11, 1.851342e-11, 
    1.847625e-11, 1.843551e-11, 1.856137e-11, 1.869584e-11, 1.869872e-11, 
    1.874193e-11, 1.88639e-11, 1.865443e-11, 1.930603e-11, 1.890251e-11, 
    1.830682e-11, 1.842848e-11, 1.844589e-11, 1.83987e-11, 1.871994e-11, 
    1.860327e-11, 1.891819e-11, 1.883286e-11, 1.897276e-11, 1.890319e-11, 
    1.889296e-11, 1.880378e-11, 1.874835e-11, 1.860861e-11, 1.849524e-11, 
    1.840555e-11, 1.842639e-11, 1.852497e-11, 1.870408e-11, 1.887419e-11, 
    1.883687e-11, 1.896211e-11, 1.863138e-11, 1.876976e-11, 1.871623e-11, 
    1.885596e-11, 1.855036e-11, 1.881045e-11, 1.848412e-11, 1.851263e-11, 
    1.860096e-11, 1.877916e-11, 1.881869e-11, 1.886092e-11, 1.883486e-11, 
    1.870864e-11, 1.8688e-11, 1.859881e-11, 1.857422e-11, 1.850642e-11, 
    1.845037e-11, 1.850158e-11, 1.855542e-11, 1.870869e-11, 1.884727e-11, 
    1.899884e-11, 1.903601e-11, 1.921387e-11, 1.906903e-11, 1.930829e-11, 
    1.910478e-11, 1.945763e-11, 1.882557e-11, 1.909882e-11, 1.860499e-11, 
    1.865793e-11, 1.875384e-11, 1.897462e-11, 1.88553e-11, 1.899487e-11, 
    1.868719e-11, 1.852837e-11, 1.848738e-11, 1.841099e-11, 1.848913e-11, 
    1.848277e-11, 1.855766e-11, 1.853358e-11, 1.871379e-11, 1.86169e-11, 
    1.88927e-11, 1.899377e-11, 1.92804e-11, 1.945699e-11, 1.963743e-11, 
    1.971731e-11, 1.974164e-11, 1.975182e-11,
  1.829491e-11, 1.846854e-11, 1.843472e-11, 1.857521e-11, 1.849721e-11, 
    1.85893e-11, 1.833005e-11, 1.847545e-11, 1.838256e-11, 1.831051e-11, 
    1.884932e-11, 1.858149e-11, 1.912945e-11, 1.895721e-11, 1.939129e-11, 
    1.91026e-11, 1.944975e-11, 1.938293e-11, 1.958437e-11, 1.952655e-11, 
    1.97853e-11, 1.961107e-11, 1.992006e-11, 1.974362e-11, 1.977117e-11, 
    1.960534e-11, 1.863524e-11, 1.881587e-11, 1.862456e-11, 1.865026e-11, 
    1.863873e-11, 1.849882e-11, 1.842851e-11, 1.828167e-11, 1.830829e-11, 
    1.841616e-11, 1.866183e-11, 1.857826e-11, 1.878921e-11, 1.878443e-11, 
    1.90206e-11, 1.891395e-11, 1.9313e-11, 1.919917e-11, 1.952897e-11, 
    1.944577e-11, 1.952506e-11, 1.9501e-11, 1.952537e-11, 1.940343e-11, 
    1.945563e-11, 1.934849e-11, 1.89339e-11, 1.90553e-11, 1.869432e-11, 
    1.847886e-11, 1.833641e-11, 1.823565e-11, 1.824988e-11, 1.827702e-11, 
    1.841679e-11, 1.854867e-11, 1.864947e-11, 1.871705e-11, 1.878375e-11, 
    1.898634e-11, 1.909398e-11, 1.933605e-11, 1.929226e-11, 1.936648e-11, 
    1.943751e-11, 1.955704e-11, 1.953734e-11, 1.95901e-11, 1.936452e-11, 
    1.95143e-11, 1.926733e-11, 1.933473e-11, 1.880191e-11, 1.860078e-11, 
    1.851562e-11, 1.844122e-11, 1.826082e-11, 1.838531e-11, 1.833619e-11, 
    1.845315e-11, 1.852766e-11, 1.849079e-11, 1.87189e-11, 1.863006e-11, 
    1.910037e-11, 1.88971e-11, 1.942922e-11, 1.930124e-11, 1.945995e-11, 
    1.937889e-11, 1.951788e-11, 1.939277e-11, 1.960974e-11, 1.965714e-11, 
    1.962475e-11, 1.974933e-11, 1.938584e-11, 1.952506e-11, 1.848976e-11, 
    1.849577e-11, 1.852378e-11, 1.84008e-11, 1.839329e-11, 1.828094e-11, 
    1.838089e-11, 1.842353e-11, 1.853198e-11, 1.859628e-11, 1.86575e-11, 
    1.879244e-11, 1.89437e-11, 1.915618e-11, 1.930952e-11, 1.941264e-11, 
    1.934938e-11, 1.940523e-11, 1.93428e-11, 1.931358e-11, 1.963938e-11, 
    1.945612e-11, 1.973139e-11, 1.971611e-11, 1.959135e-11, 1.971783e-11, 
    1.849999e-11, 1.846541e-11, 1.83456e-11, 1.843933e-11, 1.826873e-11, 
    1.836413e-11, 1.84191e-11, 1.863192e-11, 1.867883e-11, 1.872238e-11, 
    1.880854e-11, 1.89194e-11, 1.911461e-11, 1.928525e-11, 1.944164e-11, 
    1.943016e-11, 1.94342e-11, 1.946922e-11, 1.938254e-11, 1.948347e-11, 
    1.950043e-11, 1.945609e-11, 1.971406e-11, 1.96402e-11, 1.971578e-11, 
    1.966767e-11, 1.847665e-11, 1.853487e-11, 1.85034e-11, 1.85626e-11, 
    1.852088e-11, 1.870672e-11, 1.876261e-11, 1.902519e-11, 1.891721e-11, 
    1.908919e-11, 1.893465e-11, 1.896199e-11, 1.909482e-11, 1.894298e-11, 
    1.927582e-11, 1.904987e-11, 1.947058e-11, 1.924386e-11, 1.948483e-11, 
    1.944097e-11, 1.951362e-11, 1.95788e-11, 1.966094e-11, 1.981295e-11, 
    1.97777e-11, 1.990514e-11, 1.862182e-11, 1.869764e-11, 1.869096e-11, 
    1.877044e-11, 1.882932e-11, 1.895726e-11, 1.916331e-11, 1.90857e-11, 
    1.92283e-11, 1.925698e-11, 1.904039e-11, 1.917324e-11, 1.874846e-11, 
    1.881678e-11, 1.877608e-11, 1.86278e-11, 1.910357e-11, 1.885869e-11, 
    1.931206e-11, 1.917852e-11, 1.95695e-11, 1.937459e-11, 1.975831e-11, 
    1.992344e-11, 2.007945e-11, 2.026251e-11, 1.873907e-11, 1.868749e-11, 
    1.87799e-11, 1.890812e-11, 1.902745e-11, 1.918666e-11, 1.920298e-11, 
    1.923289e-11, 1.931046e-11, 1.93758e-11, 1.924235e-11, 1.93922e-11, 
    1.883265e-11, 1.91249e-11, 1.866801e-11, 1.880503e-11, 1.890055e-11, 
    1.885862e-11, 1.907684e-11, 1.912845e-11, 1.933885e-11, 1.922995e-11, 
    1.988263e-11, 1.959258e-11, 2.040242e-11, 2.017453e-11, 1.866948e-11, 
    1.873889e-11, 1.898144e-11, 1.886585e-11, 1.919731e-11, 1.927932e-11, 
    1.934611e-11, 1.943165e-11, 1.944089e-11, 1.949167e-11, 1.94085e-11, 
    1.948838e-11, 1.9187e-11, 1.93214e-11, 1.895364e-11, 1.904284e-11, 
    1.900178e-11, 1.895679e-11, 1.90958e-11, 1.924445e-11, 1.924763e-11, 
    1.929541e-11, 1.943037e-11, 1.919865e-11, 1.992022e-11, 1.94731e-11, 
    1.881473e-11, 1.894904e-11, 1.896825e-11, 1.891615e-11, 1.927109e-11, 
    1.914211e-11, 1.949044e-11, 1.9396e-11, 1.955084e-11, 1.947383e-11, 
    1.946251e-11, 1.936383e-11, 1.930251e-11, 1.914802e-11, 1.902275e-11, 
    1.89237e-11, 1.894671e-11, 1.90556e-11, 1.925356e-11, 1.944173e-11, 
    1.940044e-11, 1.953906e-11, 1.917318e-11, 1.93262e-11, 1.926699e-11, 
    1.942156e-11, 1.908364e-11, 1.937122e-11, 1.901046e-11, 1.904196e-11, 
    1.913956e-11, 1.93366e-11, 1.938032e-11, 1.942706e-11, 1.939821e-11, 
    1.92586e-11, 1.923577e-11, 1.913718e-11, 1.911001e-11, 1.90351e-11, 
    1.89732e-11, 1.902976e-11, 1.908924e-11, 1.925865e-11, 1.941194e-11, 
    1.957973e-11, 1.962089e-11, 1.981801e-11, 1.965748e-11, 1.992272e-11, 
    1.969712e-11, 2.008842e-11, 1.938795e-11, 1.969049e-11, 1.914401e-11, 
    1.920252e-11, 1.930859e-11, 1.955291e-11, 1.942083e-11, 1.957534e-11, 
    1.923487e-11, 1.905936e-11, 1.901407e-11, 1.892972e-11, 1.9016e-11, 
    1.900897e-11, 1.90917e-11, 1.90651e-11, 1.926429e-11, 1.915717e-11, 
    1.946222e-11, 1.957412e-11, 1.989176e-11, 2.00877e-11, 2.028808e-11, 
    2.037684e-11, 2.04039e-11, 2.041521e-11,
  1.973493e-11, 1.991887e-11, 1.988303e-11, 2.003196e-11, 1.994926e-11, 
    2.00469e-11, 1.977214e-11, 1.99262e-11, 1.982777e-11, 1.975144e-11, 
    2.03228e-11, 2.003862e-11, 2.062037e-11, 2.043735e-11, 2.089888e-11, 
    2.059184e-11, 2.09611e-11, 2.088997e-11, 2.110445e-11, 2.104288e-11, 
    2.131863e-11, 2.113291e-11, 2.146237e-11, 2.127418e-11, 2.130357e-11, 
    2.11268e-11, 2.009561e-11, 2.02873e-11, 2.008429e-11, 2.011155e-11, 
    2.009931e-11, 1.995097e-11, 1.987647e-11, 1.97209e-11, 1.974909e-11, 
    1.986337e-11, 2.012382e-11, 2.003518e-11, 2.025897e-11, 2.02539e-11, 
    2.050469e-11, 2.039139e-11, 2.081556e-11, 2.069449e-11, 2.104544e-11, 
    2.095686e-11, 2.104128e-11, 2.101566e-11, 2.104162e-11, 2.091179e-11, 
    2.096736e-11, 2.085332e-11, 2.041258e-11, 2.054156e-11, 2.015828e-11, 
    1.992983e-11, 1.977889e-11, 1.967218e-11, 1.968724e-11, 1.971598e-11, 
    1.986404e-11, 2.000381e-11, 2.01107e-11, 2.018239e-11, 2.025317e-11, 
    2.04683e-11, 2.058267e-11, 2.08401e-11, 2.079349e-11, 2.087247e-11, 
    2.094806e-11, 2.107535e-11, 2.105437e-11, 2.111056e-11, 2.087037e-11, 
    2.102983e-11, 2.076697e-11, 2.083868e-11, 2.027248e-11, 2.005907e-11, 
    1.996879e-11, 1.988992e-11, 1.969883e-11, 1.983069e-11, 1.977865e-11, 
    1.990257e-11, 1.998154e-11, 1.994246e-11, 2.018435e-11, 2.009012e-11, 
    2.058946e-11, 2.037351e-11, 2.093924e-11, 2.080305e-11, 2.097196e-11, 
    2.088567e-11, 2.103365e-11, 2.090044e-11, 2.113149e-11, 2.118201e-11, 
    2.114748e-11, 2.128027e-11, 2.089307e-11, 2.104129e-11, 1.994136e-11, 
    1.994774e-11, 1.997743e-11, 1.984709e-11, 1.983913e-11, 1.972013e-11, 
    1.9826e-11, 1.987118e-11, 1.998612e-11, 2.00543e-11, 2.011922e-11, 
    2.02624e-11, 2.0423e-11, 2.064878e-11, 2.081186e-11, 2.09216e-11, 
    2.085427e-11, 2.09137e-11, 2.084727e-11, 2.081617e-11, 2.116307e-11, 
    2.096788e-11, 2.126114e-11, 2.124485e-11, 2.11119e-11, 2.124668e-11, 
    1.995221e-11, 1.991556e-11, 1.978862e-11, 1.988792e-11, 1.97072e-11, 
    1.980825e-11, 1.986649e-11, 2.009209e-11, 2.014184e-11, 2.018805e-11, 
    2.027949e-11, 2.039718e-11, 2.060459e-11, 2.078604e-11, 2.095247e-11, 
    2.094024e-11, 2.094455e-11, 2.098183e-11, 2.088956e-11, 2.0997e-11, 
    2.101506e-11, 2.096785e-11, 2.124267e-11, 2.116394e-11, 2.12445e-11, 
    2.119322e-11, 1.992747e-11, 1.998918e-11, 1.995582e-11, 2.001858e-11, 
    1.997436e-11, 2.017144e-11, 2.023075e-11, 2.050957e-11, 2.039486e-11, 
    2.057758e-11, 2.041338e-11, 2.044242e-11, 2.058357e-11, 2.042223e-11, 
    2.077602e-11, 2.05358e-11, 2.098328e-11, 2.074203e-11, 2.099845e-11, 
    2.095174e-11, 2.10291e-11, 2.109853e-11, 2.118605e-11, 2.134811e-11, 
    2.131052e-11, 2.144645e-11, 2.008138e-11, 2.01618e-11, 2.015471e-11, 
    2.023904e-11, 2.030155e-11, 2.043739e-11, 2.065636e-11, 2.057386e-11, 
    2.072546e-11, 2.075597e-11, 2.052571e-11, 2.066692e-11, 2.021572e-11, 
    2.028824e-11, 2.024504e-11, 2.008772e-11, 2.059287e-11, 2.033273e-11, 
    2.081457e-11, 2.067253e-11, 2.108862e-11, 2.08811e-11, 2.128984e-11, 
    2.1466e-11, 2.163252e-11, 2.182811e-11, 2.020576e-11, 2.015103e-11, 
    2.024908e-11, 2.038521e-11, 2.051196e-11, 2.068118e-11, 2.069853e-11, 
    2.073034e-11, 2.081286e-11, 2.088238e-11, 2.074041e-11, 2.089983e-11, 
    2.03051e-11, 2.061553e-11, 2.013037e-11, 2.027578e-11, 2.037717e-11, 
    2.033265e-11, 2.056444e-11, 2.061929e-11, 2.084307e-11, 2.072721e-11, 
    2.142245e-11, 2.111322e-11, 2.19777e-11, 2.173409e-11, 2.013193e-11, 
    2.020557e-11, 2.046308e-11, 2.034032e-11, 2.06925e-11, 2.077973e-11, 
    2.085078e-11, 2.094183e-11, 2.095167e-11, 2.100574e-11, 2.091718e-11, 
    2.100223e-11, 2.068154e-11, 2.08245e-11, 2.043354e-11, 2.052831e-11, 
    2.048468e-11, 2.043689e-11, 2.05846e-11, 2.074265e-11, 2.074602e-11, 
    2.079685e-11, 2.094051e-11, 2.069393e-11, 2.146258e-11, 2.0986e-11, 
    2.028605e-11, 2.042867e-11, 2.044907e-11, 2.039373e-11, 2.077097e-11, 
    2.063383e-11, 2.100442e-11, 2.090388e-11, 2.106875e-11, 2.098673e-11, 
    2.097468e-11, 2.086964e-11, 2.08044e-11, 2.064011e-11, 2.050697e-11, 
    2.040175e-11, 2.042619e-11, 2.054187e-11, 2.075234e-11, 2.095257e-11, 
    2.090861e-11, 2.105619e-11, 2.066685e-11, 2.082961e-11, 2.076662e-11, 
    2.093108e-11, 2.057167e-11, 2.087755e-11, 2.049391e-11, 2.052738e-11, 
    2.063111e-11, 2.084068e-11, 2.088719e-11, 2.093694e-11, 2.090623e-11, 
    2.075769e-11, 2.073341e-11, 2.062858e-11, 2.05997e-11, 2.052009e-11, 
    2.045432e-11, 2.051441e-11, 2.057762e-11, 2.075775e-11, 2.092086e-11, 
    2.109952e-11, 2.114337e-11, 2.135353e-11, 2.118238e-11, 2.146525e-11, 
    2.122465e-11, 2.164213e-11, 2.089533e-11, 2.121757e-11, 2.063583e-11, 
    2.069805e-11, 2.081088e-11, 2.107097e-11, 2.093031e-11, 2.109486e-11, 
    2.073246e-11, 2.054588e-11, 2.049774e-11, 2.040814e-11, 2.049979e-11, 
    2.049233e-11, 2.058024e-11, 2.055196e-11, 2.076374e-11, 2.064983e-11, 
    2.097438e-11, 2.109355e-11, 2.143218e-11, 2.164133e-11, 2.185542e-11, 
    2.195034e-11, 2.197928e-11, 2.199138e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
