netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/21/14 13:05:54" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/21/14" ;

 time_written =
  "13:05:54" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.006537e-14, 5.020265e-14, 5.017598e-14, 5.028662e-14, 5.022528e-14, 
    5.029769e-14, 5.009324e-14, 5.020808e-14, 5.013479e-14, 5.007777e-14, 
    5.050107e-14, 5.029156e-14, 5.071864e-14, 5.058518e-14, 5.092029e-14, 
    5.069785e-14, 5.096511e-14, 5.091392e-14, 5.106806e-14, 5.102392e-14, 
    5.122079e-14, 5.108843e-14, 5.132283e-14, 5.118922e-14, 5.121011e-14, 
    5.108405e-14, 5.033379e-14, 5.047498e-14, 5.032541e-14, 5.034555e-14, 
    5.033653e-14, 5.022653e-14, 5.017103e-14, 5.005491e-14, 5.007601e-14, 
    5.016131e-14, 5.035461e-14, 5.028905e-14, 5.045433e-14, 5.04506e-14, 
    5.06344e-14, 5.055155e-14, 5.086021e-14, 5.077255e-14, 5.102576e-14, 
    5.096211e-14, 5.102276e-14, 5.100438e-14, 5.1023e-14, 5.092965e-14, 
    5.096965e-14, 5.088749e-14, 5.056706e-14, 5.066128e-14, 5.038009e-14, 
    5.021072e-14, 5.009827e-14, 5.001838e-14, 5.002968e-14, 5.00512e-14, 
    5.016181e-14, 5.026579e-14, 5.034497e-14, 5.039791e-14, 5.045006e-14, 
    5.060771e-14, 5.06912e-14, 5.08779e-14, 5.084426e-14, 5.090128e-14, 
    5.095578e-14, 5.104719e-14, 5.103216e-14, 5.107241e-14, 5.08998e-14, 
    5.101452e-14, 5.082509e-14, 5.087692e-14, 5.046407e-14, 5.030675e-14, 
    5.023969e-14, 5.01811e-14, 5.003836e-14, 5.013694e-14, 5.009808e-14, 
    5.019055e-14, 5.024925e-14, 5.022023e-14, 5.039936e-14, 5.032973e-14, 
    5.069615e-14, 5.053841e-14, 5.094942e-14, 5.085117e-14, 5.097297e-14, 
    5.091084e-14, 5.101727e-14, 5.092149e-14, 5.10874e-14, 5.112348e-14, 
    5.109882e-14, 5.119359e-14, 5.091617e-14, 5.102275e-14, 5.021941e-14, 
    5.022414e-14, 5.024621e-14, 5.014918e-14, 5.014325e-14, 5.005432e-14, 
    5.013346e-14, 5.016714e-14, 5.025267e-14, 5.030321e-14, 5.035125e-14, 
    5.045684e-14, 5.057466e-14, 5.073932e-14, 5.085754e-14, 5.093673e-14, 
    5.088819e-14, 5.093105e-14, 5.088313e-14, 5.086068e-14, 5.110995e-14, 
    5.097001e-14, 5.117996e-14, 5.116836e-14, 5.107336e-14, 5.116967e-14, 
    5.022747e-14, 5.020022e-14, 5.010555e-14, 5.017964e-14, 5.004464e-14, 
    5.01202e-14, 5.016362e-14, 5.033115e-14, 5.036798e-14, 5.040207e-14, 
    5.046942e-14, 5.055579e-14, 5.07072e-14, 5.083885e-14, 5.095896e-14, 
    5.095017e-14, 5.095326e-14, 5.098006e-14, 5.091364e-14, 5.099097e-14, 
    5.100393e-14, 5.097002e-14, 5.11668e-14, 5.111061e-14, 5.116811e-14, 
    5.113153e-14, 5.020908e-14, 5.025493e-14, 5.023015e-14, 5.027673e-14, 
    5.024391e-14, 5.038977e-14, 5.043348e-14, 5.063791e-14, 5.055408e-14, 
    5.068752e-14, 5.056766e-14, 5.058889e-14, 5.06918e-14, 5.057415e-14, 
    5.083156e-14, 5.065702e-14, 5.09811e-14, 5.08069e-14, 5.099201e-14, 
    5.095844e-14, 5.101404e-14, 5.106379e-14, 5.11264e-14, 5.124181e-14, 
    5.12151e-14, 5.131159e-14, 5.032327e-14, 5.038268e-14, 5.037748e-14, 
    5.043966e-14, 5.048562e-14, 5.058524e-14, 5.074485e-14, 5.068486e-14, 
    5.079501e-14, 5.081711e-14, 5.064976e-14, 5.07525e-14, 5.042246e-14, 
    5.047579e-14, 5.044406e-14, 5.032794e-14, 5.069864e-14, 5.050848e-14, 
    5.085949e-14, 5.07566e-14, 5.10567e-14, 5.090749e-14, 5.120039e-14, 
    5.132534e-14, 5.1443e-14, 5.158021e-14, 5.041513e-14, 5.037477e-14, 
    5.044706e-14, 5.054697e-14, 5.063971e-14, 5.076287e-14, 5.077549e-14, 
    5.079854e-14, 5.085828e-14, 5.090847e-14, 5.08058e-14, 5.092105e-14, 
    5.048809e-14, 5.071515e-14, 5.035948e-14, 5.046661e-14, 5.05411e-14, 
    5.050846e-14, 5.0678e-14, 5.071793e-14, 5.088006e-14, 5.079629e-14, 
    5.129449e-14, 5.107426e-14, 5.16847e-14, 5.151434e-14, 5.036066e-14, 
    5.041501e-14, 5.060398e-14, 5.05141e-14, 5.077111e-14, 5.08343e-14, 
    5.088568e-14, 5.095127e-14, 5.095838e-14, 5.099724e-14, 5.093355e-14, 
    5.099473e-14, 5.076314e-14, 5.086668e-14, 5.058243e-14, 5.065164e-14, 
    5.061982e-14, 5.058488e-14, 5.069268e-14, 5.080741e-14, 5.080991e-14, 
    5.084667e-14, 5.095012e-14, 5.077215e-14, 5.132279e-14, 5.098287e-14, 
    5.047425e-14, 5.057878e-14, 5.059377e-14, 5.055328e-14, 5.082796e-14, 
    5.072848e-14, 5.09963e-14, 5.092397e-14, 5.104247e-14, 5.098359e-14, 
    5.097493e-14, 5.089928e-14, 5.085215e-14, 5.073303e-14, 5.063607e-14, 
    5.055916e-14, 5.057705e-14, 5.066152e-14, 5.081443e-14, 5.0959e-14, 
    5.092734e-14, 5.103347e-14, 5.075249e-14, 5.087034e-14, 5.082478e-14, 
    5.094356e-14, 5.068325e-14, 5.090479e-14, 5.062656e-14, 5.065098e-14, 
    5.072651e-14, 5.08783e-14, 5.091194e-14, 5.094775e-14, 5.092566e-14, 
    5.081832e-14, 5.080075e-14, 5.072468e-14, 5.070365e-14, 5.064567e-14, 
    5.059763e-14, 5.064151e-14, 5.068757e-14, 5.081839e-14, 5.093617e-14, 
    5.10645e-14, 5.10959e-14, 5.124555e-14, 5.112367e-14, 5.132467e-14, 
    5.11537e-14, 5.144959e-14, 5.091769e-14, 5.114877e-14, 5.072996e-14, 
    5.077514e-14, 5.085678e-14, 5.104398e-14, 5.0943e-14, 5.106111e-14, 
    5.080007e-14, 5.066441e-14, 5.062935e-14, 5.056382e-14, 5.063085e-14, 
    5.06254e-14, 5.068951e-14, 5.066891e-14, 5.082273e-14, 5.074013e-14, 
    5.09747e-14, 5.106019e-14, 5.130146e-14, 5.144914e-14, 5.15994e-14, 
    5.166566e-14, 5.168583e-14, 5.169425e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.151354e-15, -7.140393e-15, -7.142523e-15, -7.133691e-15, -7.13859e-15, 
    -7.132808e-15, -7.149133e-15, -7.139957e-15, -7.145814e-15, 
    -7.150369e-15, -7.116579e-15, -7.133297e-15, -7.099275e-15, 
    -7.109901e-15, -7.083245e-15, -7.100925e-15, -7.079687e-15, 
    -7.083759e-15, -7.071522e-15, -7.075025e-15, -7.059392e-15, 
    -7.069905e-15, -7.05131e-15, -7.061903e-15, -7.060243e-15, -7.070252e-15, 
    -7.129933e-15, -7.118656e-15, -7.130601e-15, -7.128992e-15, 
    -7.129714e-15, -7.138488e-15, -7.142911e-15, -7.152195e-15, -7.15051e-15, 
    -7.143692e-15, -7.128268e-15, -7.133502e-15, -7.120327e-15, 
    -7.120624e-15, -7.105984e-15, -7.112581e-15, -7.088026e-15, 
    -7.094997e-15, -7.074879e-15, -7.079932e-15, -7.075115e-15, 
    -7.076576e-15, -7.075096e-15, -7.082509e-15, -7.079332e-15, 
    -7.085859e-15, -7.111344e-15, -7.103843e-15, -7.12624e-15, -7.139738e-15, 
    -7.148729e-15, -7.155113e-15, -7.154211e-15, -7.152489e-15, 
    -7.143652e-15, -7.135358e-15, -7.129043e-15, -7.124823e-15, 
    -7.120667e-15, -7.108094e-15, -7.101457e-15, -7.086616e-15, 
    -7.089295e-15, -7.08476e-15, -7.080435e-15, -7.073176e-15, -7.07437e-15, 
    -7.071173e-15, -7.084882e-15, -7.075767e-15, -7.090821e-15, 
    -7.086699e-15, -7.119525e-15, -7.132091e-15, -7.137428e-15, 
    -7.142113e-15, -7.153516e-15, -7.145639e-15, -7.148743e-15, 
    -7.141364e-15, -7.136677e-15, -7.138995e-15, -7.124708e-15, 
    -7.130258e-15, -7.101064e-15, -7.113622e-15, -7.080939e-15, 
    -7.088745e-15, -7.07907e-15, -7.084006e-15, -7.07555e-15, -7.08316e-15, 
    -7.069985e-15, -7.067119e-15, -7.069077e-15, -7.061562e-15, 
    -7.083582e-15, -7.075114e-15, -7.13906e-15, -7.138681e-15, -7.136921e-15, 
    -7.144661e-15, -7.145135e-15, -7.152241e-15, -7.14592e-15, -7.143229e-15, 
    -7.136407e-15, -7.132372e-15, -7.128541e-15, -7.120124e-15, 
    -7.110736e-15, -7.097633e-15, -7.088239e-15, -7.081949e-15, 
    -7.085806e-15, -7.0824e-15, -7.086207e-15, -7.087993e-15, -7.068191e-15, 
    -7.079301e-15, -7.062642e-15, -7.063563e-15, -7.071097e-15, 
    -7.063459e-15, -7.138416e-15, -7.140592e-15, -7.148148e-15, 
    -7.142234e-15, -7.153015e-15, -7.146977e-15, -7.143507e-15, 
    -7.130139e-15, -7.127209e-15, -7.124489e-15, -7.119124e-15, 
    -7.112243e-15, -7.100189e-15, -7.089722e-15, -7.080184e-15, 
    -7.080882e-15, -7.080636e-15, -7.078506e-15, -7.083783e-15, -7.07764e-15, 
    -7.076609e-15, -7.079304e-15, -7.063686e-15, -7.068144e-15, 
    -7.063583e-15, -7.066485e-15, -7.139885e-15, -7.136225e-15, 
    -7.138202e-15, -7.134484e-15, -7.137102e-15, -7.125464e-15, 
    -7.121978e-15, -7.105698e-15, -7.112377e-15, -7.101753e-15, 
    -7.111298e-15, -7.109606e-15, -7.101401e-15, -7.110783e-15, 
    -7.090296e-15, -7.104174e-15, -7.078423e-15, -7.09225e-15, -7.077557e-15, 
    -7.080225e-15, -7.07581e-15, -7.071858e-15, -7.066891e-15, -7.057733e-15, 
    -7.059853e-15, -7.052205e-15, -7.130773e-15, -7.126032e-15, 
    -7.126452e-15, -7.121495e-15, -7.117831e-15, -7.1099e-15, -7.097197e-15, 
    -7.101971e-15, -7.093211e-15, -7.091453e-15, -7.104765e-15, 
    -7.096586e-15, -7.122863e-15, -7.118607e-15, -7.121142e-15, 
    -7.130398e-15, -7.100867e-15, -7.116004e-15, -7.088084e-15, 
    -7.096263e-15, -7.072421e-15, -7.084264e-15, -7.06102e-15, -7.051103e-15, 
    -7.041797e-15, -7.030925e-15, -7.123448e-15, -7.126668e-15, 
    -7.120906e-15, -7.112939e-15, -7.105561e-15, -7.095764e-15, 
    -7.094763e-15, -7.092929e-15, -7.088183e-15, -7.084194e-15, 
    -7.092347e-15, -7.083194e-15, -7.117616e-15, -7.099556e-15, 
    -7.127884e-15, -7.119337e-15, -7.113409e-15, -7.116011e-15, 
    -7.102518e-15, -7.099341e-15, -7.086446e-15, -7.09311e-15, -7.053547e-15, 
    -7.07102e-15, -7.022669e-15, -7.03614e-15, -7.127793e-15, -7.123461e-15, 
    -7.108402e-15, -7.115563e-15, -7.095111e-15, -7.090086e-15, 
    -7.086006e-15, -7.08079e-15, -7.080229e-15, -7.077141e-15, -7.082202e-15, 
    -7.077342e-15, -7.095743e-15, -7.087513e-15, -7.110124e-15, 
    -7.104612e-15, -7.107149e-15, -7.109929e-15, -7.10135e-15, -7.092217e-15, 
    -7.092026e-15, -7.0891e-15, -7.080855e-15, -7.095029e-15, -7.051288e-15, 
    -7.078258e-15, -7.118739e-15, -7.110404e-15, -7.109219e-15, 
    -7.112445e-15, -7.090589e-15, -7.098499e-15, -7.077217e-15, 
    -7.082963e-15, -7.073552e-15, -7.078227e-15, -7.078914e-15, 
    -7.084924e-15, -7.088668e-15, -7.098136e-15, -7.105851e-15, 
    -7.111977e-15, -7.110553e-15, -7.103825e-15, -7.09166e-15, -7.080176e-15, 
    -7.08269e-15, -7.074267e-15, -7.096592e-15, -7.087219e-15, -7.090838e-15, 
    -7.081406e-15, -7.102097e-15, -7.084461e-15, -7.106612e-15, 
    -7.104668e-15, -7.098657e-15, -7.086581e-15, -7.083919e-15, -7.08107e-15, 
    -7.082828e-15, -7.091353e-15, -7.092752e-15, -7.098804e-15, 
    -7.100473e-15, -7.105091e-15, -7.108915e-15, -7.10542e-15, -7.101752e-15, 
    -7.091351e-15, -7.08199e-15, -7.071801e-15, -7.069312e-15, -7.057423e-15, 
    -7.067094e-15, -7.051138e-15, -7.064692e-15, -7.041252e-15, 
    -7.083446e-15, -7.065099e-15, -7.098385e-15, -7.094791e-15, 
    -7.088293e-15, -7.073422e-15, -7.08145e-15, -7.072064e-15, -7.092807e-15, 
    -7.103591e-15, -7.106389e-15, -7.111604e-15, -7.106269e-15, 
    -7.106704e-15, -7.101603e-15, -7.103242e-15, -7.091005e-15, 
    -7.097575e-15, -7.07893e-15, -7.072139e-15, -7.053004e-15, -7.041301e-15, 
    -7.029418e-15, -7.024178e-15, -7.022584e-15, -7.021918e-15 ;

 CH4_SURF_DIFF_UNSAT =
  1.652079e-14, 1.610252e-14, 1.618385e-14, 1.584641e-14, 1.603362e-14, 
    1.581264e-14, 1.643601e-14, 1.608591e-14, 1.630942e-14, 1.648316e-14, 
    1.519127e-14, 1.583136e-14, 1.452615e-14, 1.493461e-14, 1.390829e-14, 
    1.458971e-14, 1.377084e-14, 1.392798e-14, 1.345502e-14, 1.359054e-14, 
    1.298532e-14, 1.339247e-14, 1.26715e-14, 1.308258e-14, 1.301827e-14, 
    1.34059e-14, 1.570259e-14, 1.527097e-14, 1.572815e-14, 1.566662e-14, 
    1.569423e-14, 1.602974e-14, 1.619877e-14, 1.655277e-14, 1.648851e-14, 
    1.622851e-14, 1.563895e-14, 1.583912e-14, 1.533462e-14, 1.534601e-14, 
    1.47841e-14, 1.503748e-14, 1.409267e-14, 1.436129e-14, 1.358488e-14, 
    1.378019e-14, 1.359405e-14, 1.36505e-14, 1.359332e-14, 1.387975e-14, 
    1.375704e-14, 1.400905e-14, 1.499003e-14, 1.47018e-14, 1.556122e-14, 
    1.607767e-14, 1.642066e-14, 1.666397e-14, 1.662957e-14, 1.6564e-14, 
    1.622699e-14, 1.591009e-14, 1.566852e-14, 1.550691e-14, 1.534765e-14, 
    1.48654e-14, 1.461014e-14, 1.403834e-14, 1.414157e-14, 1.396669e-14, 
    1.379962e-14, 1.351904e-14, 1.356523e-14, 1.344159e-14, 1.397132e-14, 
    1.361928e-14, 1.420037e-14, 1.404147e-14, 1.530427e-14, 1.578513e-14, 
    1.598939e-14, 1.616822e-14, 1.660312e-14, 1.63028e-14, 1.642119e-14, 
    1.613952e-14, 1.59605e-14, 1.604904e-14, 1.550249e-14, 1.5715e-14, 
    1.459501e-14, 1.507755e-14, 1.381911e-14, 1.412039e-14, 1.374689e-14, 
    1.39375e-14, 1.361087e-14, 1.390484e-14, 1.339558e-14, 1.328465e-14, 
    1.336046e-14, 1.306926e-14, 1.392113e-14, 1.359405e-14, 1.605152e-14, 
    1.603708e-14, 1.596981e-14, 1.62655e-14, 1.628359e-14, 1.655453e-14, 
    1.631346e-14, 1.621078e-14, 1.595013e-14, 1.579591e-14, 1.56493e-14, 
    1.53269e-14, 1.496672e-14, 1.446292e-14, 1.410086e-14, 1.385808e-14, 
    1.400696e-14, 1.387552e-14, 1.402245e-14, 1.409132e-14, 1.332621e-14, 
    1.375589e-14, 1.311115e-14, 1.314684e-14, 1.343865e-14, 1.314282e-14, 
    1.602694e-14, 1.611004e-14, 1.63985e-14, 1.617276e-14, 1.658403e-14, 
    1.635383e-14, 1.622144e-14, 1.571054e-14, 1.559828e-14, 1.549416e-14, 
    1.52885e-14, 1.502452e-14, 1.456128e-14, 1.41581e-14, 1.37899e-14, 
    1.381689e-14, 1.380739e-14, 1.372511e-14, 1.392889e-14, 1.369165e-14, 
    1.365182e-14, 1.375595e-14, 1.315162e-14, 1.332431e-14, 1.31476e-14, 
    1.326004e-14, 1.608303e-14, 1.59432e-14, 1.601876e-14, 1.587667e-14, 
    1.597677e-14, 1.553158e-14, 1.539807e-14, 1.47732e-14, 1.502971e-14, 
    1.462147e-14, 1.498825e-14, 1.492327e-14, 1.460812e-14, 1.496844e-14, 
    1.418031e-14, 1.471466e-14, 1.372191e-14, 1.425572e-14, 1.368845e-14, 
    1.37915e-14, 1.362089e-14, 1.346806e-14, 1.327578e-14, 1.292087e-14, 
    1.300307e-14, 1.270621e-14, 1.573472e-14, 1.55533e-14, 1.556929e-14, 
    1.537941e-14, 1.523896e-14, 1.493452e-14, 1.444605e-14, 1.462977e-14, 
    1.42925e-14, 1.422477e-14, 1.473717e-14, 1.442258e-14, 1.543187e-14, 
    1.526884e-14, 1.536593e-14, 1.57204e-14, 1.458741e-14, 1.516898e-14, 
    1.409487e-14, 1.441009e-14, 1.348985e-14, 1.394759e-14, 1.304831e-14, 
    1.26636e-14, 1.230148e-14, 1.187803e-14, 1.545429e-14, 1.557757e-14, 
    1.535683e-14, 1.505133e-14, 1.476786e-14, 1.439086e-14, 1.435229e-14, 
    1.428165e-14, 1.409866e-14, 1.394476e-14, 1.425929e-14, 1.390618e-14, 
    1.5231e-14, 1.453693e-14, 1.562416e-14, 1.529685e-14, 1.506935e-14, 
    1.516917e-14, 1.465076e-14, 1.452854e-14, 1.403175e-14, 1.42886e-14, 
    1.275855e-14, 1.343575e-14, 1.155555e-14, 1.208133e-14, 1.562064e-14, 
    1.545472e-14, 1.487706e-14, 1.515195e-14, 1.43657e-14, 1.417208e-14, 
    1.401467e-14, 1.381338e-14, 1.379166e-14, 1.367238e-14, 1.386784e-14, 
    1.368011e-14, 1.439006e-14, 1.407287e-14, 1.494312e-14, 1.473136e-14, 
    1.482879e-14, 1.493564e-14, 1.460583e-14, 1.425434e-14, 1.424686e-14, 
    1.413412e-14, 1.381632e-14, 1.436252e-14, 1.267106e-14, 1.371594e-14, 
    1.527376e-14, 1.495403e-14, 1.490839e-14, 1.503225e-14, 1.41915e-14, 
    1.44962e-14, 1.36753e-14, 1.389723e-14, 1.353358e-14, 1.37143e-14, 
    1.374088e-14, 1.397294e-14, 1.411739e-14, 1.448222e-14, 1.477899e-14, 
    1.501429e-14, 1.495958e-14, 1.47011e-14, 1.423284e-14, 1.378968e-14, 
    1.388677e-14, 1.356122e-14, 1.442273e-14, 1.406156e-14, 1.420116e-14, 
    1.383712e-14, 1.463464e-14, 1.395547e-14, 1.480817e-14, 1.473344e-14, 
    1.450224e-14, 1.403704e-14, 1.393413e-14, 1.382418e-14, 1.389203e-14, 
    1.422096e-14, 1.427485e-14, 1.450787e-14, 1.457219e-14, 1.474971e-14, 
    1.489665e-14, 1.476239e-14, 1.462137e-14, 1.422083e-14, 1.385972e-14, 
    1.346588e-14, 1.336949e-14, 1.290904e-14, 1.328384e-14, 1.266524e-14, 
    1.319114e-14, 1.228063e-14, 1.391614e-14, 1.320665e-14, 1.449173e-14, 
    1.435337e-14, 1.410304e-14, 1.35287e-14, 1.383883e-14, 1.347614e-14, 
    1.427696e-14, 1.469217e-14, 1.479961e-14, 1.499998e-14, 1.479503e-14, 
    1.48117e-14, 1.461555e-14, 1.467859e-14, 1.420753e-14, 1.446058e-14, 
    1.374154e-14, 1.347901e-14, 1.273731e-14, 1.228235e-14, 1.181906e-14, 
    1.161444e-14, 1.155215e-14, 1.152611e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931951e-23, 1.931952e-23, 1.93195e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.93195e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.93195e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931946e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931946e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.931951e-23, 
    1.93195e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931943e-23, 1.931942e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 
    1.931944e-23, 1.931946e-23, 1.931942e-23, 1.931943e-23, 1.931951e-23, 
    1.931951e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.93195e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931944e-23, 
    1.931945e-23, 1.931943e-23, 1.931947e-23, 1.931946e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975384e-24, 1.975386e-24, 1.975381e-24, 1.975383e-24, 1.975379e-24, 
    1.975382e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975376e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 1.975377e-24, 
    1.975378e-24, 1.975385e-24, 1.975384e-24, 1.975385e-24, 1.975385e-24, 
    1.975385e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975386e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.975381e-24, 1.975378e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 1.975385e-24, 
    1.975387e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975383e-24, 1.975382e-24, 1.97538e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.97538e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975384e-24, 1.975386e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975382e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 
    1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975379e-24, 1.975386e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975377e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975382e-24, 1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975376e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975383e-24, 1.975381e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975382e-24, 1.975381e-24, 1.975384e-24, 
    1.975384e-24, 1.975384e-24, 1.975385e-24, 1.975382e-24, 1.975384e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 
    1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975384e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975384e-24, 1.975381e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975384e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.975376e-24, 1.975378e-24, 1.975372e-24, 1.975373e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975375e-24, 1.975379e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975382e-24, 1.97538e-24, 1.975382e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975378e-24, 1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975375e-24, 
    1.975377e-24, 1.975374e-24, 1.975379e-24, 1.975377e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24 ;

 CONC_CH4_SAT =
  3.275211e-08, 3.27318e-08, 3.273576e-08, 3.271936e-08, 3.272847e-08, 
    3.271772e-08, 3.274801e-08, 3.273098e-08, 3.274186e-08, 3.275031e-08, 
    3.268748e-08, 3.271863e-08, 3.265533e-08, 3.267515e-08, 3.262545e-08, 
    3.265839e-08, 3.261881e-08, 3.262644e-08, 3.26036e-08, 3.261014e-08, 
    3.258086e-08, 3.260058e-08, 3.256577e-08, 3.258559e-08, 3.258248e-08, 
    3.260122e-08, 3.27124e-08, 3.269135e-08, 3.271364e-08, 3.271063e-08, 
    3.271199e-08, 3.272827e-08, 3.273644e-08, 3.275369e-08, 3.275057e-08, 
    3.273791e-08, 3.270929e-08, 3.271903e-08, 3.269456e-08, 3.269511e-08, 
    3.266786e-08, 3.268014e-08, 3.26344e-08, 3.26474e-08, 3.260987e-08, 
    3.26193e-08, 3.261031e-08, 3.261304e-08, 3.261027e-08, 3.26241e-08, 
    3.261817e-08, 3.263036e-08, 3.267783e-08, 3.266386e-08, 3.270553e-08, 
    3.273054e-08, 3.274726e-08, 3.275909e-08, 3.275742e-08, 3.275422e-08, 
    3.273784e-08, 3.272248e-08, 3.271075e-08, 3.270291e-08, 3.269519e-08, 
    3.267172e-08, 3.26594e-08, 3.263175e-08, 3.263677e-08, 3.262829e-08, 
    3.262024e-08, 3.260668e-08, 3.260892e-08, 3.260293e-08, 3.262854e-08, 
    3.261151e-08, 3.263963e-08, 3.263193e-08, 3.269295e-08, 3.271641e-08, 
    3.272626e-08, 3.273499e-08, 3.275613e-08, 3.274152e-08, 3.274728e-08, 
    3.273362e-08, 3.272492e-08, 3.272923e-08, 3.27027e-08, 3.2713e-08, 
    3.265867e-08, 3.268206e-08, 3.262118e-08, 3.263574e-08, 3.261769e-08, 
    3.262691e-08, 3.261111e-08, 3.262533e-08, 3.260072e-08, 3.259535e-08, 
    3.259902e-08, 3.258498e-08, 3.262612e-08, 3.261029e-08, 3.272934e-08, 
    3.272864e-08, 3.272538e-08, 3.273971e-08, 3.274059e-08, 3.275377e-08, 
    3.274206e-08, 3.273706e-08, 3.272443e-08, 3.271693e-08, 3.270981e-08, 
    3.269417e-08, 3.267668e-08, 3.265229e-08, 3.26348e-08, 3.262307e-08, 
    3.263027e-08, 3.262391e-08, 3.263101e-08, 3.263435e-08, 3.259735e-08, 
    3.261811e-08, 3.2587e-08, 3.258872e-08, 3.260279e-08, 3.258853e-08, 
    3.272815e-08, 3.273219e-08, 3.274619e-08, 3.273523e-08, 3.275521e-08, 
    3.274401e-08, 3.273756e-08, 3.271276e-08, 3.270734e-08, 3.270228e-08, 
    3.269231e-08, 3.267951e-08, 3.265706e-08, 3.263755e-08, 3.261978e-08, 
    3.262108e-08, 3.262062e-08, 3.261664e-08, 3.262649e-08, 3.261502e-08, 
    3.261308e-08, 3.261813e-08, 3.258895e-08, 3.259728e-08, 3.258876e-08, 
    3.259419e-08, 3.273088e-08, 3.272408e-08, 3.272775e-08, 3.272084e-08, 
    3.27257e-08, 3.270407e-08, 3.269758e-08, 3.266729e-08, 3.267976e-08, 
    3.265997e-08, 3.267776e-08, 3.26746e-08, 3.265926e-08, 3.267681e-08, 
    3.26386e-08, 3.266445e-08, 3.261648e-08, 3.264222e-08, 3.261487e-08, 
    3.261985e-08, 3.261161e-08, 3.260422e-08, 3.259494e-08, 3.257779e-08, 
    3.258177e-08, 3.256746e-08, 3.271396e-08, 3.270514e-08, 3.270594e-08, 
    3.269672e-08, 3.26899e-08, 3.267516e-08, 3.265149e-08, 3.26604e-08, 
    3.264408e-08, 3.264079e-08, 3.26656e-08, 3.265034e-08, 3.269925e-08, 
    3.269132e-08, 3.269606e-08, 3.271325e-08, 3.265831e-08, 3.268648e-08, 
    3.26345e-08, 3.264975e-08, 3.260527e-08, 3.262736e-08, 3.258395e-08, 
    3.256535e-08, 3.254797e-08, 3.252753e-08, 3.270035e-08, 3.270634e-08, 
    3.269563e-08, 3.268078e-08, 3.266707e-08, 3.264882e-08, 3.264697e-08, 
    3.264354e-08, 3.26347e-08, 3.262726e-08, 3.264244e-08, 3.262539e-08, 
    3.268942e-08, 3.265588e-08, 3.270858e-08, 3.269267e-08, 3.268167e-08, 
    3.268652e-08, 3.266142e-08, 3.26555e-08, 3.263144e-08, 3.264389e-08, 
    3.256991e-08, 3.260262e-08, 3.251207e-08, 3.253733e-08, 3.270843e-08, 
    3.270038e-08, 3.267235e-08, 3.268569e-08, 3.264762e-08, 3.263824e-08, 
    3.263064e-08, 3.262089e-08, 3.261986e-08, 3.261409e-08, 3.262354e-08, 
    3.261447e-08, 3.264878e-08, 3.263345e-08, 3.267558e-08, 3.266531e-08, 
    3.267004e-08, 3.267522e-08, 3.265924e-08, 3.264219e-08, 3.264187e-08, 
    3.263639e-08, 3.26209e-08, 3.264746e-08, 3.256562e-08, 3.261607e-08, 
    3.269161e-08, 3.267606e-08, 3.267388e-08, 3.26799e-08, 3.263918e-08, 
    3.265392e-08, 3.261423e-08, 3.262496e-08, 3.260739e-08, 3.261612e-08, 
    3.26174e-08, 3.262862e-08, 3.26356e-08, 3.265324e-08, 3.266761e-08, 
    3.267903e-08, 3.267638e-08, 3.266383e-08, 3.264116e-08, 3.261975e-08, 
    3.262443e-08, 3.260873e-08, 3.265037e-08, 3.263288e-08, 3.263963e-08, 
    3.262205e-08, 3.266062e-08, 3.262765e-08, 3.266904e-08, 3.266542e-08, 
    3.265421e-08, 3.263167e-08, 3.262674e-08, 3.262141e-08, 3.262471e-08, 
    3.264059e-08, 3.264321e-08, 3.26545e-08, 3.26576e-08, 3.266621e-08, 
    3.267333e-08, 3.266682e-08, 3.265997e-08, 3.26406e-08, 3.262313e-08, 
    3.260411e-08, 3.259947e-08, 3.257716e-08, 3.259526e-08, 3.256533e-08, 
    3.259069e-08, 3.254685e-08, 3.26258e-08, 3.259152e-08, 3.265372e-08, 
    3.264702e-08, 3.263487e-08, 3.26071e-08, 3.262213e-08, 3.260458e-08, 
    3.264331e-08, 3.266338e-08, 3.266863e-08, 3.267833e-08, 3.26684e-08, 
    3.266921e-08, 3.265972e-08, 3.266277e-08, 3.263996e-08, 3.265221e-08, 
    3.261742e-08, 3.260472e-08, 3.256894e-08, 3.2547e-08, 3.252476e-08, 
    3.251492e-08, 3.251193e-08, 3.251068e-08,
  5.417225e-11, 5.419688e-11, 5.419213e-11, 5.4212e-11, 5.420099e-11, 
    5.42145e-11, 5.417732e-11, 5.419779e-11, 5.418476e-11, 5.417457e-11, 
    5.425991e-11, 5.421313e-11, 5.430903e-11, 5.42792e-11, 5.435422e-11, 
    5.430429e-11, 5.436429e-11, 5.435294e-11, 5.438746e-11, 5.437759e-11, 
    5.442129e-11, 5.439201e-11, 5.444416e-11, 5.44144e-11, 5.441899e-11, 
    5.439102e-11, 5.422271e-11, 5.425405e-11, 5.422082e-11, 5.42253e-11, 
    5.422332e-11, 5.420116e-11, 5.419109e-11, 5.417048e-11, 5.417425e-11, 
    5.418945e-11, 5.422732e-11, 5.421266e-11, 5.424988e-11, 5.424905e-11, 
    5.429027e-11, 5.427169e-11, 5.434091e-11, 5.432131e-11, 5.437801e-11, 
    5.436375e-11, 5.43773e-11, 5.437322e-11, 5.437736e-11, 5.435645e-11, 
    5.43654e-11, 5.434704e-11, 5.427514e-11, 5.429626e-11, 5.42331e-11, 
    5.419812e-11, 5.417819e-11, 5.416391e-11, 5.416593e-11, 5.416975e-11, 
    5.418953e-11, 5.420826e-11, 5.422528e-11, 5.423718e-11, 5.424892e-11, 
    5.428399e-11, 5.430287e-11, 5.434479e-11, 5.433737e-11, 5.435005e-11, 
    5.436233e-11, 5.438275e-11, 5.437941e-11, 5.438837e-11, 5.434981e-11, 
    5.43754e-11, 5.433312e-11, 5.434468e-11, 5.425157e-11, 5.421665e-11, 
    5.420334e-11, 5.419302e-11, 5.416747e-11, 5.418509e-11, 5.417813e-11, 
    5.419479e-11, 5.420529e-11, 5.420012e-11, 5.423751e-11, 5.422182e-11, 
    5.430399e-11, 5.426866e-11, 5.43609e-11, 5.433891e-11, 5.436619e-11, 
    5.43523e-11, 5.437604e-11, 5.435468e-11, 5.439174e-11, 5.439974e-11, 
    5.439426e-11, 5.441547e-11, 5.435348e-11, 5.437725e-11, 5.419995e-11, 
    5.420079e-11, 5.420477e-11, 5.418727e-11, 5.418623e-11, 5.417035e-11, 
    5.418453e-11, 5.419052e-11, 5.420594e-11, 5.421584e-11, 5.422665e-11, 
    5.42504e-11, 5.427678e-11, 5.431374e-11, 5.434033e-11, 5.435809e-11, 
    5.434724e-11, 5.435682e-11, 5.434609e-11, 5.434108e-11, 5.439671e-11, 
    5.436545e-11, 5.441242e-11, 5.440984e-11, 5.438856e-11, 5.441014e-11, 
    5.420139e-11, 5.419654e-11, 5.417951e-11, 5.419284e-11, 5.416862e-11, 
    5.418211e-11, 5.418983e-11, 5.422203e-11, 5.423045e-11, 5.423807e-11, 
    5.425325e-11, 5.427264e-11, 5.430656e-11, 5.433609e-11, 5.436307e-11, 
    5.436111e-11, 5.436179e-11, 5.436776e-11, 5.43529e-11, 5.43702e-11, 
    5.437304e-11, 5.436552e-11, 5.440949e-11, 5.439695e-11, 5.440979e-11, 
    5.440164e-11, 5.419813e-11, 5.420632e-11, 5.420189e-11, 5.421019e-11, 
    5.420429e-11, 5.423519e-11, 5.424499e-11, 5.429092e-11, 5.427223e-11, 
    5.430212e-11, 5.427531e-11, 5.428004e-11, 5.430286e-11, 5.42768e-11, 
    5.433436e-11, 5.429515e-11, 5.436799e-11, 5.432872e-11, 5.437043e-11, 
    5.436295e-11, 5.437539e-11, 5.438646e-11, 5.440047e-11, 5.442613e-11, 
    5.442021e-11, 5.444174e-11, 5.422037e-11, 5.423366e-11, 5.423259e-11, 
    5.424656e-11, 5.425686e-11, 5.427928e-11, 5.431505e-11, 5.430164e-11, 
    5.432636e-11, 5.433128e-11, 5.429378e-11, 5.431672e-11, 5.424262e-11, 
    5.425451e-11, 5.424751e-11, 5.422136e-11, 5.430459e-11, 5.426187e-11, 
    5.434075e-11, 5.431771e-11, 5.438486e-11, 5.43514e-11, 5.441693e-11, 
    5.444458e-11, 5.447104e-11, 5.450132e-11, 5.424102e-11, 5.423199e-11, 
    5.424825e-11, 5.427053e-11, 5.429147e-11, 5.431909e-11, 5.432197e-11, 
    5.432711e-11, 5.434054e-11, 5.435176e-11, 5.432864e-11, 5.435459e-11, 
    5.425706e-11, 5.430834e-11, 5.422847e-11, 5.425243e-11, 5.426927e-11, 
    5.426199e-11, 5.430013e-11, 5.430907e-11, 5.43453e-11, 5.432665e-11, 
    5.443767e-11, 5.438865e-11, 5.452468e-11, 5.448673e-11, 5.42288e-11, 
    5.424104e-11, 5.428339e-11, 5.426327e-11, 5.432099e-11, 5.433512e-11, 
    5.434668e-11, 5.436127e-11, 5.436292e-11, 5.437158e-11, 5.435738e-11, 
    5.437106e-11, 5.431915e-11, 5.434239e-11, 5.427868e-11, 5.429415e-11, 
    5.428707e-11, 5.427922e-11, 5.430341e-11, 5.432898e-11, 5.432969e-11, 
    5.433784e-11, 5.43605e-11, 5.432123e-11, 5.444367e-11, 5.436789e-11, 
    5.425435e-11, 5.427764e-11, 5.428117e-11, 5.427212e-11, 5.43337e-11, 
    5.431139e-11, 5.437139e-11, 5.435524e-11, 5.438174e-11, 5.436856e-11, 
    5.436661e-11, 5.434971e-11, 5.433913e-11, 5.431238e-11, 5.429064e-11, 
    5.427345e-11, 5.427746e-11, 5.429634e-11, 5.433057e-11, 5.4363e-11, 
    5.435588e-11, 5.437972e-11, 5.431681e-11, 5.434314e-11, 5.433291e-11, 
    5.435959e-11, 5.430125e-11, 5.435044e-11, 5.428858e-11, 5.429406e-11, 
    5.431095e-11, 5.434481e-11, 5.435254e-11, 5.436048e-11, 5.435562e-11, 
    5.433147e-11, 5.432759e-11, 5.431058e-11, 5.43058e-11, 5.429288e-11, 
    5.428209e-11, 5.42919e-11, 5.430217e-11, 5.433155e-11, 5.435788e-11, 
    5.438659e-11, 5.439367e-11, 5.44267e-11, 5.439959e-11, 5.444406e-11, 
    5.440591e-11, 5.447206e-11, 5.435353e-11, 5.440513e-11, 5.431178e-11, 
    5.432191e-11, 5.434003e-11, 5.438186e-11, 5.435947e-11, 5.438573e-11, 
    5.432745e-11, 5.42969e-11, 5.42892e-11, 5.427447e-11, 5.428953e-11, 
    5.428832e-11, 5.430271e-11, 5.42981e-11, 5.433253e-11, 5.431405e-11, 
    5.436652e-11, 5.438556e-11, 5.443942e-11, 5.447223e-11, 5.450581e-11, 
    5.452051e-11, 5.4525e-11, 5.452687e-11,
  2.415998e-14, 2.419375e-14, 2.418721e-14, 2.421624e-14, 2.419936e-14, 
    2.421962e-14, 2.416687e-14, 2.419505e-14, 2.417709e-14, 2.416309e-14, 
    2.428143e-14, 2.421775e-14, 2.434811e-14, 2.430739e-14, 2.440986e-14, 
    2.43417e-14, 2.442363e-14, 2.440802e-14, 2.44553e-14, 2.444176e-14, 
    2.450202e-14, 2.446156e-14, 2.453346e-14, 2.449242e-14, 2.449879e-14, 
    2.44602e-14, 2.423068e-14, 2.427346e-14, 2.422812e-14, 2.423422e-14, 
    2.423151e-14, 2.419963e-14, 2.418589e-14, 2.415748e-14, 2.416265e-14, 
    2.418356e-14, 2.423697e-14, 2.421706e-14, 2.426748e-14, 2.426635e-14, 
    2.432244e-14, 2.429714e-14, 2.439156e-14, 2.436474e-14, 2.444233e-14, 
    2.44228e-14, 2.444139e-14, 2.443577e-14, 2.444147e-14, 2.441283e-14, 
    2.442509e-14, 2.439993e-14, 2.430186e-14, 2.433063e-14, 2.424477e-14, 
    2.41956e-14, 2.416809e-14, 2.41485e-14, 2.415126e-14, 2.415652e-14, 
    2.418368e-14, 2.421045e-14, 2.423412e-14, 2.425026e-14, 2.426618e-14, 
    2.431409e-14, 2.433972e-14, 2.439692e-14, 2.43867e-14, 2.440409e-14, 
    2.442086e-14, 2.444887e-14, 2.444428e-14, 2.44566e-14, 2.440371e-14, 
    2.443882e-14, 2.438085e-14, 2.439669e-14, 2.427011e-14, 2.422245e-14, 
    2.420304e-14, 2.418845e-14, 2.415339e-14, 2.417757e-14, 2.416803e-14, 
    2.419083e-14, 2.420585e-14, 2.419814e-14, 2.42507e-14, 2.422946e-14, 
    2.434123e-14, 2.429307e-14, 2.44189e-14, 2.43888e-14, 2.442613e-14, 
    2.44071e-14, 2.443968e-14, 2.441036e-14, 2.446122e-14, 2.447225e-14, 
    2.44647e-14, 2.449383e-14, 2.440873e-14, 2.444135e-14, 2.419792e-14, 
    2.419908e-14, 2.420502e-14, 2.418058e-14, 2.417913e-14, 2.415732e-14, 
    2.417676e-14, 2.418502e-14, 2.420683e-14, 2.422136e-14, 2.423601e-14, 
    2.426821e-14, 2.430413e-14, 2.435449e-14, 2.439075e-14, 2.441504e-14, 
    2.440017e-14, 2.441329e-14, 2.439861e-14, 2.439175e-14, 2.446809e-14, 
    2.442518e-14, 2.448964e-14, 2.448608e-14, 2.445688e-14, 2.448648e-14, 
    2.41999e-14, 2.419322e-14, 2.416989e-14, 2.418815e-14, 2.415495e-14, 
    2.417347e-14, 2.418411e-14, 2.422981e-14, 2.424113e-14, 2.42515e-14, 
    2.427207e-14, 2.429843e-14, 2.434468e-14, 2.438499e-14, 2.442185e-14, 
    2.441916e-14, 2.44201e-14, 2.44283e-14, 2.440795e-14, 2.443164e-14, 
    2.443558e-14, 2.442522e-14, 2.44856e-14, 2.446836e-14, 2.448601e-14, 
    2.447478e-14, 2.41954e-14, 2.420743e-14, 2.420057e-14, 2.421347e-14, 
    2.420434e-14, 2.424767e-14, 2.426098e-14, 2.432343e-14, 2.429789e-14, 
    2.433864e-14, 2.430206e-14, 2.430852e-14, 2.43398e-14, 2.430407e-14, 
    2.438269e-14, 2.432923e-14, 2.442862e-14, 2.437506e-14, 2.443196e-14, 
    2.442169e-14, 2.443874e-14, 2.445396e-14, 2.44732e-14, 2.450857e-14, 
    2.45004e-14, 2.453005e-14, 2.422749e-14, 2.424555e-14, 2.424403e-14, 
    2.426299e-14, 2.427699e-14, 2.430745e-14, 2.435623e-14, 2.43379e-14, 
    2.437163e-14, 2.437837e-14, 2.432719e-14, 2.435854e-14, 2.425769e-14, 
    2.42739e-14, 2.426431e-14, 2.422887e-14, 2.434202e-14, 2.428389e-14, 
    2.439134e-14, 2.435984e-14, 2.445178e-14, 2.440598e-14, 2.449588e-14, 
    2.453413e-14, 2.45705e-14, 2.461259e-14, 2.425549e-14, 2.424321e-14, 
    2.426526e-14, 2.429565e-14, 2.432407e-14, 2.436175e-14, 2.436564e-14, 
    2.437268e-14, 2.439101e-14, 2.440637e-14, 2.437483e-14, 2.441023e-14, 
    2.427751e-14, 2.43471e-14, 2.423849e-14, 2.427109e-14, 2.429389e-14, 
    2.428397e-14, 2.433583e-14, 2.434803e-14, 2.43976e-14, 2.437202e-14, 
    2.452462e-14, 2.445708e-14, 2.464491e-14, 2.459234e-14, 2.42389e-14, 
    2.425548e-14, 2.431311e-14, 2.42857e-14, 2.43643e-14, 2.438363e-14, 
    2.43994e-14, 2.441944e-14, 2.442166e-14, 2.443355e-14, 2.441406e-14, 
    2.443281e-14, 2.436183e-14, 2.439356e-14, 2.430661e-14, 2.432772e-14, 
    2.431803e-14, 2.430735e-14, 2.434031e-14, 2.437531e-14, 2.437618e-14, 
    2.438738e-14, 2.441874e-14, 2.436462e-14, 2.453312e-14, 2.442883e-14, 
    2.427356e-14, 2.430535e-14, 2.431004e-14, 2.42977e-14, 2.438169e-14, 
    2.435123e-14, 2.443328e-14, 2.441113e-14, 2.444745e-14, 2.442939e-14, 
    2.442672e-14, 2.440356e-14, 2.43891e-14, 2.43526e-14, 2.432295e-14, 
    2.42995e-14, 2.430496e-14, 2.433072e-14, 2.437748e-14, 2.442181e-14, 
    2.441208e-14, 2.444469e-14, 2.43586e-14, 2.439463e-14, 2.438066e-14, 
    2.441711e-14, 2.433739e-14, 2.440491e-14, 2.43201e-14, 2.432756e-14, 
    2.435063e-14, 2.4397e-14, 2.440744e-14, 2.441836e-14, 2.441165e-14, 
    2.437869e-14, 2.437335e-14, 2.435009e-14, 2.434362e-14, 2.432594e-14, 
    2.431125e-14, 2.432464e-14, 2.433868e-14, 2.437876e-14, 2.441481e-14, 
    2.445416e-14, 2.446384e-14, 2.450954e-14, 2.447217e-14, 2.453368e-14, 
    2.448113e-14, 2.457223e-14, 2.4409e-14, 2.447983e-14, 2.435172e-14, 
    2.436554e-14, 2.439043e-14, 2.444777e-14, 2.441694e-14, 2.445306e-14, 
    2.437315e-14, 2.433155e-14, 2.432094e-14, 2.43009e-14, 2.43214e-14, 
    2.431974e-14, 2.433935e-14, 2.433305e-14, 2.438009e-14, 2.435482e-14, 
    2.442663e-14, 2.44528e-14, 2.45269e-14, 2.457227e-14, 2.461866e-14, 
    2.463908e-14, 2.464531e-14, 2.46479e-14,
  3.207574e-18, 3.214927e-18, 3.213501e-18, 3.219791e-18, 3.216147e-18, 
    3.220486e-18, 3.209072e-18, 3.215211e-18, 3.211295e-18, 3.208247e-18, 
    3.233226e-18, 3.220102e-18, 3.246986e-18, 3.23857e-18, 3.259766e-18, 
    3.245663e-18, 3.262618e-18, 3.259379e-18, 3.269185e-18, 3.266375e-18, 
    3.279338e-18, 3.270483e-18, 3.28629e-18, 3.27721e-18, 3.278622e-18, 
    3.270202e-18, 3.222759e-18, 3.231584e-18, 3.222233e-18, 3.223491e-18, 
    3.222931e-18, 3.216208e-18, 3.213218e-18, 3.207026e-18, 3.208153e-18, 
    3.212708e-18, 3.224057e-18, 3.219956e-18, 3.230338e-18, 3.230104e-18, 
    3.241678e-18, 3.236455e-18, 3.25597e-18, 3.250419e-18, 3.266492e-18, 
    3.262442e-18, 3.266299e-18, 3.265131e-18, 3.266314e-18, 3.260376e-18, 
    3.262918e-18, 3.257704e-18, 3.237429e-18, 3.243371e-18, 3.225662e-18, 
    3.215337e-18, 3.209337e-18, 3.205073e-18, 3.205675e-18, 3.20682e-18, 
    3.212735e-18, 3.218545e-18, 3.223466e-18, 3.22679e-18, 3.23007e-18, 
    3.239962e-18, 3.245251e-18, 3.257083e-18, 3.254963e-18, 3.258569e-18, 
    3.26204e-18, 3.267851e-18, 3.266897e-18, 3.269455e-18, 3.258486e-18, 
    3.265767e-18, 3.253752e-18, 3.257033e-18, 3.230894e-18, 3.221065e-18, 
    3.216952e-18, 3.213772e-18, 3.206137e-18, 3.211404e-18, 3.209325e-18, 
    3.214287e-18, 3.217552e-18, 3.215881e-18, 3.226881e-18, 3.222507e-18, 
    3.245564e-18, 3.235618e-18, 3.261635e-18, 3.2554e-18, 3.263134e-18, 
    3.259189e-18, 3.265945e-18, 3.259864e-18, 3.270413e-18, 3.272752e-18, 
    3.271137e-18, 3.277518e-18, 3.259526e-18, 3.266292e-18, 3.215834e-18, 
    3.216087e-18, 3.217372e-18, 3.212058e-18, 3.211743e-18, 3.206992e-18, 
    3.211225e-18, 3.213024e-18, 3.217762e-18, 3.220843e-18, 3.223856e-18, 
    3.23049e-18, 3.2379e-18, 3.248303e-18, 3.255803e-18, 3.260833e-18, 
    3.257753e-18, 3.260471e-18, 3.257429e-18, 3.256007e-18, 3.271842e-18, 
    3.262938e-18, 3.276592e-18, 3.275806e-18, 3.269513e-18, 3.275895e-18, 
    3.216266e-18, 3.214808e-18, 3.209729e-18, 3.213703e-18, 3.206475e-18, 
    3.21051e-18, 3.212828e-18, 3.222584e-18, 3.22491e-18, 3.227046e-18, 
    3.231284e-18, 3.236722e-18, 3.246273e-18, 3.254612e-18, 3.262245e-18, 
    3.261687e-18, 3.261883e-18, 3.263583e-18, 3.259364e-18, 3.264276e-18, 
    3.265095e-18, 3.262945e-18, 3.2757e-18, 3.271895e-18, 3.275789e-18, 
    3.273309e-18, 3.215284e-18, 3.217894e-18, 3.216412e-18, 3.219199e-18, 
    3.217227e-18, 3.226261e-18, 3.229004e-18, 3.241885e-18, 3.236611e-18, 
    3.245027e-18, 3.23747e-18, 3.238804e-18, 3.245273e-18, 3.237883e-18, 
    3.254138e-18, 3.243085e-18, 3.263649e-18, 3.252562e-18, 3.264343e-18, 
    3.262212e-18, 3.265747e-18, 3.268908e-18, 3.272959e-18, 3.280782e-18, 
    3.278972e-18, 3.285533e-18, 3.222103e-18, 3.225822e-18, 3.225507e-18, 
    3.229413e-18, 3.2323e-18, 3.238581e-18, 3.24866e-18, 3.244871e-18, 
    3.251843e-18, 3.25324e-18, 3.242656e-18, 3.249139e-18, 3.228323e-18, 
    3.231666e-18, 3.229685e-18, 3.222388e-18, 3.245726e-18, 3.233725e-18, 
    3.255925e-18, 3.249406e-18, 3.268456e-18, 3.258959e-18, 3.277973e-18, 
    3.286445e-18, 3.294492e-18, 3.303841e-18, 3.227868e-18, 3.225337e-18, 
    3.229881e-18, 3.236151e-18, 3.242014e-18, 3.249801e-18, 3.250606e-18, 
    3.252063e-18, 3.255854e-18, 3.259038e-18, 3.252511e-18, 3.259837e-18, 
    3.232416e-18, 3.246776e-18, 3.224369e-18, 3.231086e-18, 3.235787e-18, 
    3.233737e-18, 3.244442e-18, 3.246964e-18, 3.257223e-18, 3.251924e-18, 
    3.284342e-18, 3.269558e-18, 3.311015e-18, 3.299344e-18, 3.22445e-18, 
    3.227865e-18, 3.239753e-18, 3.234094e-18, 3.250328e-18, 3.254328e-18, 
    3.257593e-18, 3.261748e-18, 3.262206e-18, 3.264672e-18, 3.260631e-18, 
    3.264518e-18, 3.249818e-18, 3.256384e-18, 3.238407e-18, 3.242768e-18, 
    3.240766e-18, 3.238561e-18, 3.245368e-18, 3.25261e-18, 3.252786e-18, 
    3.255107e-18, 3.261617e-18, 3.250395e-18, 3.286234e-18, 3.263706e-18, 
    3.231591e-18, 3.238153e-18, 3.239117e-18, 3.236568e-18, 3.253926e-18, 
    3.247626e-18, 3.264615e-18, 3.260022e-18, 3.267555e-18, 3.263809e-18, 
    3.263256e-18, 3.258454e-18, 3.255462e-18, 3.247911e-18, 3.241783e-18, 
    3.23694e-18, 3.238067e-18, 3.243389e-18, 3.253059e-18, 3.262239e-18, 
    3.260223e-18, 3.266983e-18, 3.249148e-18, 3.256608e-18, 3.253717e-18, 
    3.261263e-18, 3.244766e-18, 3.258748e-18, 3.241192e-18, 3.242733e-18, 
    3.247501e-18, 3.257101e-18, 3.259258e-18, 3.261525e-18, 3.26013e-18, 
    3.253308e-18, 3.252201e-18, 3.24739e-18, 3.246053e-18, 3.242399e-18, 
    3.239366e-18, 3.242132e-18, 3.245034e-18, 3.25332e-18, 3.260787e-18, 
    3.26895e-18, 3.270958e-18, 3.281007e-18, 3.272743e-18, 3.286358e-18, 
    3.274737e-18, 3.294893e-18, 3.25959e-18, 3.274438e-18, 3.247725e-18, 
    3.250585e-18, 3.25574e-18, 3.267627e-18, 3.261228e-18, 3.268723e-18, 
    3.252159e-18, 3.243562e-18, 3.241367e-18, 3.237231e-18, 3.241461e-18, 
    3.241118e-18, 3.245169e-18, 3.243868e-18, 3.253595e-18, 3.248368e-18, 
    3.263237e-18, 3.268669e-18, 3.284838e-18, 3.294892e-18, 3.30518e-18, 
    3.309717e-18, 3.311101e-18, 3.311678e-18,
  1.341941e-22, 1.346684e-22, 1.345763e-22, 1.349729e-22, 1.347471e-22, 
    1.350149e-22, 1.342905e-22, 1.346869e-22, 1.34434e-22, 1.342373e-22, 
    1.357853e-22, 1.349917e-22, 1.36618e-22, 1.36108e-22, 1.373933e-22, 
    1.365379e-22, 1.375665e-22, 1.373695e-22, 1.379674e-22, 1.377945e-22, 
    1.386118e-22, 1.380494e-22, 1.390534e-22, 1.384763e-22, 1.385661e-22, 
    1.380317e-22, 1.35152e-22, 1.35686e-22, 1.351202e-22, 1.351963e-22, 
    1.351623e-22, 1.347511e-22, 1.345584e-22, 1.341585e-22, 1.342312e-22, 
    1.345253e-22, 1.352305e-22, 1.349827e-22, 1.356098e-22, 1.355957e-22, 
    1.362961e-22, 1.359799e-22, 1.371626e-22, 1.368258e-22, 1.378016e-22, 
    1.375555e-22, 1.377899e-22, 1.377189e-22, 1.377908e-22, 1.374301e-22, 
    1.375845e-22, 1.372678e-22, 1.360389e-22, 1.363988e-22, 1.353274e-22, 
    1.346954e-22, 1.343077e-22, 1.340326e-22, 1.340715e-22, 1.341454e-22, 
    1.34527e-22, 1.34896e-22, 1.351946e-22, 1.353954e-22, 1.355936e-22, 
    1.361927e-22, 1.365128e-22, 1.372303e-22, 1.371014e-22, 1.373204e-22, 
    1.375311e-22, 1.378843e-22, 1.378263e-22, 1.379846e-22, 1.373153e-22, 
    1.377577e-22, 1.370278e-22, 1.37227e-22, 1.356443e-22, 1.350496e-22, 
    1.347981e-22, 1.345939e-22, 1.341013e-22, 1.344411e-22, 1.34307e-22, 
    1.34627e-22, 1.348347e-22, 1.347298e-22, 1.354009e-22, 1.351367e-22, 
    1.365318e-22, 1.359294e-22, 1.375065e-22, 1.371279e-22, 1.375975e-22, 
    1.373579e-22, 1.377684e-22, 1.373989e-22, 1.380451e-22, 1.381933e-22, 
    1.380909e-22, 1.384956e-22, 1.373784e-22, 1.377896e-22, 1.347268e-22, 
    1.347432e-22, 1.348235e-22, 1.344833e-22, 1.34463e-22, 1.341564e-22, 
    1.344294e-22, 1.345456e-22, 1.348475e-22, 1.350362e-22, 1.352182e-22, 
    1.356191e-22, 1.360675e-22, 1.366977e-22, 1.371524e-22, 1.374577e-22, 
    1.372707e-22, 1.374358e-22, 1.372511e-22, 1.371647e-22, 1.381356e-22, 
    1.375857e-22, 1.384369e-22, 1.383869e-22, 1.379883e-22, 1.383926e-22, 
    1.347547e-22, 1.346605e-22, 1.343329e-22, 1.345892e-22, 1.341231e-22, 
    1.343834e-22, 1.345331e-22, 1.351415e-22, 1.352818e-22, 1.354109e-22, 
    1.356671e-22, 1.359961e-22, 1.365746e-22, 1.370802e-22, 1.375435e-22, 
    1.375096e-22, 1.375215e-22, 1.376248e-22, 1.373686e-22, 1.37667e-22, 
    1.377168e-22, 1.375861e-22, 1.383802e-22, 1.381387e-22, 1.383859e-22, 
    1.382284e-22, 1.346912e-22, 1.348557e-22, 1.347641e-22, 1.349364e-22, 
    1.348147e-22, 1.353637e-22, 1.355295e-22, 1.363089e-22, 1.359894e-22, 
    1.364991e-22, 1.360414e-22, 1.361222e-22, 1.365144e-22, 1.360663e-22, 
    1.370517e-22, 1.363817e-22, 1.376289e-22, 1.369563e-22, 1.37671e-22, 
    1.375415e-22, 1.377563e-22, 1.3795e-22, 1.382062e-22, 1.387032e-22, 
    1.385882e-22, 1.390051e-22, 1.351123e-22, 1.353371e-22, 1.353179e-22, 
    1.355539e-22, 1.357286e-22, 1.361086e-22, 1.367192e-22, 1.364895e-22, 
    1.369121e-22, 1.369969e-22, 1.363553e-22, 1.367483e-22, 1.354882e-22, 
    1.356905e-22, 1.355705e-22, 1.351296e-22, 1.365416e-22, 1.35815e-22, 
    1.371598e-22, 1.367644e-22, 1.379214e-22, 1.373442e-22, 1.385247e-22, 
    1.390636e-22, 1.395751e-22, 1.401713e-22, 1.354606e-22, 1.353076e-22, 
    1.355822e-22, 1.359618e-22, 1.363165e-22, 1.367884e-22, 1.368371e-22, 
    1.369255e-22, 1.371555e-22, 1.373487e-22, 1.369529e-22, 1.373973e-22, 
    1.357362e-22, 1.366051e-22, 1.352492e-22, 1.356555e-22, 1.359396e-22, 
    1.358155e-22, 1.364634e-22, 1.366163e-22, 1.372388e-22, 1.36917e-22, 
    1.389299e-22, 1.379914e-22, 1.406287e-22, 1.398845e-22, 1.35254e-22, 
    1.354604e-22, 1.361797e-22, 1.358371e-22, 1.368203e-22, 1.370629e-22, 
    1.37261e-22, 1.375135e-22, 1.375412e-22, 1.376911e-22, 1.374455e-22, 
    1.376816e-22, 1.367894e-22, 1.371876e-22, 1.36098e-22, 1.363622e-22, 
    1.362408e-22, 1.361073e-22, 1.365196e-22, 1.369589e-22, 1.369693e-22, 
    1.371103e-22, 1.375064e-22, 1.368243e-22, 1.390509e-22, 1.376332e-22, 
    1.356856e-22, 1.36083e-22, 1.36141e-22, 1.359867e-22, 1.370386e-22, 
    1.366565e-22, 1.376876e-22, 1.374085e-22, 1.378662e-22, 1.376385e-22, 
    1.37605e-22, 1.373133e-22, 1.371317e-22, 1.366738e-22, 1.363025e-22, 
    1.360092e-22, 1.360774e-22, 1.363998e-22, 1.369861e-22, 1.375433e-22, 
    1.374209e-22, 1.378314e-22, 1.367487e-22, 1.372014e-22, 1.37026e-22, 
    1.374839e-22, 1.364832e-22, 1.37332e-22, 1.362666e-22, 1.363599e-22, 
    1.366489e-22, 1.372315e-22, 1.373621e-22, 1.374999e-22, 1.37415e-22, 
    1.370012e-22, 1.369339e-22, 1.366421e-22, 1.365612e-22, 1.363397e-22, 
    1.36156e-22, 1.363235e-22, 1.364995e-22, 1.370018e-22, 1.374551e-22, 
    1.379527e-22, 1.380795e-22, 1.387181e-22, 1.381931e-22, 1.390588e-22, 
    1.383205e-22, 1.396016e-22, 1.373828e-22, 1.383008e-22, 1.366624e-22, 
    1.368358e-22, 1.371488e-22, 1.37871e-22, 1.374818e-22, 1.379386e-22, 
    1.369313e-22, 1.364105e-22, 1.362772e-22, 1.360268e-22, 1.362829e-22, 
    1.362621e-22, 1.365075e-22, 1.364286e-22, 1.370185e-22, 1.367014e-22, 
    1.376039e-22, 1.379351e-22, 1.38961e-22, 1.396009e-22, 1.402562e-22, 
    1.405457e-22, 1.40634e-22, 1.406708e-22,
  1.832321e-27, 1.841509e-27, 1.83972e-27, 1.847307e-27, 1.843033e-27, 
    1.84809e-27, 1.834178e-27, 1.84187e-27, 1.836959e-27, 1.833146e-27, 
    1.862512e-27, 1.847657e-27, 1.878116e-27, 1.868547e-27, 1.892685e-27, 
    1.876616e-27, 1.895942e-27, 1.892233e-27, 1.903495e-27, 1.900231e-27, 
    1.915548e-27, 1.905049e-27, 1.923766e-27, 1.913024e-27, 1.914696e-27, 
    1.904714e-27, 1.850651e-27, 1.860653e-27, 1.850057e-27, 1.85148e-27, 
    1.850844e-27, 1.843114e-27, 1.839378e-27, 1.831652e-27, 1.833028e-27, 
    1.838733e-27, 1.852121e-27, 1.847486e-27, 1.859214e-27, 1.858948e-27, 
    1.872074e-27, 1.866145e-27, 1.888342e-27, 1.882012e-27, 1.900365e-27, 
    1.895733e-27, 1.900145e-27, 1.898808e-27, 1.900163e-27, 1.893373e-27, 
    1.896279e-27, 1.890319e-27, 1.867251e-27, 1.874e-27, 1.853931e-27, 
    1.842038e-27, 1.834513e-27, 1.829296e-27, 1.830024e-27, 1.831408e-27, 
    1.838766e-27, 1.845853e-27, 1.851446e-27, 1.855201e-27, 1.85891e-27, 
    1.870142e-27, 1.876142e-27, 1.889617e-27, 1.887191e-27, 1.891312e-27, 
    1.895273e-27, 1.901924e-27, 1.90083e-27, 1.903823e-27, 1.891212e-27, 
    1.89954e-27, 1.885807e-27, 1.889553e-27, 1.859874e-27, 1.848738e-27, 
    1.844012e-27, 1.840062e-27, 1.830582e-27, 1.8371e-27, 1.834499e-27, 
    1.840702e-27, 1.844696e-27, 1.842697e-27, 1.855304e-27, 1.850365e-27, 
    1.876499e-27, 1.865201e-27, 1.894811e-27, 1.88769e-27, 1.896523e-27, 
    1.892013e-27, 1.899742e-27, 1.892785e-27, 1.904968e-27, 1.907761e-27, 
    1.905838e-27, 1.913381e-27, 1.892399e-27, 1.900141e-27, 1.84264e-27, 
    1.842958e-27, 1.844484e-27, 1.837919e-27, 1.837523e-27, 1.831613e-27, 
    1.836871e-27, 1.839126e-27, 1.844938e-27, 1.848487e-27, 1.851889e-27, 
    1.859389e-27, 1.86779e-27, 1.87961e-27, 1.88815e-27, 1.893892e-27, 
    1.890372e-27, 1.893479e-27, 1.890005e-27, 1.88838e-27, 1.906686e-27, 
    1.896303e-27, 1.912288e-27, 1.911359e-27, 1.903894e-27, 1.911464e-27, 
    1.843182e-27, 1.841352e-27, 1.835001e-27, 1.83997e-27, 1.830989e-27, 
    1.83598e-27, 1.838885e-27, 1.850458e-27, 1.853077e-27, 1.855493e-27, 
    1.860286e-27, 1.866448e-27, 1.877299e-27, 1.886794e-27, 1.895506e-27, 
    1.894867e-27, 1.895092e-27, 1.897037e-27, 1.892214e-27, 1.897831e-27, 
    1.89877e-27, 1.896307e-27, 1.911234e-27, 1.906743e-27, 1.911339e-27, 
    1.908411e-27, 1.841948e-27, 1.845094e-27, 1.843363e-27, 1.846617e-27, 
    1.844319e-27, 1.854613e-27, 1.857717e-27, 1.872317e-27, 1.866324e-27, 
    1.875883e-27, 1.867296e-27, 1.868813e-27, 1.876176e-27, 1.867762e-27, 
    1.886261e-27, 1.873684e-27, 1.897113e-27, 1.884472e-27, 1.897907e-27, 
    1.895468e-27, 1.899512e-27, 1.903166e-27, 1.908e-27, 1.917245e-27, 
    1.915103e-27, 1.922864e-27, 1.849908e-27, 1.854114e-27, 1.853751e-27, 
    1.858168e-27, 1.861438e-27, 1.868555e-27, 1.880012e-27, 1.875699e-27, 
    1.883634e-27, 1.885227e-27, 1.873181e-27, 1.88056e-27, 1.85694e-27, 
    1.860729e-27, 1.858478e-27, 1.850234e-27, 1.87668e-27, 1.86306e-27, 
    1.88829e-27, 1.88086e-27, 1.902625e-27, 1.89176e-27, 1.913923e-27, 
    1.923959e-27, 1.933487e-27, 1.944874e-27, 1.856422e-27, 1.853559e-27, 
    1.858696e-27, 1.865809e-27, 1.872456e-27, 1.881311e-27, 1.882224e-27, 
    1.883886e-27, 1.888206e-27, 1.891841e-27, 1.884403e-27, 1.892754e-27, 
    1.861591e-27, 1.877871e-27, 1.85247e-27, 1.860074e-27, 1.865393e-27, 
    1.863067e-27, 1.875209e-27, 1.878078e-27, 1.889775e-27, 1.883726e-27, 
    1.92147e-27, 1.903955e-27, 1.953658e-27, 1.939366e-27, 1.852558e-27, 
    1.856416e-27, 1.869891e-27, 1.86347e-27, 1.881909e-27, 1.886469e-27, 
    1.89019e-27, 1.894942e-27, 1.895463e-27, 1.898285e-27, 1.893661e-27, 
    1.898106e-27, 1.88133e-27, 1.888812e-27, 1.868357e-27, 1.873312e-27, 
    1.871034e-27, 1.868531e-27, 1.876263e-27, 1.884518e-27, 1.884708e-27, 
    1.88736e-27, 1.894824e-27, 1.881984e-27, 1.923731e-27, 1.897209e-27, 
    1.860632e-27, 1.868081e-27, 1.869165e-27, 1.866271e-27, 1.88601e-27, 
    1.878834e-27, 1.898218e-27, 1.892965e-27, 1.901583e-27, 1.897295e-27, 
    1.896664e-27, 1.891175e-27, 1.887761e-27, 1.87916e-27, 1.872193e-27, 
    1.866692e-27, 1.867971e-27, 1.874019e-27, 1.885027e-27, 1.895503e-27, 
    1.893202e-27, 1.900927e-27, 1.880565e-27, 1.889073e-27, 1.885776e-27, 
    1.894385e-27, 1.875582e-27, 1.891541e-27, 1.871517e-27, 1.873268e-27, 
    1.878692e-27, 1.889642e-27, 1.892092e-27, 1.894687e-27, 1.893088e-27, 
    1.88531e-27, 1.884044e-27, 1.878564e-27, 1.877046e-27, 1.872888e-27, 
    1.869444e-27, 1.872586e-27, 1.875889e-27, 1.885319e-27, 1.893845e-27, 
    1.903218e-27, 1.905619e-27, 1.917529e-27, 1.907764e-27, 1.923881e-27, 
    1.910142e-27, 1.933992e-27, 1.89249e-27, 1.909768e-27, 1.878944e-27, 
    1.8822e-27, 1.888087e-27, 1.901678e-27, 1.894345e-27, 1.902954e-27, 
    1.883996e-27, 1.874221e-27, 1.871716e-27, 1.867024e-27, 1.871824e-27, 
    1.871433e-27, 1.876035e-27, 1.874556e-27, 1.885633e-27, 1.879676e-27, 
    1.896644e-27, 1.902886e-27, 1.922044e-27, 1.933973e-27, 1.946497e-27, 
    1.952061e-27, 1.953758e-27, 1.954467e-27,
  8.06339e-33, 8.118358e-33, 8.107643e-33, 8.15271e-33, 8.127482e-33, 
    8.157306e-33, 8.074477e-33, 8.120527e-33, 8.091114e-33, 8.068299e-33, 
    8.242991e-33, 8.154762e-33, 8.337307e-33, 8.279387e-33, 8.425708e-33, 
    8.328233e-33, 8.445504e-33, 8.422942e-33, 8.491361e-33, 8.471579e-33, 
    8.562953e-33, 8.500693e-33, 8.611592e-33, 8.548006e-33, 8.557901e-33, 
    8.498683e-33, 8.172321e-33, 8.231767e-33, 8.168835e-33, 8.177199e-33, 
    8.173458e-33, 8.127972e-33, 8.105616e-33, 8.059411e-33, 8.067596e-33, 
    8.101738e-33, 8.180964e-33, 8.153746e-33, 8.223016e-33, 8.221415e-33, 
    8.300711e-33, 8.264866e-33, 8.399303e-33, 8.360892e-33, 8.472397e-33, 
    8.444212e-33, 8.47106e-33, 8.462919e-33, 8.471167e-33, 8.429871e-33, 
    8.447537e-33, 8.411306e-33, 8.271556e-33, 8.312373e-33, 8.19159e-33, 
    8.121555e-33, 8.076481e-33, 8.045438e-33, 8.049752e-33, 8.057973e-33, 
    8.101937e-33, 8.144133e-33, 8.176983e-33, 8.199041e-33, 8.221184e-33, 
    8.289073e-33, 8.325356e-33, 8.407061e-33, 8.39231e-33, 8.417352e-33, 
    8.441416e-33, 8.481896e-33, 8.475228e-33, 8.493338e-33, 8.416728e-33, 
    8.46739e-33, 8.383907e-33, 8.406656e-33, 8.227072e-33, 8.16109e-33, 
    8.133314e-33, 8.109694e-33, 8.053067e-33, 8.091961e-33, 8.076401e-33, 
    8.113511e-33, 8.137314e-33, 8.125459e-33, 8.199645e-33, 8.17064e-33, 
    8.327512e-33, 8.259175e-33, 8.438606e-33, 8.39534e-33, 8.449016e-33, 
    8.421595e-33, 8.468615e-33, 8.426287e-33, 8.500213e-33, 8.516904e-33, 
    8.505443e-33, 8.550102e-33, 8.423941e-33, 8.471041e-33, 8.125123e-33, 
    8.127027e-33, 8.136065e-33, 8.096867e-33, 8.094495e-33, 8.05918e-33, 
    8.090586e-33, 8.104087e-33, 8.138733e-33, 8.15962e-33, 8.179588e-33, 
    8.22408e-33, 8.274821e-33, 8.346347e-33, 8.398136e-33, 8.433012e-33, 
    8.411624e-33, 8.430502e-33, 8.409393e-33, 8.399526e-33, 8.510539e-33, 
    8.447689e-33, 8.543641e-33, 8.538147e-33, 8.493768e-33, 8.538767e-33, 
    8.128369e-33, 8.117406e-33, 8.079398e-33, 8.109128e-33, 8.055477e-33, 
    8.08526e-33, 8.102655e-33, 8.171201e-33, 8.186561e-33, 8.200765e-33, 
    8.22949e-33, 8.266695e-33, 8.332346e-33, 8.389914e-33, 8.442827e-33, 
    8.438943e-33, 8.440308e-33, 8.452147e-33, 8.422821e-33, 8.456973e-33, 
    8.462698e-33, 8.447706e-33, 8.537411e-33, 8.510866e-33, 8.538031e-33, 
    8.520731e-33, 8.120973e-33, 8.139656e-33, 8.129454e-33, 8.148641e-33, 
    8.1351e-33, 8.195605e-33, 8.214016e-33, 8.302203e-33, 8.26595e-33, 
    8.323775e-33, 8.271822e-33, 8.280993e-33, 8.325582e-33, 8.274635e-33, 
    8.386691e-33, 8.310484e-33, 8.452608e-33, 8.375851e-33, 8.457436e-33, 
    8.442597e-33, 8.4672e-33, 8.489397e-33, 8.518303e-33, 8.572976e-33, 
    8.560295e-33, 8.606239e-33, 8.167956e-33, 8.192664e-33, 8.190524e-33, 
    8.216711e-33, 8.236446e-33, 8.279428e-33, 8.348777e-33, 8.322645e-33, 
    8.370723e-33, 8.380394e-33, 8.307399e-33, 8.352106e-33, 8.209318e-33, 
    8.232185e-33, 8.21859e-33, 8.16988e-33, 8.328607e-33, 8.246254e-33, 
    8.398987e-33, 8.353916e-33, 8.486148e-33, 8.420081e-33, 8.553313e-33, 
    8.612755e-33, 8.669236e-33, 8.73726e-33, 8.206222e-33, 8.189393e-33, 
    8.219894e-33, 8.262855e-33, 8.303019e-33, 8.356651e-33, 8.362178e-33, 
    8.372258e-33, 8.39847e-33, 8.420549e-33, 8.37541e-33, 8.426096e-33, 
    8.237422e-33, 8.335811e-33, 8.183005e-33, 8.228236e-33, 8.260333e-33, 
    8.246277e-33, 8.319673e-33, 8.33705e-33, 8.408016e-33, 8.371281e-33, 
    8.598014e-33, 8.494152e-33, 8.790544e-33, 8.704308e-33, 8.183512e-33, 
    8.206181e-33, 8.287517e-33, 8.24871e-33, 8.360263e-33, 8.387929e-33, 
    8.410517e-33, 8.439412e-33, 8.442566e-33, 8.459743e-33, 8.431609e-33, 
    8.458644e-33, 8.356765e-33, 8.402154e-33, 8.278222e-33, 8.308199e-33, 
    8.294409e-33, 8.279279e-33, 8.326055e-33, 8.37611e-33, 8.377244e-33, 
    8.393347e-33, 8.438771e-33, 8.36072e-33, 8.611452e-33, 8.453265e-33, 
    8.231571e-33, 8.27659e-33, 8.283114e-33, 8.265621e-33, 8.385149e-33, 
    8.341639e-33, 8.459333e-33, 8.427381e-33, 8.479811e-33, 8.453712e-33, 
    8.449877e-33, 8.416501e-33, 8.395769e-33, 8.343617e-33, 8.301434e-33, 
    8.268164e-33, 8.275892e-33, 8.312482e-33, 8.379196e-33, 8.442824e-33, 
    8.428837e-33, 8.475815e-33, 8.352123e-33, 8.403746e-33, 8.383737e-33, 
    8.436015e-33, 8.321938e-33, 8.4188e-33, 8.297332e-33, 8.307926e-33, 
    8.340778e-33, 8.407217e-33, 8.422076e-33, 8.437858e-33, 8.428129e-33, 
    8.380907e-33, 8.373222e-33, 8.339993e-33, 8.330811e-33, 8.305623e-33, 
    8.284797e-33, 8.303807e-33, 8.323805e-33, 8.380953e-33, 8.43274e-33, 
    8.489712e-33, 8.504119e-33, 8.574691e-33, 8.516945e-33, 8.612342e-33, 
    8.531043e-33, 8.672298e-33, 8.424537e-33, 8.528791e-33, 8.342297e-33, 
    8.362029e-33, 8.397769e-33, 8.480425e-33, 8.43577e-33, 8.488138e-33, 
    8.372927e-33, 8.313717e-33, 8.29854e-33, 8.270171e-33, 8.29919e-33, 
    8.296829e-33, 8.324678e-33, 8.315722e-33, 8.382857e-33, 8.346732e-33, 
    8.449763e-33, 8.487727e-33, 8.60139e-33, 8.672146e-33, 8.746944e-33, 
    8.780739e-33, 8.791143e-33, 8.795492e-33,
  1.162231e-38, 1.173476e-38, 1.17128e-38, 1.180474e-38, 1.175345e-38, 
    1.181406e-38, 1.164497e-38, 1.173922e-38, 1.167898e-38, 1.163235e-38, 
    1.198878e-38, 1.18089e-38, 1.21827e-38, 1.206338e-38, 1.236963e-38, 
    1.216399e-38, 1.241184e-38, 1.236369e-38, 1.250969e-38, 1.246751e-38, 
    1.266018e-38, 1.252943e-38, 1.276247e-38, 1.262877e-38, 1.264955e-38, 
    1.252518e-38, 1.184452e-38, 1.19658e-38, 1.183744e-38, 1.185444e-38, 
    1.184683e-38, 1.175447e-38, 1.170869e-38, 1.161406e-38, 1.163092e-38, 
    1.170073e-38, 1.186209e-38, 1.180682e-38, 1.194776e-38, 1.194449e-38, 
    1.210723e-38, 1.203354e-38, 1.231339e-38, 1.223186e-38, 1.246926e-38, 
    1.240904e-38, 1.246641e-38, 1.244899e-38, 1.246664e-38, 1.237846e-38, 
    1.241614e-38, 1.233891e-38, 1.204729e-38, 1.213126e-38, 1.188368e-38, 
    1.174136e-38, 1.164907e-38, 1.158519e-38, 1.15941e-38, 1.16111e-38, 
    1.170114e-38, 1.17873e-38, 1.185397e-38, 1.189882e-38, 1.194402e-38, 
    1.208335e-38, 1.215804e-38, 1.232991e-38, 1.229852e-38, 1.235181e-38, 
    1.240307e-38, 1.248961e-38, 1.247533e-38, 1.251389e-38, 1.235045e-38, 
    1.245858e-38, 1.228066e-38, 1.232902e-38, 1.195619e-38, 1.182171e-38, 
    1.176539e-38, 1.171701e-38, 1.160095e-38, 1.168072e-38, 1.164892e-38, 
    1.172481e-38, 1.177345e-38, 1.174929e-38, 1.190005e-38, 1.18411e-38, 
    1.216249e-38, 1.202188e-38, 1.239708e-38, 1.230496e-38, 1.241929e-38, 
    1.236081e-38, 1.246119e-38, 1.237081e-38, 1.252843e-38, 1.256364e-38, 
    1.25395e-38, 1.263314e-38, 1.236581e-38, 1.246638e-38, 1.174861e-38, 
    1.175251e-38, 1.177091e-38, 1.169076e-38, 1.16859e-38, 1.161359e-38, 
    1.167789e-38, 1.170553e-38, 1.177632e-38, 1.181873e-38, 1.185927e-38, 
    1.194995e-38, 1.205401e-38, 1.220135e-38, 1.23109e-38, 1.238514e-38, 
    1.233958e-38, 1.237979e-38, 1.233484e-38, 1.231384e-38, 1.255031e-38, 
    1.241648e-38, 1.26196e-38, 1.260808e-38, 1.25148e-38, 1.260938e-38, 
    1.175526e-38, 1.173278e-38, 1.165503e-38, 1.171583e-38, 1.160593e-38, 
    1.166701e-38, 1.170261e-38, 1.184226e-38, 1.187344e-38, 1.190234e-38, 
    1.196102e-38, 1.20373e-38, 1.217244e-38, 1.229345e-38, 1.240608e-38, 
    1.239779e-38, 1.24007e-38, 1.242598e-38, 1.236343e-38, 1.243629e-38, 
    1.244854e-38, 1.24165e-38, 1.260654e-38, 1.255097e-38, 1.260784e-38, 
    1.257161e-38, 1.174009e-38, 1.17782e-38, 1.175749e-38, 1.179646e-38, 
    1.176896e-38, 1.189187e-38, 1.192941e-38, 1.211033e-38, 1.203577e-38, 
    1.215476e-38, 1.204782e-38, 1.206668e-38, 1.215855e-38, 1.205359e-38, 
    1.228663e-38, 1.21274e-38, 1.242697e-38, 1.226366e-38, 1.243728e-38, 
    1.240558e-38, 1.245814e-38, 1.250555e-38, 1.256654e-38, 1.268119e-38, 
    1.265454e-38, 1.275117e-38, 1.183565e-38, 1.188587e-38, 1.188149e-38, 
    1.193487e-38, 1.197527e-38, 1.206344e-38, 1.220635e-38, 1.21524e-38, 
    1.22527e-38, 1.227322e-38, 1.212098e-38, 1.221328e-38, 1.191977e-38, 
    1.196658e-38, 1.193872e-38, 1.183957e-38, 1.216474e-38, 1.19954e-38, 
    1.231272e-38, 1.221709e-38, 1.249869e-38, 1.235763e-38, 1.263989e-38, 
    1.276497e-38, 1.288428e-38, 1.302888e-38, 1.191344e-38, 1.187919e-38, 
    1.194138e-38, 1.202945e-38, 1.211198e-38, 1.222289e-38, 1.223459e-38, 
    1.225596e-38, 1.23116e-38, 1.235858e-38, 1.226268e-38, 1.23704e-38, 
    1.197736e-38, 1.217959e-38, 1.186622e-38, 1.19585e-38, 1.202426e-38, 
    1.199541e-38, 1.214627e-38, 1.218212e-38, 1.233194e-38, 1.225388e-38, 
    1.273391e-38, 1.251565e-38, 1.314408e-38, 1.295819e-38, 1.186724e-38, 
    1.191335e-38, 1.20801e-38, 1.20004e-38, 1.223053e-38, 1.228922e-38, 
    1.233722e-38, 1.239881e-38, 1.240552e-38, 1.244222e-38, 1.238215e-38, 
    1.243986e-38, 1.222313e-38, 1.231944e-38, 1.206096e-38, 1.212264e-38, 
    1.209424e-38, 1.206313e-38, 1.215943e-38, 1.226417e-38, 1.226653e-38, 
    1.230074e-38, 1.239759e-38, 1.223149e-38, 1.276231e-38, 1.242851e-38, 
    1.196528e-38, 1.205766e-38, 1.207103e-38, 1.203508e-38, 1.228332e-38, 
    1.21916e-38, 1.244133e-38, 1.237314e-38, 1.248513e-38, 1.242932e-38, 
    1.242113e-38, 1.234996e-38, 1.230587e-38, 1.21957e-38, 1.210872e-38, 
    1.20403e-38, 1.205617e-38, 1.213147e-38, 1.227071e-38, 1.240609e-38, 
    1.237627e-38, 1.247658e-38, 1.221329e-38, 1.232285e-38, 1.228034e-38, 
    1.239155e-38, 1.215095e-38, 1.2355e-38, 1.210025e-38, 1.212207e-38, 
    1.218983e-38, 1.233026e-38, 1.236184e-38, 1.23955e-38, 1.237473e-38, 
    1.227433e-38, 1.225801e-38, 1.218819e-38, 1.216926e-38, 1.211732e-38, 
    1.207447e-38, 1.211359e-38, 1.215481e-38, 1.227441e-38, 1.238458e-38, 
    1.250623e-38, 1.253669e-38, 1.268486e-38, 1.256378e-38, 1.27642e-38, 
    1.259338e-38, 1.289089e-38, 1.236716e-38, 1.258858e-38, 1.219295e-38, 
    1.223427e-38, 1.231016e-38, 1.248651e-38, 1.239103e-38, 1.250293e-38, 
    1.225738e-38, 1.213404e-38, 1.210274e-38, 1.204443e-38, 1.210408e-38, 
    1.209922e-38, 1.215659e-38, 1.213812e-38, 1.227845e-38, 1.220211e-38, 
    1.24209e-38, 1.250205e-38, 1.274097e-38, 1.289049e-38, 1.304969e-38, 
    1.31228e-38, 1.314536e-38, 1.31548e-38,
  5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 7.006492e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 5.605194e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  9.311208e-06, 9.153605e-06, 9.184262e-06, 9.057017e-06, 9.127622e-06, 
    9.044275e-06, 9.279276e-06, 9.147341e-06, 9.231584e-06, 9.297032e-06, 
    8.809661e-06, 9.051337e-06, 8.558091e-06, 8.712626e-06, 8.324022e-06, 
    8.58215e-06, 8.2719e-06, 8.331484e-06, 8.152067e-06, 8.203497e-06, 
    7.973681e-06, 8.128322e-06, 7.854369e-06, 8.010635e-06, 7.986201e-06, 
    8.133419e-06, 9.002747e-06, 8.839776e-06, 9.012395e-06, 8.989172e-06, 
    8.999594e-06, 9.126162e-06, 9.189887e-06, 9.323248e-06, 9.299049e-06, 
    9.201096e-06, 8.978727e-06, 9.054264e-06, 8.863806e-06, 8.868111e-06, 
    8.655701e-06, 8.751522e-06, 8.393909e-06, 8.495666e-06, 8.20135e-06, 
    8.275442e-06, 8.204831e-06, 8.226248e-06, 8.204552e-06, 8.313196e-06, 
    8.26666e-06, 8.362215e-06, 8.733581e-06, 8.624565e-06, 8.949387e-06, 
    9.144242e-06, 9.273492e-06, 9.365116e-06, 9.352168e-06, 9.327478e-06, 
    9.200523e-06, 9.081034e-06, 8.989888e-06, 8.928876e-06, 8.86873e-06, 
    8.68646e-06, 8.589881e-06, 8.373317e-06, 8.412437e-06, 8.346159e-06, 
    8.282811e-06, 8.176366e-06, 8.193894e-06, 8.146971e-06, 8.347913e-06, 
    8.214405e-06, 8.434712e-06, 8.374501e-06, 8.852355e-06, 9.033892e-06, 
    9.11095e-06, 9.178369e-06, 9.34221e-06, 9.229088e-06, 9.273695e-06, 
    9.167548e-06, 9.100047e-06, 9.133439e-06, 8.927208e-06, 9.007429e-06, 
    8.584154e-06, 8.766669e-06, 8.290202e-06, 8.40441e-06, 8.26281e-06, 
    8.335089e-06, 8.211213e-06, 8.322707e-06, 8.129504e-06, 8.087387e-06, 
    8.11617e-06, 8.005571e-06, 8.328883e-06, 8.204829e-06, 9.134373e-06, 
    9.128928e-06, 9.103558e-06, 9.215034e-06, 9.221851e-06, 9.323911e-06, 
    9.233104e-06, 9.194411e-06, 9.096135e-06, 9.037962e-06, 8.982634e-06, 
    8.860892e-06, 8.72477e-06, 8.534153e-06, 8.39701e-06, 8.304978e-06, 
    8.361421e-06, 8.311591e-06, 8.367293e-06, 8.393392e-06, 8.103169e-06, 
    8.266225e-06, 8.021485e-06, 8.035043e-06, 8.145854e-06, 8.033515e-06, 
    9.125105e-06, 9.156436e-06, 9.265145e-06, 9.180079e-06, 9.33502e-06, 
    9.248316e-06, 9.19843e-06, 9.005749e-06, 8.963376e-06, 8.924064e-06, 
    8.846388e-06, 8.746619e-06, 8.571387e-06, 8.4187e-06, 8.279125e-06, 
    8.289358e-06, 8.285755e-06, 8.25455e-06, 8.331827e-06, 8.241859e-06, 
    8.226751e-06, 8.266246e-06, 8.036858e-06, 8.102442e-06, 8.035331e-06, 
    8.078038e-06, 9.146253e-06, 9.093525e-06, 9.12202e-06, 9.068429e-06, 
    9.106186e-06, 8.938196e-06, 8.887781e-06, 8.651581e-06, 8.748583e-06, 
    8.594169e-06, 8.732909e-06, 8.708336e-06, 8.589122e-06, 8.725417e-06, 
    8.42712e-06, 8.629436e-06, 8.253338e-06, 8.45569e-06, 8.240644e-06, 
    8.279729e-06, 8.215012e-06, 8.157016e-06, 8.084015e-06, 7.949182e-06, 
    7.980419e-06, 7.867569e-06, 9.014872e-06, 8.946394e-06, 8.952428e-06, 
    8.880727e-06, 8.82767e-06, 8.712589e-06, 8.527765e-06, 8.597304e-06, 
    8.469612e-06, 8.443959e-06, 8.637943e-06, 8.518877e-06, 8.900544e-06, 
    8.838964e-06, 8.875635e-06, 9.00947e-06, 8.581278e-06, 8.801229e-06, 
    8.394741e-06, 8.514148e-06, 8.165286e-06, 8.33892e-06, 7.997612e-06, 
    7.85137e-06, 7.713575e-06, 7.552298e-06, 8.909007e-06, 8.955556e-06, 
    8.872198e-06, 8.756761e-06, 8.649556e-06, 8.506868e-06, 8.49226e-06, 
    8.465504e-06, 8.396174e-06, 8.337842e-06, 8.457039e-06, 8.323214e-06, 
    8.824672e-06, 8.562168e-06, 8.973147e-06, 8.849545e-06, 8.76357e-06, 
    8.801297e-06, 8.60525e-06, 8.558993e-06, 8.370821e-06, 8.468138e-06, 
    7.887478e-06, 8.144757e-06, 7.429353e-06, 7.629749e-06, 8.971815e-06, 
    8.909169e-06, 8.690864e-06, 8.794786e-06, 8.497338e-06, 8.423998e-06, 
    8.364344e-06, 8.288031e-06, 8.279792e-06, 8.23455e-06, 8.308678e-06, 
    8.23748e-06, 8.506564e-06, 8.386402e-06, 8.715842e-06, 8.635746e-06, 
    8.672601e-06, 8.713012e-06, 8.588246e-06, 8.455163e-06, 8.452324e-06, 
    8.409615e-06, 8.289157e-06, 8.496131e-06, 7.854216e-06, 8.251082e-06, 
    8.840818e-06, 8.719972e-06, 8.702708e-06, 8.749542e-06, 8.431353e-06, 
    8.546748e-06, 8.235654e-06, 8.319822e-06, 8.181882e-06, 8.250448e-06, 
    8.260531e-06, 8.348526e-06, 8.403272e-06, 8.541459e-06, 8.653768e-06, 
    8.742752e-06, 8.722067e-06, 8.6243e-06, 8.447019e-06, 8.279043e-06, 
    8.315861e-06, 8.192372e-06, 8.518932e-06, 8.382118e-06, 8.435016e-06, 
    8.297031e-06, 8.599151e-06, 8.341915e-06, 8.664803e-06, 8.636533e-06, 
    8.549037e-06, 8.372827e-06, 8.333812e-06, 8.292126e-06, 8.317851e-06, 
    8.442516e-06, 8.462928e-06, 8.551167e-06, 8.575514e-06, 8.642689e-06, 
    8.69827e-06, 8.647487e-06, 8.59413e-06, 8.442466e-06, 8.305602e-06, 
    8.156189e-06, 8.119597e-06, 7.944692e-06, 8.087084e-06, 7.852001e-06, 
    8.051885e-06, 7.705649e-06, 8.326998e-06, 8.05777e-06, 8.545057e-06, 
    8.492667e-06, 8.397839e-06, 8.180036e-06, 8.29768e-06, 8.160087e-06, 
    8.463729e-06, 8.620923e-06, 8.661566e-06, 8.737343e-06, 8.659832e-06, 
    8.666138e-06, 8.591924e-06, 8.615778e-06, 8.437427e-06, 8.533265e-06, 
    8.260783e-06, 8.161176e-06, 7.879399e-06, 7.706298e-06, 7.529819e-06, 
    7.451811e-06, 7.428057e-06, 7.418126e-06,
  3.99803e-06, 3.863622e-06, 3.889628e-06, 3.782136e-06, 3.841638e-06, 
    3.771439e-06, 3.970658e-06, 3.858313e-06, 3.929905e-06, 3.985873e-06, 
    3.576616e-06, 3.777368e-06, 3.372439e-06, 3.497294e-06, 3.186959e-06, 
    3.391749e-06, 3.146266e-06, 3.192811e-06, 3.053564e-06, 3.093207e-06, 
    2.917772e-06, 3.035336e-06, 2.828481e-06, 2.945685e-06, 2.927218e-06, 
    3.039244e-06, 3.736663e-06, 3.601387e-06, 3.744731e-06, 3.725316e-06, 
    3.734026e-06, 3.840401e-06, 3.894399e-06, 4.008378e-06, 3.987604e-06, 
    3.903934e-06, 3.716598e-06, 3.779832e-06, 3.621233e-06, 3.624787e-06, 
    3.451087e-06, 3.529014e-06, 3.241882e-06, 3.322552e-06, 3.091548e-06, 
    3.149032e-06, 3.094237e-06, 3.110814e-06, 3.094021e-06, 3.178496e-06, 
    3.142193e-06, 3.21693e-06, 3.514368e-06, 3.425919e-06, 3.692156e-06, 
    3.85568e-06, 3.965704e-06, 4.044418e-06, 4.033258e-06, 4.012009e-06, 
    3.903446e-06, 3.80234e-06, 3.725921e-06, 3.675112e-06, 3.625298e-06, 
    3.476008e-06, 3.397968e-06, 3.225656e-06, 3.25651e-06, 3.204316e-06, 
    3.154774e-06, 3.072264e-06, 3.085787e-06, 3.049644e-06, 3.205697e-06, 
    3.101639e-06, 3.274132e-06, 3.226593e-06, 3.611753e-06, 3.762737e-06, 
    3.827542e-06, 3.884623e-06, 4.024683e-06, 3.927773e-06, 3.965878e-06, 
    3.875447e-06, 3.81836e-06, 3.846559e-06, 3.673726e-06, 3.740579e-06, 
    3.393364e-06, 3.541393e-06, 3.160537e-06, 3.250169e-06, 3.1392e-06, 
    3.19564e-06, 3.09917e-06, 3.18594e-06, 3.03624e-06, 3.004017e-06, 
    3.026021e-06, 2.941859e-06, 3.190777e-06, 3.094233e-06, 3.847348e-06, 
    3.842743e-06, 3.821322e-06, 3.915797e-06, 3.921605e-06, 4.008946e-06, 
    3.931201e-06, 3.898252e-06, 3.815064e-06, 3.766149e-06, 3.719863e-06, 
    3.618824e-06, 3.507181e-06, 3.353272e-06, 3.244329e-06, 3.172075e-06, 
    3.216309e-06, 3.177244e-06, 3.220924e-06, 3.241478e-06, 3.016072e-06, 
    3.141853e-06, 2.953906e-06, 2.964186e-06, 3.048786e-06, 2.963027e-06, 
    3.839512e-06, 3.866027e-06, 3.958566e-06, 3.88608e-06, 4.018499e-06, 
    3.944181e-06, 3.901665e-06, 3.739167e-06, 3.703807e-06, 3.671113e-06, 
    3.606862e-06, 3.52501e-06, 3.383112e-06, 3.261456e-06, 3.151903e-06, 
    3.159881e-06, 3.157071e-06, 3.132777e-06, 3.193083e-06, 3.12292e-06, 
    3.1112e-06, 3.141873e-06, 2.965564e-06, 3.015521e-06, 2.964405e-06, 
    2.99689e-06, 3.857402e-06, 3.812861e-06, 3.836906e-06, 3.791733e-06, 
    3.823534e-06, 3.682845e-06, 3.641035e-06, 3.447746e-06, 3.526612e-06, 
    3.401422e-06, 3.513822e-06, 3.493803e-06, 3.397349e-06, 3.507716e-06, 
    3.268111e-06, 3.429842e-06, 3.131834e-06, 3.290745e-06, 3.121977e-06, 
    3.152373e-06, 3.102114e-06, 3.057366e-06, 3.001447e-06, 2.899344e-06, 
    2.922862e-06, 2.838304e-06, 3.746807e-06, 3.689666e-06, 3.694692e-06, 
    3.635211e-06, 3.591446e-06, 3.497268e-06, 3.348168e-06, 3.403951e-06, 
    3.301819e-06, 3.281456e-06, 3.436729e-06, 3.341063e-06, 3.651608e-06, 
    3.600736e-06, 3.631e-06, 3.742283e-06, 3.391054e-06, 3.56971e-06, 
    3.242539e-06, 3.337291e-06, 3.06373e-06, 3.198635e-06, 2.935839e-06, 
    2.826245e-06, 2.724702e-06, 2.607962e-06, 3.658623e-06, 3.697296e-06, 
    3.628163e-06, 3.533287e-06, 3.446115e-06, 3.33148e-06, 3.319839e-06, 
    3.298553e-06, 3.243672e-06, 3.197797e-06, 3.291826e-06, 3.186338e-06, 
    3.588958e-06, 3.375714e-06, 3.711948e-06, 3.609454e-06, 3.538858e-06, 
    3.569772e-06, 3.410351e-06, 3.373173e-06, 3.223694e-06, 3.300647e-06, 
    2.85313e-06, 3.047937e-06, 2.520551e-06, 2.663734e-06, 3.710841e-06, 
    3.65876e-06, 3.479597e-06, 3.564432e-06, 3.323884e-06, 3.265649e-06, 
    3.218606e-06, 3.158842e-06, 3.152422e-06, 3.117248e-06, 3.174966e-06, 
    3.119523e-06, 3.331237e-06, 3.235966e-06, 3.499918e-06, 3.43495e-06, 
    3.464784e-06, 3.497613e-06, 3.396665e-06, 3.290335e-06, 3.288091e-06, 
    3.254277e-06, 3.159692e-06, 3.322923e-06, 2.828345e-06, 3.130056e-06, 
    3.602274e-06, 3.503269e-06, 3.489228e-06, 3.527399e-06, 3.271469e-06, 
    3.363358e-06, 3.118105e-06, 3.183683e-06, 3.076519e-06, 3.129589e-06, 
    3.137427e-06, 3.206179e-06, 3.249271e-06, 3.359121e-06, 3.449523e-06, 
    3.521855e-06, 3.504987e-06, 3.425706e-06, 3.283876e-06, 3.151835e-06, 
    3.180578e-06, 3.084613e-06, 3.341112e-06, 3.232587e-06, 3.274365e-06, 
    3.165867e-06, 3.405436e-06, 3.200965e-06, 3.458463e-06, 3.435588e-06, 
    3.365192e-06, 3.225267e-06, 3.194638e-06, 3.162036e-06, 3.182141e-06, 
    3.280308e-06, 3.296506e-06, 3.366899e-06, 3.386428e-06, 3.440565e-06, 
    3.485622e-06, 3.444443e-06, 3.401392e-06, 3.280272e-06, 3.172558e-06, 
    3.05673e-06, 3.028648e-06, 2.895957e-06, 3.003776e-06, 2.826696e-06, 
    2.976945e-06, 2.718891e-06, 3.189285e-06, 2.981436e-06, 3.362006e-06, 
    3.320163e-06, 3.244977e-06, 3.075085e-06, 3.166374e-06, 3.059722e-06, 
    3.297142e-06, 3.422976e-06, 3.45584e-06, 3.517439e-06, 3.454436e-06, 
    3.459545e-06, 3.399623e-06, 3.418837e-06, 3.276279e-06, 3.352569e-06, 
    3.13762e-06, 3.060562e-06, 2.847114e-06, 2.719378e-06, 2.591886e-06, 
    2.53642e-06, 2.519641e-06, 2.51264e-06,
  1.84168e-06, 1.771747e-06, 1.78525e-06, 1.729531e-06, 1.760345e-06, 
    1.723999e-06, 1.827408e-06, 1.768993e-06, 1.806189e-06, 1.83534e-06, 
    1.623671e-06, 1.727065e-06, 1.519409e-06, 1.583058e-06, 1.425502e-06, 
    1.52923e-06, 1.405004e-06, 1.428454e-06, 1.358455e-06, 1.378337e-06, 
    1.290643e-06, 1.349327e-06, 1.2463e-06, 1.304545e-06, 1.295345e-06, 
    1.351283e-06, 1.706032e-06, 1.636383e-06, 1.710198e-06, 1.700175e-06, 
    1.704671e-06, 1.759703e-06, 1.787728e-06, 1.847079e-06, 1.836242e-06, 
    1.792683e-06, 1.695677e-06, 1.728339e-06, 1.646577e-06, 1.648404e-06, 
    1.559462e-06, 1.599283e-06, 1.453229e-06, 1.494076e-06, 1.377504e-06, 
    1.406397e-06, 1.378854e-06, 1.387179e-06, 1.378745e-06, 1.421236e-06, 
    1.402955e-06, 1.440624e-06, 1.591788e-06, 1.54663e-06, 1.683074e-06, 
    1.767626e-06, 1.824827e-06, 1.8659e-06, 1.860069e-06, 1.848974e-06, 
    1.79243e-06, 1.739986e-06, 1.700487e-06, 1.674294e-06, 1.648667e-06, 
    1.572181e-06, 1.532395e-06, 1.44503e-06, 1.460625e-06, 1.434257e-06, 
    1.409287e-06, 1.367829e-06, 1.374613e-06, 1.356492e-06, 1.434954e-06, 
    1.38257e-06, 1.469541e-06, 1.445504e-06, 1.641706e-06, 1.719501e-06, 
    1.753038e-06, 1.78265e-06, 1.855591e-06, 1.80508e-06, 1.824917e-06, 
    1.777885e-06, 1.748281e-06, 1.762896e-06, 1.67358e-06, 1.708054e-06, 
    1.530052e-06, 1.60562e-06, 1.412189e-06, 1.457418e-06, 1.401449e-06, 
    1.42988e-06, 1.381331e-06, 1.424989e-06, 1.349779e-06, 1.33366e-06, 
    1.344665e-06, 1.302639e-06, 1.427427e-06, 1.378852e-06, 1.763305e-06, 
    1.760918e-06, 1.749816e-06, 1.79885e-06, 1.801871e-06, 1.847376e-06, 
    1.806863e-06, 1.78973e-06, 1.746574e-06, 1.721265e-06, 1.697362e-06, 
    1.64534e-06, 1.588112e-06, 1.509669e-06, 1.454466e-06, 1.418001e-06, 
    1.44031e-06, 1.420605e-06, 1.442641e-06, 1.453025e-06, 1.339687e-06, 
    1.402784e-06, 1.308644e-06, 1.313771e-06, 1.356061e-06, 1.313192e-06, 
    1.759242e-06, 1.772996e-06, 1.821109e-06, 1.783407e-06, 1.852362e-06, 
    1.813618e-06, 1.791504e-06, 1.707325e-06, 1.68908e-06, 1.672234e-06, 
    1.639195e-06, 1.597233e-06, 1.524836e-06, 1.463126e-06, 1.407842e-06, 
    1.411859e-06, 1.410444e-06, 1.398219e-06, 1.42859e-06, 1.393262e-06, 
    1.387373e-06, 1.402794e-06, 1.314458e-06, 1.339412e-06, 1.31388e-06, 
    1.330099e-06, 1.768521e-06, 1.745433e-06, 1.757891e-06, 1.734496e-06, 
    1.750962e-06, 1.678276e-06, 1.656756e-06, 1.557757e-06, 1.598053e-06, 
    1.534153e-06, 1.591509e-06, 1.581273e-06, 1.532079e-06, 1.588386e-06, 
    1.466493e-06, 1.548628e-06, 1.397744e-06, 1.477952e-06, 1.392788e-06, 
    1.408079e-06, 1.382809e-06, 1.360361e-06, 1.332376e-06, 1.281475e-06, 
    1.293177e-06, 1.251168e-06, 1.71127e-06, 1.681791e-06, 1.684382e-06, 
    1.653762e-06, 1.631281e-06, 1.583045e-06, 1.507077e-06, 1.535441e-06, 
    1.483564e-06, 1.473249e-06, 1.55214e-06, 1.503469e-06, 1.662195e-06, 
    1.636049e-06, 1.651597e-06, 1.708934e-06, 1.528877e-06, 1.620131e-06, 
    1.453561e-06, 1.501554e-06, 1.36355e-06, 1.431391e-06, 1.299639e-06, 
    1.245192e-06, 1.195017e-06, 1.137662e-06, 1.665805e-06, 1.685724e-06, 
    1.650139e-06, 1.60147e-06, 1.556926e-06, 1.498605e-06, 1.492699e-06, 
    1.481908e-06, 1.454134e-06, 1.430968e-06, 1.4785e-06, 1.42519e-06, 
    1.630003e-06, 1.521074e-06, 1.693278e-06, 1.640526e-06, 1.604322e-06, 
    1.620163e-06, 1.5387e-06, 1.519783e-06, 1.444039e-06, 1.48297e-06, 
    1.25852e-06, 1.355636e-06, 1.094955e-06, 1.165018e-06, 1.692707e-06, 
    1.665876e-06, 1.574015e-06, 1.617425e-06, 1.494751e-06, 1.465248e-06, 
    1.44147e-06, 1.411335e-06, 1.408103e-06, 1.390411e-06, 1.419458e-06, 
    1.391555e-06, 1.498482e-06, 1.450239e-06, 1.584399e-06, 1.551233e-06, 
    1.566452e-06, 1.583221e-06, 1.531732e-06, 1.477745e-06, 1.476608e-06, 
    1.459495e-06, 1.411762e-06, 1.494264e-06, 1.246231e-06, 1.396849e-06, 
    1.636839e-06, 1.586112e-06, 1.578935e-06, 1.598456e-06, 1.468193e-06, 
    1.514794e-06, 1.390842e-06, 1.423851e-06, 1.369963e-06, 1.396616e-06, 
    1.400557e-06, 1.435197e-06, 1.456964e-06, 1.51264e-06, 1.558664e-06, 
    1.595619e-06, 1.586991e-06, 1.546521e-06, 1.474474e-06, 1.407807e-06, 
    1.422285e-06, 1.374023e-06, 1.503494e-06, 1.448532e-06, 1.469659e-06, 
    1.414873e-06, 1.536197e-06, 1.432565e-06, 1.563226e-06, 1.551559e-06, 
    1.515726e-06, 1.444834e-06, 1.429375e-06, 1.412944e-06, 1.423074e-06, 
    1.472667e-06, 1.480871e-06, 1.516594e-06, 1.526523e-06, 1.554096e-06, 
    1.577093e-06, 1.556073e-06, 1.534138e-06, 1.472649e-06, 1.418244e-06, 
    1.360041e-06, 1.345979e-06, 1.27979e-06, 1.333539e-06, 1.245415e-06, 
    1.320136e-06, 1.192153e-06, 1.426674e-06, 1.322379e-06, 1.514107e-06, 
    1.492864e-06, 1.454793e-06, 1.369243e-06, 1.415129e-06, 1.361541e-06, 
    1.481193e-06, 1.54513e-06, 1.561887e-06, 1.59336e-06, 1.561171e-06, 
    1.563778e-06, 1.533238e-06, 1.543022e-06, 1.470628e-06, 1.509312e-06, 
    1.400655e-06, 1.361962e-06, 1.255537e-06, 1.192393e-06, 1.129793e-06, 
    1.102693e-06, 1.094512e-06, 1.0911e-06,
  4.641148e-07, 4.427102e-07, 4.468269e-07, 4.298902e-07, 4.3924e-07, 
    4.28216e-07, 4.597298e-07, 4.418715e-07, 4.53226e-07, 4.621657e-07, 
    3.980869e-07, 4.291436e-07, 3.672588e-07, 3.860189e-07, 3.399304e-07, 
    3.701411e-07, 3.340223e-07, 3.407827e-07, 3.206826e-07, 3.263668e-07, 
    3.014446e-07, 3.180792e-07, 2.889934e-07, 3.053696e-07, 3.027712e-07, 
    3.186368e-07, 4.227876e-07, 4.018794e-07, 4.240451e-07, 4.210212e-07, 
    4.22377e-07, 4.390449e-07, 4.475831e-07, 4.65776e-07, 4.62443e-07, 
    4.490964e-07, 4.196655e-07, 4.295295e-07, 4.049263e-07, 4.054727e-07, 
    3.790424e-07, 3.908311e-07, 3.479547e-07, 3.598446e-07, 3.261284e-07, 
    3.344229e-07, 3.26515e-07, 3.289012e-07, 3.264839e-07, 3.386991e-07, 
    3.334328e-07, 3.443021e-07, 3.886068e-07, 3.75259e-07, 4.158722e-07, 
    4.414553e-07, 4.589377e-07, 4.715761e-07, 4.697775e-07, 4.663592e-07, 
    4.490189e-07, 4.330579e-07, 4.211153e-07, 4.132333e-07, 4.055513e-07, 
    3.827999e-07, 3.71071e-07, 3.45578e-07, 3.501015e-07, 3.424599e-07, 
    3.35255e-07, 3.233601e-07, 3.253006e-07, 3.201222e-07, 3.426615e-07, 
    3.275797e-07, 3.526933e-07, 3.457153e-07, 4.034698e-07, 4.268558e-07, 
    4.370191e-07, 4.460336e-07, 4.683972e-07, 4.528865e-07, 4.589654e-07, 
    4.445806e-07, 4.355747e-07, 4.40016e-07, 4.13019e-07, 4.233979e-07, 
    3.703825e-07, 3.927139e-07, 3.360907e-07, 3.491704e-07, 3.329997e-07, 
    3.411949e-07, 3.272245e-07, 3.397822e-07, 3.182081e-07, 3.136212e-07, 
    3.167513e-07, 3.048308e-07, 3.404863e-07, 3.265144e-07, 4.401405e-07, 
    4.394142e-07, 4.360405e-07, 4.509811e-07, 4.519048e-07, 4.658672e-07, 
    4.534324e-07, 4.481945e-07, 4.350564e-07, 4.27389e-07, 4.201731e-07, 
    4.045561e-07, 3.875167e-07, 3.644047e-07, 3.483136e-07, 3.377659e-07, 
    3.442113e-07, 3.385171e-07, 3.44886e-07, 3.478956e-07, 3.153348e-07, 
    3.333835e-07, 3.065284e-07, 3.079795e-07, 3.199995e-07, 3.078158e-07, 
    4.389047e-07, 4.430906e-07, 4.577969e-07, 4.462646e-07, 4.674024e-07, 
    4.55501e-07, 4.487361e-07, 4.231777e-07, 4.176791e-07, 4.12615e-07, 
    4.027196e-07, 3.902225e-07, 3.688511e-07, 3.508283e-07, 3.348389e-07, 
    3.359956e-07, 3.35588e-07, 3.32071e-07, 3.408223e-07, 3.306472e-07, 
    3.289568e-07, 3.333865e-07, 3.081742e-07, 3.152566e-07, 3.080104e-07, 
    3.126096e-07, 4.417277e-07, 4.347103e-07, 4.384941e-07, 4.313939e-07, 
    4.363885e-07, 4.144298e-07, 4.07973e-07, 3.785392e-07, 3.904659e-07, 
    3.715878e-07, 3.88524e-07, 3.854905e-07, 3.709783e-07, 3.875979e-07, 
    3.518069e-07, 3.758477e-07, 3.319347e-07, 3.551417e-07, 3.305111e-07, 
    3.349071e-07, 3.276482e-07, 3.212265e-07, 3.132563e-07, 2.988619e-07, 
    3.021593e-07, 2.903554e-07, 4.243689e-07, 4.154862e-07, 4.162653e-07, 
    4.070764e-07, 4.003564e-07, 3.86015e-07, 3.636458e-07, 3.719665e-07, 
    3.567771e-07, 3.537722e-07, 3.768825e-07, 3.625902e-07, 4.096029e-07, 
    4.017798e-07, 4.064282e-07, 4.236634e-07, 3.700374e-07, 3.970319e-07, 
    3.48051e-07, 3.620302e-07, 3.221373e-07, 3.416314e-07, 3.039834e-07, 
    2.886835e-07, 2.747229e-07, 2.589321e-07, 4.106855e-07, 4.166691e-07, 
    4.059919e-07, 3.914806e-07, 3.782939e-07, 3.61168e-07, 3.594427e-07, 
    3.562945e-07, 3.482172e-07, 3.415094e-07, 3.553013e-07, 3.398401e-07, 
    3.999752e-07, 3.677471e-07, 4.18943e-07, 4.031171e-07, 3.923281e-07, 
    3.970414e-07, 3.729248e-07, 3.673684e-07, 3.45291e-07, 3.566039e-07, 
    2.924145e-07, 3.198781e-07, 2.472932e-07, 2.66441e-07, 4.187711e-07, 
    4.107067e-07, 3.833422e-07, 3.96226e-07, 3.60042e-07, 3.514449e-07, 
    3.445471e-07, 3.358448e-07, 3.349141e-07, 3.298288e-07, 3.38186e-07, 
    3.30157e-07, 3.611321e-07, 3.470876e-07, 3.864163e-07, 3.766152e-07, 
    3.811063e-07, 3.860673e-07, 3.708763e-07, 3.550813e-07, 3.547503e-07, 
    3.497735e-07, 3.359677e-07, 3.598996e-07, 2.889741e-07, 3.316773e-07, 
    4.020158e-07, 3.869238e-07, 3.847982e-07, 3.905856e-07, 3.523012e-07, 
    3.659057e-07, 3.299524e-07, 3.394536e-07, 3.239703e-07, 3.316104e-07, 
    3.327432e-07, 3.427319e-07, 3.490386e-07, 3.652749e-07, 3.788069e-07, 
    3.897434e-07, 3.871844e-07, 3.75227e-07, 3.541288e-07, 3.348289e-07, 
    3.390018e-07, 3.25132e-07, 3.625976e-07, 3.465926e-07, 3.527275e-07, 
    3.368642e-07, 3.721886e-07, 3.419708e-07, 3.801535e-07, 3.767112e-07, 
    3.661789e-07, 3.45521e-07, 3.410489e-07, 3.363082e-07, 3.392293e-07, 
    3.536029e-07, 3.559922e-07, 3.664333e-07, 3.693463e-07, 3.774592e-07, 
    3.84253e-07, 3.780425e-07, 3.715834e-07, 3.535976e-07, 3.37836e-07, 
    3.211353e-07, 3.171257e-07, 2.983878e-07, 3.135868e-07, 2.887457e-07, 
    3.097827e-07, 2.7393e-07, 3.402688e-07, 3.104188e-07, 3.657045e-07, 
    3.594908e-07, 3.484084e-07, 3.237644e-07, 3.369378e-07, 3.215635e-07, 
    3.560861e-07, 3.748173e-07, 3.797581e-07, 3.890729e-07, 3.795467e-07, 
    3.803164e-07, 3.713188e-07, 3.741966e-07, 3.530094e-07, 3.643002e-07, 
    3.327712e-07, 3.216837e-07, 2.915785e-07, 2.739965e-07, 2.567798e-07, 
    2.493944e-07, 2.471729e-07, 2.462477e-07,
  4.229465e-08, 3.984172e-08, 4.031087e-08, 3.83888e-08, 3.944722e-08, 
    3.819997e-08, 4.178942e-08, 3.974629e-08, 4.104261e-08, 4.206991e-08, 
    3.483861e-08, 3.830457e-08, 3.147369e-08, 3.351221e-08, 2.855669e-08, 
    3.1785e-08, 2.793452e-08, 2.86467e-08, 2.654108e-08, 2.713291e-08, 
    2.455988e-08, 2.627099e-08, 2.329599e-08, 2.496132e-08, 2.469539e-08, 
    2.632879e-08, 3.758919e-08, 3.525784e-08, 3.773047e-08, 3.739091e-08, 
    3.754307e-08, 3.942507e-08, 4.039719e-08, 4.248642e-08, 4.210186e-08, 
    4.057005e-08, 3.723891e-08, 3.834809e-08, 3.559545e-08, 3.565608e-08, 
    3.275076e-08, 3.403972e-08, 2.940658e-08, 3.067606e-08, 2.710803e-08, 
    2.797662e-08, 2.714837e-08, 2.739771e-08, 2.714513e-08, 2.842678e-08, 
    2.787261e-08, 2.901903e-08, 3.379567e-08, 3.233948e-08, 3.681434e-08, 
    3.969896e-08, 4.16983e-08, 4.315753e-08, 4.294916e-08, 4.25538e-08, 
    4.056119e-08, 3.874666e-08, 3.740147e-08, 3.651964e-08, 3.56648e-08, 
    3.316038e-08, 3.188559e-08, 2.915427e-08, 2.963491e-08, 2.882401e-08, 
    2.806408e-08, 2.68195e-08, 2.702168e-08, 2.64829e-08, 2.884534e-08, 
    2.725957e-08, 2.991107e-08, 2.916883e-08, 3.543397e-08, 3.804671e-08, 
    3.919522e-08, 4.022036e-08, 4.278941e-08, 4.100372e-08, 4.170148e-08, 
    4.005472e-08, 3.903151e-08, 3.953536e-08, 3.649573e-08, 3.765773e-08, 
    3.181111e-08, 3.424663e-08, 2.815199e-08, 2.953583e-08, 2.782714e-08, 
    2.869025e-08, 2.722246e-08, 2.854105e-08, 2.628436e-08, 2.580993e-08, 
    2.613347e-08, 2.490612e-08, 2.86154e-08, 2.714831e-08, 3.95495e-08, 
    3.9467e-08, 3.908429e-08, 4.078557e-08, 4.089129e-08, 4.249695e-08, 
    4.106627e-08, 4.0467e-08, 3.897282e-08, 3.810677e-08, 3.729581e-08, 
    3.55544e-08, 3.36762e-08, 3.116609e-08, 2.944472e-08, 2.83284e-08, 
    2.900941e-08, 2.840758e-08, 2.90809e-08, 2.94003e-08, 2.598694e-08, 
    2.786744e-08, 2.508012e-08, 2.522905e-08, 2.647015e-08, 2.521224e-08, 
    3.940915e-08, 3.988501e-08, 4.156715e-08, 4.024672e-08, 4.267436e-08, 
    4.130349e-08, 4.052887e-08, 3.763301e-08, 3.701644e-08, 3.645066e-08, 
    3.535085e-08, 3.397291e-08, 3.164559e-08, 2.971229e-08, 2.802033e-08, 
    2.814198e-08, 2.809911e-08, 2.77297e-08, 2.865088e-08, 2.758047e-08, 
    2.740353e-08, 2.786775e-08, 2.524904e-08, 2.597885e-08, 2.523222e-08, 
    2.570556e-08, 3.972993e-08, 3.893362e-08, 3.936254e-08, 3.855858e-08, 
    3.912373e-08, 3.665319e-08, 3.593379e-08, 3.2696e-08, 3.399963e-08, 
    3.194153e-08, 3.378658e-08, 3.34544e-08, 3.187556e-08, 3.36851e-08, 
    2.981656e-08, 3.240341e-08, 2.771541e-08, 3.017249e-08, 2.756622e-08, 
    2.80275e-08, 2.726672e-08, 2.659758e-08, 2.577227e-08, 2.429651e-08, 
    2.463287e-08, 2.343352e-08, 3.776687e-08, 3.67712e-08, 3.685829e-08, 
    3.583414e-08, 3.508934e-08, 3.351179e-08, 3.108442e-08, 3.198252e-08, 
    3.034739e-08, 3.00262e-08, 3.251583e-08, 3.097089e-08, 3.611508e-08, 
    3.524681e-08, 3.576215e-08, 3.768757e-08, 3.17738e-08, 3.472219e-08, 
    2.941681e-08, 3.091071e-08, 2.669227e-08, 2.873639e-08, 2.481938e-08, 
    2.326473e-08, 2.186577e-08, 2.030673e-08, 3.623562e-08, 3.690344e-08, 
    3.57137e-08, 3.411106e-08, 3.266931e-08, 3.081809e-08, 3.063295e-08, 
    3.029576e-08, 2.943448e-08, 2.872349e-08, 3.018955e-08, 2.854716e-08, 
    3.50472e-08, 3.152638e-08, 3.715795e-08, 3.539489e-08, 3.420421e-08, 
    3.472324e-08, 3.208633e-08, 3.148551e-08, 2.912384e-08, 3.032886e-08, 
    2.364179e-08, 2.645755e-08, 1.917395e-08, 2.104496e-08, 3.71387e-08, 
    3.623797e-08, 3.32196e-08, 3.463332e-08, 3.069723e-08, 2.977798e-08, 
    2.904499e-08, 2.812612e-08, 2.802824e-08, 2.749477e-08, 2.837268e-08, 
    2.752913e-08, 3.081423e-08, 2.931448e-08, 3.35557e-08, 3.248678e-08, 
    3.297562e-08, 3.351751e-08, 3.186452e-08, 3.016604e-08, 3.013067e-08, 
    2.959999e-08, 2.813905e-08, 3.068195e-08, 2.329404e-08, 2.768843e-08, 
    3.527293e-08, 3.361126e-08, 3.337869e-08, 3.401277e-08, 2.986926e-08, 
    3.132778e-08, 2.750771e-08, 2.850637e-08, 2.688304e-08, 2.768141e-08, 
    2.780023e-08, 2.885279e-08, 2.952181e-08, 3.125981e-08, 3.272513e-08, 
    3.392033e-08, 3.36398e-08, 3.233601e-08, 3.006428e-08, 2.801929e-08, 
    2.84587e-08, 2.700409e-08, 3.097168e-08, 2.926193e-08, 2.991472e-08, 
    2.823342e-08, 3.200657e-08, 2.877228e-08, 3.287177e-08, 3.249721e-08, 
    3.135722e-08, 2.914824e-08, 2.867483e-08, 2.817489e-08, 2.84827e-08, 
    3.000813e-08, 3.026342e-08, 3.138465e-08, 3.169909e-08, 3.257852e-08, 
    3.33191e-08, 3.264195e-08, 3.194105e-08, 3.000757e-08, 2.833579e-08, 
    2.658811e-08, 2.617223e-08, 2.424824e-08, 2.580638e-08, 2.3271e-08, 
    2.541439e-08, 2.178689e-08, 2.859242e-08, 2.547984e-08, 3.130609e-08, 
    3.06381e-08, 2.94548e-08, 2.686159e-08, 2.824117e-08, 2.663261e-08, 
    3.027347e-08, 3.229155e-08, 3.28287e-08, 3.384678e-08, 3.280567e-08, 
    3.288952e-08, 3.191241e-08, 3.22242e-08, 2.99448e-08, 3.115484e-08, 
    2.780317e-08, 2.66451e-08, 2.355718e-08, 2.17935e-08, 2.009619e-08, 
    1.937741e-08, 1.916231e-08, 1.907289e-08,
  1.221174e-09, 1.13161e-09, 1.148624e-09, 1.079274e-09, 1.117346e-09, 
    1.072512e-09, 1.202605e-09, 1.128156e-09, 1.175272e-09, 1.212906e-09, 
    9.537289e-10, 1.076256e-09, 8.379684e-10, 9.077097e-10, 7.403452e-10, 
    8.485402e-10, 7.198684e-10, 7.433179e-10, 6.744663e-10, 6.936713e-10, 
    6.110435e-10, 6.657409e-10, 5.713071e-10, 6.237843e-10, 6.153381e-10, 
    6.67606e-10, 1.050703e-09, 9.683763e-10, 1.055739e-09, 1.043645e-09, 
    1.049061e-09, 1.116546e-09, 1.151761e-09, 1.228238e-09, 1.214081e-09, 
    1.158047e-09, 1.038241e-09, 1.077815e-09, 9.80207e-10, 9.823349e-10, 
    8.815176e-10, 9.259521e-10, 7.685161e-10, 8.110145e-10, 6.928615e-10, 
    7.212499e-10, 6.941745e-10, 7.023019e-10, 6.940691e-10, 7.360593e-10, 
    7.178377e-10, 7.556418e-10, 9.175025e-10, 8.674405e-10, 1.023179e-09, 
    1.126444e-09, 1.199262e-09, 1.253031e-09, 1.245322e-09, 1.230723e-09, 
    1.157725e-09, 1.092114e-09, 1.044021e-09, 1.012752e-09, 9.826411e-10, 
    8.955871e-10, 8.519623e-10, 7.601292e-10, 7.76123e-10, 7.491812e-10, 
    7.241222e-10, 6.834864e-10, 6.900529e-10, 6.725845e-10, 7.498871e-10, 
    6.977965e-10, 7.853455e-10, 7.606126e-10, 9.745447e-10, 1.06703e-09, 
    1.108255e-09, 1.145337e-09, 1.239418e-09, 1.173852e-09, 1.199379e-09, 
    1.139328e-09, 1.102358e-09, 1.120529e-09, 1.011908e-09, 1.053146e-09, 
    8.494282e-10, 9.331288e-10, 7.270116e-10, 7.728201e-10, 7.163471e-10, 
    7.447571e-10, 6.965875e-10, 7.398288e-10, 6.66172e-10, 6.509029e-10, 
    6.613076e-10, 6.220293e-10, 7.422837e-10, 6.941725e-10, 1.12104e-09, 
    1.11806e-09, 1.104259e-09, 1.165896e-09, 1.16975e-09, 1.228627e-09, 
    1.176135e-09, 1.154299e-09, 1.100246e-09, 1.069178e-09, 1.040263e-09, 
    9.787668e-10, 9.133725e-10, 8.275512e-10, 7.697856e-10, 7.328171e-10, 
    7.553227e-10, 7.354264e-10, 7.57694e-10, 7.683069e-10, 6.565911e-10, 
    7.176681e-10, 6.275658e-10, 6.323131e-10, 6.721724e-10, 6.317769e-10, 
    1.115972e-09, 1.133177e-09, 1.194455e-09, 1.146294e-09, 1.23517e-09, 
    1.184804e-09, 1.156549e-09, 1.052265e-09, 1.030343e-09, 1.010315e-09, 
    9.716324e-10, 9.236374e-10, 8.438024e-10, 7.787049e-10, 7.226852e-10, 
    7.266825e-10, 7.252732e-10, 7.131548e-10, 7.434559e-10, 7.082719e-10, 
    7.024917e-10, 7.176782e-10, 6.32951e-10, 6.563309e-10, 6.324143e-10, 
    6.475542e-10, 1.127564e-09, 1.098835e-09, 1.114289e-09, 1.085361e-09, 
    1.105679e-09, 1.017475e-09, 9.92095e-10, 8.796405e-10, 9.24563e-10, 
    8.538664e-10, 9.171883e-10, 9.057153e-10, 8.516208e-10, 9.136799e-10, 
    7.821866e-10, 8.696251e-10, 7.12687e-10, 7.940973e-10, 7.07806e-10, 
    7.229206e-10, 6.980296e-10, 6.762948e-10, 6.496944e-10, 6.027158e-10, 
    6.133558e-10, 5.756029e-10, 1.057038e-09, 1.021651e-09, 1.024736e-09, 
    9.885903e-10, 9.624831e-10, 9.076951e-10, 8.247901e-10, 8.552623e-10, 
    7.999642e-10, 7.891972e-10, 8.734703e-10, 8.209554e-10, 9.984776e-10, 
    9.679901e-10, 9.860601e-10, 1.05421e-09, 8.481592e-10, 9.496698e-10, 
    7.688565e-10, 8.18924e-10, 6.793612e-10, 7.462824e-10, 6.192731e-10, 
    5.703316e-10, 5.270528e-10, 4.797119e-10, 1.002726e-09, 1.026336e-09, 
    9.843584e-10, 9.284254e-10, 8.787257e-10, 8.158002e-10, 8.095633e-10, 
    7.982313e-10, 7.694447e-10, 7.45856e-10, 7.94669e-10, 7.400306e-10, 
    9.610106e-10, 8.397558e-10, 1.035365e-09, 9.731753e-10, 9.316565e-10, 
    9.497064e-10, 8.587999e-10, 8.383694e-10, 7.591188e-10, 7.993422e-10, 
    5.821214e-10, 6.717652e-10, 4.459314e-10, 5.020087e-10, 1.034682e-09, 
    1.002809e-09, 8.976249e-10, 9.465738e-10, 8.117275e-10, 7.808978e-10, 
    7.565025e-10, 7.261611e-10, 7.229449e-10, 7.05471e-10, 7.34276e-10, 
    7.065937e-10, 8.1567e-10, 7.654521e-10, 9.092108e-10, 8.724764e-10, 
    8.892348e-10, 9.078925e-10, 8.51245e-10, 7.93881e-10, 7.926958e-10, 
    7.749587e-10, 7.265862e-10, 8.112129e-10, 5.712461e-10, 7.118036e-10, 
    9.689042e-10, 9.111292e-10, 9.031049e-10, 9.250182e-10, 7.839476e-10, 
    8.330235e-10, 7.058939e-10, 7.386843e-10, 6.855486e-10, 7.115737e-10, 
    7.154651e-10, 7.501337e-10, 7.723531e-10, 8.30722e-10, 8.806389e-10, 
    9.218163e-10, 9.121148e-10, 8.673219e-10, 7.904719e-10, 7.226509e-10, 
    7.371119e-10, 6.894812e-10, 8.209822e-10, 7.637053e-10, 7.854676e-10, 
    7.296901e-10, 8.560818e-10, 7.474694e-10, 8.856687e-10, 8.728332e-10, 
    8.340208e-10, 7.599288e-10, 7.442473e-10, 7.277645e-10, 7.379035e-10, 
    7.885923e-10, 7.971462e-10, 8.349502e-10, 8.456199e-10, 8.756162e-10, 
    9.010513e-10, 8.777885e-10, 8.5385e-10, 7.885734e-10, 7.330605e-10, 
    6.759882e-10, 6.625564e-10, 6.011919e-10, 6.50789e-10, 5.705271e-10, 
    6.38232e-10, 5.246346e-10, 7.415251e-10, 6.403249e-10, 8.32289e-10, 
    8.097367e-10, 7.701212e-10, 6.848525e-10, 7.299452e-10, 6.774287e-10, 
    7.974833e-10, 8.658028e-10, 8.841908e-10, 9.192705e-10, 8.834009e-10, 
    8.862783e-10, 8.528749e-10, 8.635035e-10, 7.864734e-10, 8.271709e-10, 
    7.155613e-10, 6.778334e-10, 5.794714e-10, 5.248372e-10, 4.733936e-10, 
    4.519595e-10, 4.455873e-10, 4.429438e-10,
  9.840423e-12, 8.887793e-12, 9.067056e-12, 8.341541e-12, 8.738133e-12, 
    8.271547e-12, 9.641117e-12, 8.851498e-12, 9.349444e-12, 9.751567e-12, 
    7.064608e-12, 8.310289e-12, 5.932419e-12, 6.609068e-12, 5.014919e-12, 
    6.033893e-12, 4.827144e-12, 5.042317e-12, 4.41693e-12, 4.5894e-12, 
    3.858774e-12, 4.339091e-12, 3.518469e-12, 3.969452e-12, 3.895997e-12, 
    4.355702e-12, 8.046718e-12, 7.211053e-12, 8.098509e-12, 7.974257e-12, 
    8.029842e-12, 8.72976e-12, 9.100194e-12, 9.916484e-12, 9.76418e-12, 
    9.16669e-12, 7.918881e-12, 8.326432e-12, 7.329839e-12, 7.351251e-12, 
    6.352966e-12, 6.788809e-12, 5.275961e-12, 5.675528e-12, 4.582097e-12, 
    4.839759e-12, 4.59394e-12, 4.667411e-12, 4.592989e-12, 4.975477e-12, 
    4.808614e-12, 5.156278e-12, 6.705417e-12, 6.216297e-12, 7.765002e-12, 
    8.833523e-12, 9.605343e-12, 1.018447e-11, 1.010097e-11, 9.943265e-12, 
    9.16328e-12, 8.474823e-12, 7.978109e-12, 7.658888e-12, 7.354332e-12, 
    6.490245e-12, 6.066826e-12, 5.197921e-12, 5.346978e-12, 5.096462e-12, 
    4.866013e-12, 4.497741e-12, 4.556786e-12, 4.400115e-12, 5.102989e-12, 
    4.626649e-12, 5.433375e-12, 5.202412e-12, 7.272931e-12, 8.214902e-12, 
    8.643058e-12, 9.032366e-12, 1.003713e-11, 9.334349e-12, 9.606591e-12, 
    8.969005e-12, 8.581508e-12, 8.771484e-12, 7.650304e-12, 8.071829e-12, 
    6.042435e-12, 6.859824e-12, 4.892456e-12, 5.316116e-12, 4.795023e-12, 
    5.055595e-12, 4.615724e-12, 5.010162e-12, 4.342928e-12, 4.207478e-12, 
    4.299666e-12, 3.954162e-12, 5.032781e-12, 4.593922e-12, 8.776839e-12, 
    8.745614e-12, 8.601332e-12, 9.249862e-12, 9.290771e-12, 9.920668e-12, 
    9.358628e-12, 9.127026e-12, 8.559483e-12, 8.237081e-12, 7.939593e-12, 
    7.315354e-12, 6.664744e-12, 5.832822e-12, 5.287797e-12, 4.94569e-12, 
    5.15332e-12, 4.969659e-12, 5.175312e-12, 5.274011e-12, 4.257818e-12, 
    4.807067e-12, 4.002445e-12, 4.043956e-12, 4.396435e-12, 4.039262e-12, 
    8.723745e-12, 8.904272e-12, 9.553943e-12, 9.04246e-12, 9.991251e-12, 
    9.450935e-12, 9.150834e-12, 8.062768e-12, 7.838103e-12, 7.634135e-12, 
    7.243701e-12, 6.76594e-12, 5.988367e-12, 5.371132e-12, 4.852874e-12, 
    4.889443e-12, 4.876542e-12, 4.765948e-12, 5.043591e-12, 4.721555e-12, 
    4.669131e-12, 4.807159e-12, 4.049541e-12, 4.255513e-12, 4.044842e-12, 
    4.177908e-12, 8.845279e-12, 8.544787e-12, 8.706137e-12, 8.404672e-12, 
    8.616156e-12, 7.706909e-12, 7.449647e-12, 6.334702e-12, 6.775083e-12, 
    6.085168e-12, 6.70232e-12, 6.589484e-12, 6.063538e-12, 6.667769e-12, 
    5.403746e-12, 6.237462e-12, 4.76169e-12, 5.51566e-12, 4.717324e-12, 
    4.855026e-12, 4.628756e-12, 4.433284e-12, 4.196801e-12, 3.786836e-12, 
    3.878804e-12, 3.554894e-12, 8.111871e-12, 7.749434e-12, 7.780876e-12, 
    7.41428e-12, 7.152048e-12, 6.608924e-12, 5.80649e-12, 6.098623e-12, 
    5.570981e-12, 5.469553e-12, 6.274754e-12, 5.769964e-12, 7.514154e-12, 
    7.207183e-12, 7.388771e-12, 8.082769e-12, 6.030229e-12, 7.024146e-12, 
    5.279135e-12, 5.750638e-12, 4.46074e-12, 5.069676e-12, 3.930178e-12, 
    3.510209e-12, 3.148578e-12, 2.764217e-12, 7.557162e-12, 7.797196e-12, 
    7.371625e-12, 6.813264e-12, 6.325805e-12, 5.720946e-12, 5.661773e-12, 
    5.554628e-12, 5.284618e-12, 5.065739e-12, 5.521045e-12, 5.01202e-12, 
    7.137324e-12, 5.949548e-12, 7.889447e-12, 7.259183e-12, 6.845241e-12, 
    7.024511e-12, 6.132752e-12, 5.936261e-12, 5.188538e-12, 5.56511e-12, 
    3.610336e-12, 4.392799e-12, 2.497604e-12, 2.943732e-12, 7.882455e-12, 
    7.558005e-12, 6.510184e-12, 6.993322e-12, 5.68229e-12, 5.391668e-12, 
    5.16426e-12, 4.884669e-12, 4.855248e-12, 4.696134e-12, 4.959088e-12, 
    4.70632e-12, 5.719709e-12, 5.247419e-12, 6.623816e-12, 6.26511e-12, 
    6.428179e-12, 6.610864e-12, 6.059919e-12, 5.513623e-12, 5.502464e-12, 
    5.336094e-12, 4.888561e-12, 5.67741e-12, 3.517952e-12, 4.753654e-12, 
    7.216343e-12, 6.642676e-12, 6.563874e-12, 6.77958e-12, 5.420258e-12, 
    5.885093e-12, 4.699971e-12, 4.999626e-12, 4.516264e-12, 4.751563e-12, 
    4.786986e-12, 5.10527e-12, 5.311755e-12, 5.863096e-12, 6.344415e-12, 
    6.747962e-12, 6.652368e-12, 6.215148e-12, 5.481539e-12, 4.852561e-12, 
    4.985157e-12, 4.551638e-12, 5.770219e-12, 5.231163e-12, 5.434521e-12, 
    4.917e-12, 6.106525e-12, 5.080641e-12, 6.393398e-12, 6.268571e-12, 
    5.894631e-12, 5.19606e-12, 5.050891e-12, 4.899353e-12, 4.99244e-12, 
    5.463868e-12, 5.544393e-12, 5.903522e-12, 6.005822e-12, 6.295588e-12, 
    6.543741e-12, 6.316695e-12, 6.08501e-12, 5.46369e-12, 4.947924e-12, 
    4.430541e-12, 4.310763e-12, 3.773707e-12, 4.206472e-12, 3.511865e-12, 
    4.095853e-12, 3.128653e-12, 5.025789e-12, 4.114241e-12, 5.878071e-12, 
    5.663416e-12, 5.290929e-12, 4.51001e-12, 4.919338e-12, 4.443431e-12, 
    5.547572e-12, 6.200443e-12, 6.378996e-12, 6.722847e-12, 6.371301e-12, 
    6.399341e-12, 6.075614e-12, 6.178198e-12, 5.443963e-12, 5.829193e-12, 
    4.787862e-12, 4.447055e-12, 3.587772e-12, 3.130322e-12, 2.713851e-12, 
    2.544694e-12, 2.494922e-12, 2.474346e-12,
  1.242757e-14, 1.029839e-14, 1.068943e-14, 9.135775e-15, 9.975472e-15, 
    8.990046e-15, 1.197188e-14, 1.021978e-14, 1.131462e-14, 1.222376e-14, 
    6.601605e-15, 9.070615e-15, 4.598079e-15, 5.765806e-15, 3.170908e-15, 
    4.767296e-15, 2.903251e-15, 3.210692e-15, 2.350116e-15, 2.577252e-15, 
    1.672596e-15, 2.250265e-15, 1.306043e-15, 1.799651e-15, 1.714909e-15, 
    2.271433e-15, 8.527096e-15, 6.87829e-15, 8.633039e-15, 8.379588e-15, 
    8.492667e-15, 9.957503e-15, 1.076222e-14, 1.260284e-14, 1.225263e-14, 
    1.090875e-14, 8.267422e-15, 9.104251e-15, 7.105476e-15, 7.146688e-15, 
    5.313116e-15, 6.091002e-15, 3.557311e-15, 4.179457e-15, 2.567472e-15, 
    2.920956e-15, 2.58334e-15, 2.682601e-15, 2.582064e-15, 3.113959e-15, 
    2.877318e-15, 3.378125e-15, 5.93937e-15, 5.076805e-15, 7.958334e-15, 
    1.018092e-14, 1.189065e-14, 1.322638e-14, 1.30311e-14, 1.266474e-14, 
    1.090122e-14, 9.415335e-15, 8.387406e-15, 7.747443e-15, 7.152627e-15, 
    5.554194e-15, 4.822673e-15, 3.440088e-15, 3.665227e-15, 3.289851e-15, 
    2.95793e-15, 2.455541e-15, 2.533688e-15, 2.328404e-15, 3.299442e-15, 
    2.627354e-15, 3.798085e-15, 3.446794e-15, 6.996332e-15, 8.872663e-15, 
    9.772036e-15, 1.06134e-14, 1.288241e-14, 1.128093e-14, 1.189349e-14, 
    1.047498e-14, 9.641042e-15, 1.004715e-14, 7.730464e-15, 8.57841e-15, 
    4.781637e-15, 6.221147e-15, 2.995348e-15, 3.618185e-15, 2.858354e-15, 
    3.230038e-15, 2.612622e-15, 3.164019e-15, 2.255149e-15, 2.085296e-15, 
    2.200336e-15, 1.781877e-15, 3.196824e-15, 2.583316e-15, 1.005867e-14, 
    9.991535e-15, 9.683171e-15, 1.109289e-14, 1.118381e-14, 1.261251e-14, 
    1.133514e-14, 1.082127e-14, 9.594306e-15, 8.918565e-15, 8.309314e-15, 
    7.077641e-15, 5.865889e-15, 4.4341e-15, 3.575215e-15, 3.071205e-15, 
    3.37374e-15, 3.105591e-15, 3.406396e-15, 3.554364e-15, 2.147815e-15, 
    2.875157e-15, 1.838244e-15, 1.887264e-15, 2.323663e-15, 1.881695e-15, 
    9.9446e-15, 1.033415e-14, 1.177424e-14, 1.063551e-14, 1.277587e-14, 
    1.154202e-14, 1.087375e-14, 8.559885e-15, 8.104687e-15, 7.698516e-15, 
    6.940482e-15, 6.04929e-15, 4.691112e-15, 3.702198e-15, 2.939404e-15, 
    2.991076e-15, 2.972809e-15, 2.81794e-15, 3.212545e-15, 2.756656e-15, 
    2.68494e-15, 2.875286e-15, 1.893898e-15, 2.144936e-15, 1.888316e-15, 
    2.04891e-15, 1.020633e-14, 9.563162e-15, 9.906861e-15, 9.267857e-15, 
    9.714713e-15, 7.842651e-15, 7.337095e-15, 5.281322e-15, 6.065954e-15, 
    4.853612e-15, 5.933764e-15, 5.730743e-15, 4.817135e-15, 5.871341e-15, 
    3.752331e-15, 5.113159e-15, 2.812041e-15, 3.926206e-15, 2.750841e-15, 
    2.942436e-15, 2.630198e-15, 2.371307e-15, 2.072128e-15, 1.592036e-15, 
    1.695312e-15, 1.343484e-15, 8.66044e-15, 7.927279e-15, 7.99004e-15, 
    7.268465e-15, 6.766348e-15, 5.765548e-15, 4.391099e-15, 4.876351e-15, 
    4.013198e-15, 3.854226e-15, 5.177425e-15, 4.331698e-15, 7.462817e-15, 
    6.870925e-15, 7.219098e-15, 8.600797e-15, 4.761147e-15, 6.52583e-15, 
    3.562109e-15, 4.300384e-15, 2.407049e-15, 3.250602e-15, 1.754139e-15, 
    1.297615e-15, 9.515462e-16, 6.360298e-16, 7.547027e-15, 8.022681e-15, 
    7.185979e-15, 6.135715e-15, 5.265857e-15, 4.252433e-15, 4.157444e-15, 
    3.98741e-15, 3.570403e-15, 3.244846e-15, 3.934643e-15, 3.16671e-15, 
    6.738515e-15, 4.626492e-15, 8.208003e-15, 6.970044e-15, 6.194346e-15, 
    6.52651e-15, 4.934199e-15, 4.604445e-15, 3.42609e-15, 4.003933e-15, 
    1.401315e-15, 2.318982e-15, 4.515406e-16, 7.763729e-16, 8.193907e-15, 
    7.548681e-15, 5.589513e-15, 6.468301e-15, 4.190293e-15, 3.733736e-15, 
    3.38997e-15, 2.984311e-15, 2.942748e-15, 2.721792e-15, 3.090409e-15, 
    2.735742e-15, 4.250441e-15, 3.514271e-15, 5.792258e-15, 5.160778e-15, 
    5.444741e-15, 5.769024e-15, 4.811039e-15, 3.923015e-15, 3.905554e-15, 
    3.648611e-15, 2.989827e-15, 4.182472e-15, 1.305515e-15, 2.800918e-15, 
    6.888348e-15, 5.826149e-15, 5.685e-15, 6.074156e-15, 3.777805e-15, 
    4.519897e-15, 2.727043e-15, 3.148781e-15, 2.479955e-15, 2.798026e-15, 
    2.847161e-15, 3.302796e-15, 3.611556e-15, 4.483722e-15, 5.298221e-15, 
    6.016566e-15, 5.84359e-15, 5.074836e-15, 3.872892e-15, 2.938964e-15, 
    3.1279e-15, 2.526837e-15, 4.332111e-15, 3.489845e-15, 3.79986e-15, 
    3.030234e-15, 4.889724e-15, 3.266649e-15, 5.383735e-15, 5.16675e-15, 
    4.535615e-15, 3.437309e-15, 3.22318e-15, 3.005135e-15, 3.138404e-15, 
    3.845385e-15, 3.971303e-15, 4.550285e-15, 4.720269e-15, 5.213451e-15, 
    5.649129e-15, 5.250037e-15, 4.853345e-15, 3.845109e-15, 3.074405e-15, 
    2.367748e-15, 2.214345e-15, 1.577508e-15, 2.084053e-15, 1.299302e-15, 
    1.949268e-15, 9.338249e-16, 3.186671e-15, 1.971426e-15, 4.508337e-15, 
    4.160072e-15, 3.579958e-15, 2.471701e-15, 3.033567e-15, 2.384493e-15, 
    3.976303e-15, 5.049636e-15, 5.358543e-15, 5.970955e-15, 5.345101e-15, 
    5.394141e-15, 4.837488e-15, 5.011597e-15, 3.814486e-15, 4.428164e-15, 
    2.84838e-15, 2.389209e-15, 1.377657e-15, 9.353039e-16, 5.989441e-16, 
    4.819759e-16, 4.498357e-16, 4.368566e-16,
  4.204027e-20, 3.491363e-20, 3.622382e-20, 3.101438e-20, 3.38312e-20, 
    3.052519e-20, 4.051648e-20, 3.465017e-20, 3.831726e-20, 4.135884e-20, 
    2.249192e-20, 3.079566e-20, 1.572527e-20, 1.967273e-20, 1.088431e-20, 
    1.6298e-20, 9.97377e-21, 1.101956e-20, 8.088746e-21, 8.863382e-21, 
    5.772404e-21, 7.74793e-21, 4.514845e-21, 6.207517e-21, 5.917352e-21, 
    7.820194e-21, 2.897047e-20, 2.342417e-20, 2.932635e-20, 2.847488e-20, 
    2.885481e-20, 3.377095e-20, 3.646764e-20, 4.262621e-20, 4.145536e-20, 
    3.695836e-20, 2.809795e-20, 3.090857e-20, 2.41893e-20, 2.432807e-20, 
    1.814372e-20, 2.077019e-20, 1.219717e-20, 1.43074e-20, 8.830046e-21, 
    1.003403e-20, 8.884131e-21, 9.222388e-21, 8.879783e-21, 1.069065e-20, 
    9.885497e-21, 1.158859e-20, 2.025856e-20, 1.734492e-20, 2.705894e-20, 
    3.451992e-20, 4.024476e-20, 4.470975e-20, 4.405738e-20, 4.283309e-20, 
    3.693315e-20, 3.195254e-20, 2.850115e-20, 2.634973e-20, 2.434807e-20, 
    1.895818e-20, 1.648537e-20, 1.179908e-20, 1.256351e-20, 1.128863e-20, 
    1.015986e-20, 8.448396e-21, 8.714873e-21, 8.014652e-21, 1.132123e-20, 
    9.03414e-21, 1.301434e-20, 1.182186e-20, 2.382177e-20, 3.013109e-20, 
    3.314905e-20, 3.596913e-20, 4.356054e-20, 3.820447e-20, 4.025423e-20, 
    3.550536e-20, 3.270971e-20, 3.40715e-20, 2.629261e-20, 2.914285e-20, 
    1.634652e-20, 2.12092e-20, 1.028718e-20, 1.240383e-20, 9.820938e-21, 
    1.108533e-20, 8.983934e-21, 1.086088e-20, 7.764604e-21, 7.184452e-21, 
    7.577441e-21, 6.146668e-21, 1.097242e-20, 8.884049e-21, 3.411014e-20, 
    3.388505e-20, 3.285101e-20, 3.757496e-20, 3.787937e-20, 4.265851e-20, 
    3.838594e-20, 3.66654e-20, 3.255294e-20, 3.028521e-20, 2.823874e-20, 
    2.409558e-20, 2.001057e-20, 1.517002e-20, 1.225796e-20, 1.054524e-20, 
    1.157369e-20, 1.06622e-20, 1.168463e-20, 1.218716e-20, 7.398056e-21, 
    9.878142e-21, 6.339608e-21, 6.507344e-21, 7.998471e-21, 6.48829e-21, 
    3.372769e-20, 3.503345e-20, 3.985532e-20, 3.604318e-20, 4.320452e-20, 
    3.907831e-20, 3.684117e-20, 2.908062e-20, 2.755097e-20, 2.618515e-20, 
    2.363366e-20, 2.062947e-20, 1.604017e-20, 1.268898e-20, 1.009682e-20, 
    1.027265e-20, 1.021049e-20, 9.683345e-21, 1.102586e-20, 9.474647e-21, 
    9.230357e-21, 9.87858e-21, 6.53004e-21, 7.388222e-21, 6.510943e-21, 
    7.060099e-21, 3.460508e-20, 3.244847e-20, 3.360116e-20, 3.145767e-20, 
    3.29568e-20, 2.666993e-20, 2.496905e-20, 1.803627e-20, 2.068569e-20, 
    1.659004e-20, 2.023965e-20, 1.955436e-20, 1.646663e-20, 2.002897e-20, 
    1.28591e-20, 1.746783e-20, 9.663256e-21, 1.344891e-20, 9.454843e-21, 
    1.010713e-20, 9.043832e-21, 8.161052e-21, 7.139455e-21, 5.496323e-21, 
    5.850226e-21, 4.643466e-21, 2.941839e-20, 2.695451e-20, 2.716554e-20, 
    2.473804e-20, 2.304706e-20, 1.967186e-20, 1.502438e-20, 1.666697e-20, 
    1.374388e-20, 1.320478e-20, 1.76851e-20, 1.482316e-20, 2.539216e-20, 
    2.339937e-20, 2.457185e-20, 2.921805e-20, 1.627719e-20, 2.223652e-20, 
    1.221346e-20, 1.47171e-20, 8.282992e-21, 1.115523e-20, 6.051697e-21, 
    4.485883e-21, 3.294765e-21, 2.204597e-21, 2.567551e-20, 2.727529e-20, 
    2.446035e-20, 2.092103e-20, 1.7984e-20, 1.455466e-20, 1.423281e-20, 
    1.365644e-20, 1.224162e-20, 1.113567e-20, 1.347752e-20, 1.087003e-20, 
    2.295328e-20, 1.582145e-20, 2.789825e-20, 2.373323e-20, 2.11188e-20, 
    2.223881e-20, 1.686265e-20, 1.574682e-20, 1.175153e-20, 1.371247e-20, 
    4.84205e-21, 7.982496e-21, 1.564588e-21, 2.690079e-21, 2.785087e-20, 
    2.568108e-20, 1.907746e-20, 2.204259e-20, 1.434412e-20, 1.279601e-20, 
    1.162883e-20, 1.024963e-20, 1.01082e-20, 9.355897e-21, 1.061056e-20, 
    9.403413e-21, 1.454791e-20, 1.205102e-20, 1.976203e-20, 1.762882e-20, 
    1.858846e-20, 1.968359e-20, 1.644601e-20, 1.343809e-20, 1.337887e-20, 
    1.250711e-20, 1.02684e-20, 1.431761e-20, 4.51303e-21, 9.625384e-21, 
    2.345806e-20, 1.987643e-20, 1.939991e-20, 2.071336e-20, 1.294553e-20, 
    1.546057e-20, 9.373783e-21, 1.080907e-20, 8.531659e-21, 9.615536e-21, 
    9.782832e-21, 1.133262e-20, 1.238133e-20, 1.533807e-20, 1.809338e-20, 
    2.051906e-20, 1.99353e-20, 1.733826e-20, 1.32681e-20, 1.009532e-20, 
    1.073806e-20, 8.691515e-21, 1.482456e-20, 1.196807e-20, 1.302036e-20, 
    1.040587e-20, 1.671221e-20, 1.120977e-20, 1.838234e-20, 1.764901e-20, 
    1.551379e-20, 1.178964e-20, 1.106201e-20, 1.032048e-20, 1.077378e-20, 
    1.317479e-20, 1.360183e-20, 1.556346e-20, 1.613885e-20, 1.780688e-20, 
    1.927879e-20, 1.793053e-20, 1.658914e-20, 1.317386e-20, 1.055613e-20, 
    8.148907e-21, 7.625283e-21, 5.446519e-21, 7.180206e-21, 4.491682e-21, 
    6.719432e-21, 3.233653e-21, 1.09379e-20, 6.795208e-21, 1.542142e-20, 
    1.424171e-20, 1.227406e-20, 8.503511e-21, 1.041721e-20, 8.206042e-21, 
    1.361879e-20, 1.725305e-20, 1.829722e-20, 2.036515e-20, 1.82518e-20, 
    1.84175e-20, 1.653549e-20, 1.712442e-20, 1.306998e-20, 1.514992e-20, 
    9.786984e-21, 8.222131e-21, 4.760825e-21, 3.238754e-21, 2.076125e-21, 
    1.670337e-21, 1.558662e-21, 1.513542e-21,
  3.086726e-26, 2.565605e-26, 2.661439e-26, 2.28031e-26, 2.486421e-26, 
    2.244508e-26, 2.975332e-26, 2.546333e-26, 2.814535e-26, 3.036913e-26, 
    1.656212e-26, 2.264303e-26, 1.159973e-26, 1.449558e-26, 8.043276e-27, 
    1.202007e-26, 7.373578e-27, 8.142735e-27, 5.986152e-27, 6.55648e-27, 
    4.278932e-27, 5.73514e-27, 3.350597e-27, 4.599864e-27, 4.385857e-27, 
    5.788367e-27, 2.130709e-26, 1.724523e-26, 2.15676e-26, 2.094427e-26, 
    2.122242e-26, 2.482013e-26, 2.679271e-26, 3.129555e-26, 3.043969e-26, 
    2.71516e-26, 2.066832e-26, 2.272567e-26, 1.78058e-26, 1.790746e-26, 
    1.337424e-26, 1.530019e-26, 9.008419e-27, 1.055875e-26, 6.531942e-27, 
    7.417909e-27, 6.571754e-27, 6.820713e-27, 6.568553e-27, 7.900868e-27, 
    7.308638e-27, 8.561088e-27, 1.492511e-26, 1.278826e-26, 1.990756e-26, 
    2.536805e-26, 2.955467e-26, 3.281835e-26, 3.234159e-26, 3.144677e-26, 
    2.713316e-26, 2.348965e-26, 2.096351e-26, 1.938822e-26, 1.79221e-26, 
    1.39716e-26, 1.215757e-26, 8.715819e-27, 9.277641e-27, 8.340569e-27, 
    7.510471e-27, 6.250979e-27, 6.447161e-27, 5.931587e-27, 8.364533e-27, 
    6.682166e-27, 9.608907e-27, 8.732562e-27, 1.753654e-26, 2.215664e-26, 
    2.436513e-26, 2.642811e-26, 3.197847e-26, 2.806287e-26, 2.956159e-26, 
    2.608889e-26, 2.404368e-26, 2.504001e-26, 1.934639e-26, 2.143327e-26, 
    1.205568e-26, 1.5622e-26, 7.604125e-27, 9.1603e-27, 7.261142e-27, 
    8.191092e-27, 6.645214e-27, 8.026051e-27, 5.747422e-27, 5.32001e-27, 
    5.609553e-27, 4.55499e-27, 8.108067e-27, 6.571693e-27, 2.506827e-26, 
    2.490361e-26, 2.414707e-26, 2.760253e-26, 2.782514e-26, 3.131916e-26, 
    2.819557e-26, 2.693735e-26, 2.392898e-26, 2.226944e-26, 2.077139e-26, 
    1.773714e-26, 1.474329e-26, 1.119215e-26, 9.053095e-27, 7.793929e-27, 
    8.550136e-27, 7.879941e-27, 8.631692e-27, 9.001065e-27, 5.477397e-27, 
    7.303226e-27, 4.697267e-27, 4.82094e-27, 5.91967e-27, 4.806893e-27, 
    2.478848e-26, 2.57437e-26, 2.926994e-26, 2.648227e-26, 3.171825e-26, 
    2.870183e-26, 2.706589e-26, 2.138772e-26, 2.026784e-26, 1.926769e-26, 
    1.739872e-26, 1.519703e-26, 1.183085e-26, 9.369845e-27, 7.464095e-27, 
    7.593433e-27, 7.547713e-27, 7.15991e-27, 8.147367e-27, 7.006348e-27, 
    6.826579e-27, 7.303549e-27, 4.837673e-27, 5.470152e-27, 4.823593e-27, 
    5.228374e-27, 2.543034e-26, 2.385254e-26, 2.469591e-26, 2.312751e-26, 
    2.422448e-26, 1.962271e-26, 1.8377e-26, 1.329543e-26, 1.523825e-26, 
    1.223438e-26, 1.491124e-26, 1.440878e-26, 1.214382e-26, 1.475678e-26, 
    9.494848e-27, 1.287843e-26, 7.145128e-27, 9.928174e-27, 6.991776e-27, 
    7.471684e-27, 6.689301e-27, 6.0394e-27, 5.286852e-27, 4.075233e-27, 
    4.336342e-27, 3.445606e-27, 2.163497e-26, 1.98311e-26, 1.998562e-26, 
    1.820778e-26, 1.696891e-26, 1.449494e-26, 1.108522e-26, 1.229083e-26, 
    1.014485e-26, 9.748828e-27, 1.303782e-26, 1.09375e-26, 1.868691e-26, 
    1.722706e-26, 1.808604e-26, 2.148832e-26, 1.200479e-26, 1.637495e-26, 
    9.02039e-27, 1.085961e-26, 6.129192e-27, 8.242486e-27, 4.484948e-27, 
    3.329202e-27, 2.448524e-27, 1.640798e-27, 1.889445e-26, 2.006598e-26, 
    1.800436e-26, 1.541077e-26, 1.325709e-26, 1.074033e-26, 1.050396e-26, 
    1.008063e-26, 9.041086e-27, 8.228104e-27, 9.949192e-27, 8.03278e-27, 
    1.69002e-26, 1.167032e-26, 2.052211e-26, 1.747167e-26, 1.555574e-26, 
    1.637663e-26, 1.243441e-26, 1.161554e-26, 8.680869e-27, 1.012178e-26, 
    3.592265e-27, 5.907905e-27, 1.165494e-27, 2.000755e-27, 2.048742e-26, 
    1.889852e-26, 1.405907e-26, 1.623283e-26, 1.058571e-26, 9.448487e-27, 
    8.590669e-27, 7.576501e-27, 7.472466e-27, 6.918964e-27, 7.841965e-27, 
    6.953931e-27, 1.073537e-26, 8.901007e-27, 1.456106e-26, 1.299654e-26, 
    1.370044e-26, 1.450355e-26, 1.212868e-26, 9.920224e-27, 9.876723e-27, 
    9.236198e-27, 7.590309e-27, 1.056625e-26, 3.349257e-27, 7.117263e-27, 
    1.727006e-26, 1.464494e-26, 1.429553e-26, 1.525853e-26, 9.558353e-27, 
    1.140543e-26, 6.932127e-27, 7.987949e-27, 6.31228e-27, 7.110017e-27, 
    7.233106e-27, 8.372913e-27, 9.143763e-27, 1.131551e-26, 1.333732e-26, 
    1.511609e-26, 1.46881e-26, 1.278337e-26, 9.795341e-27, 7.462992e-27, 
    7.935733e-27, 6.429966e-27, 1.093853e-26, 8.840037e-27, 9.613329e-27, 
    7.691425e-27, 1.232402e-26, 8.28259e-27, 1.354927e-26, 1.301135e-26, 
    1.14445e-26, 8.708883e-27, 8.173949e-27, 7.628619e-27, 7.962002e-27, 
    9.726794e-27, 1.004051e-26, 1.148096e-26, 1.190327e-26, 1.312715e-26, 
    1.420671e-26, 1.321787e-26, 1.223372e-26, 9.726107e-27, 7.801933e-27, 
    6.030456e-27, 5.644796e-27, 4.03848e-27, 5.316881e-27, 3.333486e-27, 
    4.97729e-27, 2.403294e-27, 8.082684e-27, 5.033145e-27, 1.13767e-26, 
    1.05105e-26, 9.064928e-27, 6.291557e-27, 7.699762e-27, 6.07253e-27, 
    1.005297e-26, 1.272085e-26, 1.348683e-26, 1.500325e-26, 1.345352e-26, 
    1.357506e-26, 1.219435e-26, 1.262648e-26, 9.649786e-27, 1.117739e-26, 
    7.23616e-27, 6.084377e-27, 3.532282e-27, 2.407069e-27, 1.545465e-27, 
    1.244101e-27, 1.161089e-27, 1.127538e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004395003, 0.004392459, 0.004392955, 0.0043909, 0.004392041, 0.004390695, 
    0.004394489, 0.004392356, 0.004393719, 0.004394777, 0.004386907, 
    0.004390809, 0.004382877, 0.004385361, 0.004379131, 0.00438326, 
    0.0043783, 0.004379255, 0.004376392, 0.004377213, 0.004373542, 
    0.004376014, 0.004371648, 0.004374135, 0.004373744, 0.004376095, 
    0.004390028, 0.00438739, 0.004390183, 0.004389808, 0.004389978, 
    0.004392016, 0.00439304, 0.004395201, 0.00439481, 0.004393225, 
    0.004389639, 0.00439086, 0.004387793, 0.004387863, 0.004384447, 
    0.004385986, 0.004380254, 0.004381883, 0.004377179, 0.004378361, 
    0.004377233, 0.004377576, 0.004377229, 0.004378963, 0.00437822, 
    0.004379747, 0.004385697, 0.004383946, 0.004389167, 0.004392301, 
    0.004394395, 0.004395877, 0.004395668, 0.004395267, 0.004393215, 
    0.004391291, 0.004389822, 0.00438884, 0.004387872, 0.004384932, 
    0.004383387, 0.004379922, 0.004380551, 0.004379488, 0.004378479, 
    0.004376778, 0.004377059, 0.004376309, 0.004379519, 0.004377384, 
    0.004380909, 0.004379944, 0.004387592, 0.004390531, 0.004391765, 
    0.004392859, 0.004395506, 0.004393677, 0.004394398, 0.004392687, 
    0.004391597, 0.004392137, 0.004388813, 0.004390105, 0.004383295, 
    0.004386227, 0.004378596, 0.004380422, 0.00437816, 0.004379315, 
    0.004377334, 0.004379116, 0.004376031, 0.004375358, 0.004375818, 
    0.004374058, 0.004379215, 0.004377231, 0.004392151, 0.004392063, 
    0.004391654, 0.00439345, 0.00439356, 0.004395211, 0.004393744, 
    0.004393118, 0.004391535, 0.004390596, 0.004389705, 0.004387744, 
    0.004385553, 0.004382496, 0.004380303, 0.004378833, 0.004379736, 
    0.004378939, 0.004379829, 0.004380248, 0.004375609, 0.004378212, 
    0.00437431, 0.004374527, 0.00437629, 0.004374503, 0.004392001, 
    0.004392507, 0.004394261, 0.004392889, 0.004395391, 0.004393988, 
    0.00439318, 0.004390074, 0.004389395, 0.004388761, 0.004387512, 
    0.004385908, 0.004383094, 0.004380649, 0.004378421, 0.004378584, 
    0.004378526, 0.004378027, 0.004379262, 0.004377824, 0.004377582, 
    0.004378214, 0.004374556, 0.004375601, 0.004374532, 0.004375212, 
    0.004392344, 0.004391492, 0.004391952, 0.004391087, 0.004391695, 
    0.004388985, 0.004388172, 0.004384377, 0.004385938, 0.004383458, 
    0.004385688, 0.004385292, 0.00438337, 0.004385568, 0.00438078, 
    0.004384019, 0.004378008, 0.004381234, 0.004377805, 0.00437843, 
    0.004377397, 0.00437647, 0.004375307, 0.004373157, 0.004373655, 
    0.004371861, 0.004390225, 0.004389119, 0.004389219, 0.004388065, 
    0.00438721, 0.004385362, 0.004382396, 0.004383512, 0.004381467, 
    0.004381055, 0.004384165, 0.004382252, 0.004388381, 0.004387387, 
    0.004387981, 0.004390135, 0.004383251, 0.004386781, 0.004380267, 
    0.004382179, 0.004376601, 0.004379371, 0.004373929, 0.004371596, 
    0.004369417, 0.004366853, 0.004388519, 0.00438927, 0.004387928, 
    0.004386066, 0.004384349, 0.004382061, 0.004381829, 0.0043814, 
    0.004380292, 0.004379359, 0.004381261, 0.004379125, 0.00438715, 
    0.004382946, 0.004389551, 0.004387557, 0.004386178, 0.004386786, 
    0.00438364, 0.004382899, 0.004379882, 0.004381443, 0.004372169, 
    0.004376269, 0.004364914, 0.004368082, 0.004389531, 0.004388523, 
    0.00438501, 0.004386682, 0.00438191, 0.004380735, 0.004379783, 
    0.00437856, 0.004378431, 0.004377707, 0.004378892, 0.004377755, 
    0.004382056, 0.004380134, 0.004385415, 0.004384127, 0.004384721, 
    0.004385369, 0.004383367, 0.00438123, 0.00438119, 0.004380504, 
    0.004378561, 0.004381891, 0.00437163, 0.004377955, 0.004387423, 
    0.004385474, 0.004385203, 0.004385956, 0.004380853, 0.004382701, 
    0.004377725, 0.004379071, 0.004376868, 0.004377962, 0.004378123, 
    0.00437953, 0.004380404, 0.004382615, 0.004384416, 0.004385848, 
    0.004385515, 0.004383943, 0.004381101, 0.004378417, 0.004379004, 
    0.004377035, 0.004382256, 0.004380064, 0.004380909, 0.004378706, 
    0.004383541, 0.004379407, 0.004384596, 0.004384142, 0.004382737, 
    0.004379911, 0.004379294, 0.004378626, 0.004379039, 0.004381029, 
    0.004381358, 0.004382773, 0.004383161, 0.004384241, 0.004385133, 
    0.004384317, 0.004383459, 0.004381031, 0.004378841, 0.004376456, 
    0.004375875, 0.004373077, 0.004375346, 0.004371594, 0.004374773, 
    0.004369277, 0.004379175, 0.004374878, 0.004382675, 0.004381836, 
    0.004380313, 0.004376831, 0.004378716, 0.004376514, 0.004381371, 
    0.004383886, 0.004384543, 0.00438576, 0.004384516, 0.004384617, 
    0.004383427, 0.004383809, 0.00438095, 0.004382486, 0.004378125, 
    0.004376533, 0.004372047, 0.004369296, 0.004366505, 0.004365271, 
    0.004364896, 0.004364739,
  8.322729e-06, 8.322773e-06, 8.322771e-06, 8.322805e-06, 8.322788e-06, 
    8.322892e-06, 8.32275e-06, 8.322766e-06, 8.322763e-06, 8.322748e-06, 
    8.324379e-06, 8.322845e-06, 8.326019e-06, 8.325065e-06, 8.32745e-06, 
    8.325857e-06, 8.327767e-06, 8.32743e-06, 8.328498e-06, 8.328196e-06, 
    8.329477e-06, 8.328636e-06, 8.330163e-06, 8.329292e-06, 8.32942e-06, 
    8.328604e-06, 8.323182e-06, 8.324184e-06, 8.323116e-06, 8.323262e-06, 
    8.323202e-06, 8.32278e-06, 8.322747e-06, 8.322741e-06, 8.322747e-06, 
    8.32276e-06, 8.323328e-06, 8.322841e-06, 8.324105e-06, 8.324077e-06, 
    8.325429e-06, 8.324824e-06, 8.327053e-06, 8.326437e-06, 8.328209e-06, 
    8.327767e-06, 8.328184e-06, 8.328061e-06, 8.328186e-06, 8.327537e-06, 
    8.327816e-06, 8.327248e-06, 8.324933e-06, 8.325619e-06, 8.323529e-06, 
    8.322743e-06, 8.322746e-06, 8.322723e-06, 8.322727e-06, 8.322729e-06, 
    8.32276e-06, 8.322799e-06, 8.323274e-06, 8.323676e-06, 8.324073e-06, 
    8.325189e-06, 8.325821e-06, 8.327164e-06, 8.326946e-06, 8.327331e-06, 
    8.327725e-06, 8.328348e-06, 8.328249e-06, 8.328517e-06, 8.327336e-06, 
    8.328117e-06, 8.326816e-06, 8.327174e-06, 8.324098e-06, 8.322977e-06, 
    8.322755e-06, 8.32277e-06, 8.322728e-06, 8.322754e-06, 8.322743e-06, 
    8.322784e-06, 8.322794e-06, 8.322793e-06, 8.323687e-06, 8.323154e-06, 
    8.325858e-06, 8.324714e-06, 8.327679e-06, 8.326992e-06, 8.327845e-06, 
    8.327416e-06, 8.32814e-06, 8.327489e-06, 8.328623e-06, 8.328856e-06, 
    8.328695e-06, 8.329336e-06, 8.327451e-06, 8.328177e-06, 8.32279e-06, 
    8.322789e-06, 8.322797e-06, 8.322756e-06, 8.322758e-06, 8.322737e-06, 
    8.322763e-06, 8.322766e-06, 8.322801e-06, 8.322949e-06, 8.323316e-06, 
    8.324116e-06, 8.324979e-06, 8.32618e-06, 8.327036e-06, 8.327596e-06, 
    8.32726e-06, 8.327556e-06, 8.327221e-06, 8.327067e-06, 8.328763e-06, 
    8.327813e-06, 8.329244e-06, 8.32917e-06, 8.32852e-06, 8.329178e-06, 
    8.322791e-06, 8.322789e-06, 8.322751e-06, 8.322781e-06, 8.322735e-06, 
    8.322753e-06, 8.322755e-06, 8.323147e-06, 8.323449e-06, 8.323701e-06, 
    8.324215e-06, 8.324855e-06, 8.325952e-06, 8.326896e-06, 8.327751e-06, 
    8.32769e-06, 8.327711e-06, 8.327891e-06, 8.327432e-06, 8.327966e-06, 
    8.328047e-06, 8.327823e-06, 8.329159e-06, 8.328783e-06, 8.329168e-06, 
    8.328926e-06, 8.322791e-06, 8.322797e-06, 8.322792e-06, 8.322795e-06, 
    8.322787e-06, 8.32359e-06, 8.323916e-06, 8.325434e-06, 8.324838e-06, 
    8.325806e-06, 8.324944e-06, 8.325093e-06, 8.325802e-06, 8.324996e-06, 
    8.326829e-06, 8.325564e-06, 8.327898e-06, 8.326635e-06, 8.327974e-06, 
    8.327746e-06, 8.32813e-06, 8.32846e-06, 8.328888e-06, 8.329639e-06, 
    8.32947e-06, 8.330103e-06, 8.323105e-06, 8.323546e-06, 8.323523e-06, 
    8.323991e-06, 8.32433e-06, 8.325077e-06, 8.32623e-06, 8.325805e-06, 
    8.3266e-06, 8.326751e-06, 8.325553e-06, 8.326278e-06, 8.32385e-06, 
    8.324235e-06, 8.324018e-06, 8.323131e-06, 8.325882e-06, 8.324481e-06, 
    8.327048e-06, 8.326318e-06, 8.328411e-06, 8.327369e-06, 8.329373e-06, 
    8.330157e-06, 8.33095e-06, 8.331769e-06, 8.323802e-06, 8.323503e-06, 
    8.32405e-06, 8.32477e-06, 8.32547e-06, 8.32636e-06, 8.326459e-06, 
    8.326619e-06, 8.327049e-06, 8.327398e-06, 8.326654e-06, 8.327487e-06, 
    8.324293e-06, 8.326008e-06, 8.323374e-06, 8.324163e-06, 8.324734e-06, 
    8.3245e-06, 8.32576e-06, 8.326047e-06, 8.327183e-06, 8.326609e-06, 
    8.329951e-06, 8.328508e-06, 8.33243e-06, 8.33137e-06, 8.323394e-06, 
    8.323808e-06, 8.325198e-06, 8.324545e-06, 8.326428e-06, 8.326871e-06, 
    8.327242e-06, 8.327685e-06, 8.327744e-06, 8.328006e-06, 8.327574e-06, 
    8.327995e-06, 8.326362e-06, 8.327102e-06, 8.32506e-06, 8.325557e-06, 
    8.325334e-06, 8.325078e-06, 8.325865e-06, 8.326661e-06, 8.326704e-06, 
    8.326952e-06, 8.327595e-06, 8.326435e-06, 8.330087e-06, 8.327833e-06, 
    8.324254e-06, 8.324999e-06, 8.325135e-06, 8.324843e-06, 8.326826e-06, 
    8.326115e-06, 8.328003e-06, 8.327507e-06, 8.328322e-06, 8.327917e-06, 
    8.327856e-06, 8.327334e-06, 8.327e-06, 8.326143e-06, 8.325441e-06, 
    8.324889e-06, 8.32502e-06, 8.325625e-06, 8.326716e-06, 8.327738e-06, 
    8.327513e-06, 8.328261e-06, 8.326292e-06, 8.327118e-06, 8.326792e-06, 
    8.327639e-06, 8.325788e-06, 8.327293e-06, 8.325384e-06, 8.325561e-06, 
    8.326101e-06, 8.327156e-06, 8.327423e-06, 8.32766e-06, 8.327519e-06, 
    8.326748e-06, 8.326631e-06, 8.326094e-06, 8.325932e-06, 8.325525e-06, 
    8.325172e-06, 8.325488e-06, 8.325812e-06, 8.326759e-06, 8.327578e-06, 
    8.328461e-06, 8.328684e-06, 8.329622e-06, 8.328826e-06, 8.330094e-06, 
    8.328966e-06, 8.330921e-06, 8.327415e-06, 8.328984e-06, 8.326134e-06, 
    8.326458e-06, 8.327011e-06, 8.328298e-06, 8.327635e-06, 8.328422e-06, 
    8.326629e-06, 8.325633e-06, 8.325403e-06, 8.324918e-06, 8.325414e-06, 
    8.325374e-06, 8.325843e-06, 8.325695e-06, 8.32679e-06, 8.326207e-06, 
    8.327847e-06, 8.328422e-06, 8.330027e-06, 8.330961e-06, 8.331923e-06, 
    8.332326e-06, 8.332449e-06, 8.332499e-06,
  1.678844e-10, 1.679383e-10, 1.679279e-10, 1.679826e-10, 1.679474e-10, 
    1.679914e-10, 1.678956e-10, 1.679401e-10, 1.679118e-10, 1.678897e-10, 
    1.681511e-10, 1.679865e-10, 1.68326e-10, 1.682199e-10, 1.684879e-10, 
    1.68309e-10, 1.685242e-10, 1.684835e-10, 1.686079e-10, 1.685723e-10, 
    1.687302e-10, 1.686244e-10, 1.688136e-10, 1.687053e-10, 1.68722e-10, 
    1.686207e-10, 1.680203e-10, 1.681304e-10, 1.680136e-10, 1.680293e-10, 
    1.680225e-10, 1.679477e-10, 1.679253e-10, 1.678808e-10, 1.67889e-10, 
    1.679219e-10, 1.680364e-10, 1.67985e-10, 1.681162e-10, 1.681132e-10, 
    1.682593e-10, 1.681933e-10, 1.684403e-10, 1.683701e-10, 1.685738e-10, 
    1.685223e-10, 1.685712e-10, 1.685565e-10, 1.685714e-10, 1.684961e-10, 
    1.685283e-10, 1.684623e-10, 1.682055e-10, 1.682806e-10, 1.680568e-10, 
    1.679405e-10, 1.678974e-10, 1.678665e-10, 1.678709e-10, 1.67879e-10, 
    1.679221e-10, 1.679703e-10, 1.680294e-10, 1.680713e-10, 1.681128e-10, 
    1.682367e-10, 1.683041e-10, 1.684541e-10, 1.684276e-10, 1.68473e-10, 
    1.685173e-10, 1.685908e-10, 1.685788e-10, 1.686111e-10, 1.684723e-10, 
    1.685643e-10, 1.684124e-10, 1.684538e-10, 1.681215e-10, 1.67999e-10, 
    1.679538e-10, 1.679298e-10, 1.678742e-10, 1.679124e-10, 1.678972e-10, 
    1.679339e-10, 1.679605e-10, 1.679456e-10, 1.680725e-10, 1.680172e-10, 
    1.68308e-10, 1.681825e-10, 1.685121e-10, 1.684331e-10, 1.685311e-10, 
    1.684812e-10, 1.685666e-10, 1.684898e-10, 1.686234e-10, 1.686522e-10, 
    1.686324e-10, 1.687093e-10, 1.684854e-10, 1.68571e-10, 1.679452e-10, 
    1.67947e-10, 1.679588e-10, 1.679172e-10, 1.679149e-10, 1.678805e-10, 
    1.679113e-10, 1.679243e-10, 1.679627e-10, 1.679962e-10, 1.680342e-10, 
    1.681179e-10, 1.682113e-10, 1.683429e-10, 1.684382e-10, 1.68502e-10, 
    1.684631e-10, 1.684975e-10, 1.684589e-10, 1.68441e-10, 1.686412e-10, 
    1.685284e-10, 1.686982e-10, 1.686889e-10, 1.686118e-10, 1.6869e-10, 
    1.679484e-10, 1.679378e-10, 1.679003e-10, 1.679296e-10, 1.678768e-10, 
    1.67906e-10, 1.679226e-10, 1.680178e-10, 1.680476e-10, 1.680744e-10, 
    1.681281e-10, 1.681967e-10, 1.683173e-10, 1.68423e-10, 1.685199e-10, 
    1.685129e-10, 1.685154e-10, 1.685368e-10, 1.684834e-10, 1.685456e-10, 
    1.685558e-10, 1.685287e-10, 1.686876e-10, 1.686422e-10, 1.686887e-10, 
    1.686592e-10, 1.679413e-10, 1.679639e-10, 1.679495e-10, 1.679766e-10, 
    1.679572e-10, 1.680641e-10, 1.680987e-10, 1.682615e-10, 1.681952e-10, 
    1.683015e-10, 1.682062e-10, 1.682229e-10, 1.683039e-10, 1.682115e-10, 
    1.684166e-10, 1.682765e-10, 1.685376e-10, 1.683963e-10, 1.685464e-10, 
    1.685195e-10, 1.685643e-10, 1.686042e-10, 1.686549e-10, 1.687479e-10, 
    1.687265e-10, 1.688048e-10, 1.680121e-10, 1.680588e-10, 1.680552e-10, 
    1.681044e-10, 1.681408e-10, 1.682203e-10, 1.683477e-10, 1.682999e-10, 
    1.683882e-10, 1.684058e-10, 1.682719e-10, 1.683536e-10, 1.680904e-10, 
    1.681323e-10, 1.681077e-10, 1.680155e-10, 1.683102e-10, 1.681584e-10, 
    1.684397e-10, 1.683572e-10, 1.685985e-10, 1.684778e-10, 1.687146e-10, 
    1.68815e-10, 1.689119e-10, 1.690228e-10, 1.680848e-10, 1.68053e-10, 
    1.681104e-10, 1.681891e-10, 1.682636e-10, 1.683621e-10, 1.683725e-10, 
    1.683908e-10, 1.68439e-10, 1.684793e-10, 1.683962e-10, 1.684894e-10, 
    1.681411e-10, 1.683236e-10, 1.680406e-10, 1.681249e-10, 1.681846e-10, 
    1.681589e-10, 1.682945e-10, 1.683264e-10, 1.68456e-10, 1.683892e-10, 
    1.687897e-10, 1.68612e-10, 1.69109e-10, 1.689693e-10, 1.680418e-10, 
    1.680849e-10, 1.682348e-10, 1.681635e-10, 1.68369e-10, 1.684195e-10, 
    1.68461e-10, 1.685134e-10, 1.685194e-10, 1.685505e-10, 1.684995e-10, 
    1.685487e-10, 1.683623e-10, 1.684456e-10, 1.682182e-10, 1.682731e-10, 
    1.68248e-10, 1.682201e-10, 1.683062e-10, 1.683974e-10, 1.684001e-10, 
    1.684292e-10, 1.685101e-10, 1.683698e-10, 1.688113e-10, 1.685368e-10, 
    1.68132e-10, 1.682143e-10, 1.68227e-10, 1.681949e-10, 1.684144e-10, 
    1.683346e-10, 1.685499e-10, 1.684918e-10, 1.685872e-10, 1.685397e-10, 
    1.685327e-10, 1.684719e-10, 1.684339e-10, 1.683381e-10, 1.682606e-10, 
    1.681996e-10, 1.682139e-10, 1.682809e-10, 1.684031e-10, 1.685196e-10, 
    1.68494e-10, 1.6858e-10, 1.68354e-10, 1.684482e-10, 1.684115e-10, 
    1.685074e-10, 1.682984e-10, 1.68474e-10, 1.682534e-10, 1.682729e-10, 
    1.683331e-10, 1.684541e-10, 1.684821e-10, 1.685106e-10, 1.684931e-10, 
    1.684064e-10, 1.683925e-10, 1.683318e-10, 1.683146e-10, 1.682687e-10, 
    1.682303e-10, 1.682652e-10, 1.683017e-10, 1.684067e-10, 1.685012e-10, 
    1.686047e-10, 1.686303e-10, 1.687498e-10, 1.686515e-10, 1.688127e-10, 
    1.68674e-10, 1.689152e-10, 1.684853e-10, 1.686715e-10, 1.683361e-10, 
    1.683722e-10, 1.68437e-10, 1.685874e-10, 1.68507e-10, 1.686015e-10, 
    1.68392e-10, 1.682828e-10, 1.682556e-10, 1.682032e-10, 1.682568e-10, 
    1.682524e-10, 1.683037e-10, 1.682873e-10, 1.684102e-10, 1.683442e-10, 
    1.685323e-10, 1.686009e-10, 1.687963e-10, 1.689161e-10, 1.690395e-10, 
    1.690937e-10, 1.691103e-10, 1.691172e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  1.093018, 1.074178, 1.077842, 1.062635, 1.071073, 1.061113, 1.0892, 
    1.073429, 1.083498, 1.091323, 1.03309, 1.061957, 1.003061, 1.021505, 
    0.975141, 1.005932, 0.9689265, 0.9760309, 0.9546425, 0.9607723, 
    0.9333884, 0.9518127, 0.9191797, 0.9377904, 0.9348798, 0.9524201, 
    1.056152, 1.036686, 1.057304, 1.05453, 1.055775, 1.070898, 1.078514, 
    1.094457, 1.091564, 1.079854, 1.053282, 1.062307, 1.039556, 1.04007, 
    1.01471, 1.026148, 0.9834754, 0.9956135, 0.9605165, 0.969349, 0.9609313, 
    0.9634842, 0.960898, 0.9738503, 0.9683019, 0.9796957, 1.024006, 1.010994, 
    1.049777, 1.073059, 1.088508, 1.099463, 1.097915, 1.094963, 1.079786, 
    1.065505, 1.054615, 1.047327, 1.040144, 1.018381, 1.006855, 0.9810195, 
    0.9856853, 0.9777809, 0.9702275, 0.9575384, 0.9596277, 0.9540351, 
    0.97799, 0.9620725, 0.9883422, 0.9811608, 1.038188, 1.059873, 1.06908, 
    1.077138, 1.096725, 1.0832, 1.088533, 1.075844, 1.067778, 1.071768, 
    1.047128, 1.056711, 1.006171, 1.027957, 0.9711086, 0.9847278, 0.9678429, 
    0.9764609, 0.961692, 0.9749844, 0.9519535, 0.9469347, 0.9503645, 
    0.9371872, 0.9757209, 0.9609311, 1.07188, 1.071229, 1.068197, 1.08152, 
    1.082335, 1.094536, 1.08368, 1.079055, 1.06731, 1.060359, 1.053749, 
    1.039208, 1.022955, 1.000205, 0.9838453, 0.9728705, 0.979601, 0.973659, 
    0.9803013, 0.9834138, 0.9488152, 0.96825, 0.939083, 0.9406982, 0.9539019, 
    0.9405162, 1.070772, 1.074516, 1.087511, 1.077342, 1.095865, 1.085499, 
    1.079535, 1.05651, 1.051448, 1.046752, 1.037476, 1.025563, 1.004648, 
    0.9864321, 0.969788, 0.9710081, 0.9705786, 0.9668583, 0.976072, 
    0.9653453, 0.9635441, 0.9682527, 0.9409145, 0.9487287, 0.9407325, 
    0.9458209, 1.073299, 1.066998, 1.070403, 1.063999, 1.068511, 1.04844, 
    1.042419, 1.014218, 1.025797, 1.007367, 1.023926, 1.020993, 1.006764, 
    1.023032, 0.9874365, 1.011575, 0.9667136, 0.9908442, 0.9652004, 
    0.9698601, 0.9621449, 0.9552323, 0.9465329, 0.9304704, 0.9341912, 
    0.9207514, 1.0576, 1.04942, 1.050141, 1.041577, 1.03524, 1.021501, 
    0.999443, 1.007741, 0.9925053, 0.9894452, 1.012591, 0.9983824, 1.043943, 
    1.036589, 1.040968, 1.056955, 1.005828, 1.032083, 0.9835747, 0.9978184, 
    0.9562179, 0.9769176, 0.936239, 0.9188224, 0.9024196, 0.8832309, 
    1.044954, 1.050514, 1.040558, 1.026774, 1.013977, 0.9969497, 0.9952071, 
    0.9920152, 0.9837456, 0.9767891, 0.9910054, 0.975045, 1.034882, 1.003548, 
    1.052616, 1.037853, 1.027587, 1.032091, 1.008689, 1.003169, 0.980722, 
    0.9923294, 0.9231219, 0.9537711, 0.8686102, 0.8924448, 1.052456, 
    1.044973, 1.018907, 1.031314, 0.9958128, 0.9870642, 0.9799495, 0.9708499, 
    0.9698676, 0.9644739, 0.9733116, 0.9648232, 0.9969135, 0.9825801, 
    1.021889, 1.012328, 1.016727, 1.021551, 1.00666, 0.9907815, 0.990443, 
    0.9853486, 0.9709836, 0.9956689, 0.9191611, 0.9664444, 1.036811, 
    1.022382, 1.020321, 1.025912, 0.9879414, 1.001708, 0.9646055, 0.9746404, 
    0.958196, 0.9663692, 0.9675713, 0.9780632, 0.9845921, 1.001077, 1.014479, 
    1.025101, 1.022632, 1.010962, 0.98981, 0.9697782, 0.974168, 0.9594462, 
    0.9983891, 0.9820692, 0.9883783, 0.9719229, 1.007961, 0.9772744, 
    1.015797, 1.012422, 1.001981, 0.9809611, 0.9763086, 0.9713381, 0.9744055, 
    0.989273, 0.9917079, 1.002235, 1.00514, 1.013157, 1.019791, 1.01373, 
    1.007362, 0.989267, 0.9729448, 0.9551337, 0.9507729, 0.9299354, 
    0.9468985, 0.9188973, 0.9427042, 0.9014761, 0.9754959, 0.9434056, 
    1.001506, 0.9952556, 0.9839441, 0.9579758, 0.9720004, 0.9555982, 
    0.9918033, 1.010559, 1.01541, 1.024456, 1.015203, 1.015956, 1.007099, 
    1.009945, 0.9886659, 1.000099, 0.9676012, 0.955728, 0.92216, 0.9015535, 
    0.8805574, 0.8712807, 0.8684563, 0.8672755,
  0.4710495, 0.455137, 0.4582155, 0.4454927, 0.4525349, 0.4442267, 0.4678084, 
    0.4545087, 0.4629835, 0.46961, 0.4211769, 0.4449283, 0.3970329, 
    0.4117954, 0.3751112, 0.3993157, 0.3703032, 0.3758026, 0.3593521, 
    0.3640348, 0.343316, 0.3571991, 0.3327746, 0.3466118, 0.3444313, 
    0.3576607, 0.4401114, 0.424107, 0.4410661, 0.4387688, 0.4397994, 
    0.4523885, 0.4587802, 0.4722748, 0.4698149, 0.459909, 0.4377372, 
    0.4452199, 0.4264545, 0.426875, 0.4063315, 0.4155467, 0.3816013, 
    0.3911356, 0.3638389, 0.3706299, 0.3641565, 0.3661148, 0.364131, 
    0.3741112, 0.3698219, 0.3786526, 0.4138146, 0.4033556, 0.4348452, 
    0.454197, 0.4672219, 0.4765425, 0.4752209, 0.4727047, 0.4598512, 
    0.4478837, 0.4388403, 0.4328286, 0.4269354, 0.4092784, 0.400051, 
    0.3796838, 0.38333, 0.377162, 0.3713083, 0.361561, 0.3631584, 0.3588892, 
    0.3773252, 0.3650309, 0.3854126, 0.3797945, 0.4253332, 0.4431969, 
    0.4508666, 0.4576229, 0.4742055, 0.4627312, 0.4672424, 0.4565367, 
    0.4497797, 0.4531173, 0.4326646, 0.4405748, 0.3995066, 0.4170107, 
    0.3719892, 0.3825806, 0.3694682, 0.3761368, 0.3647393, 0.3749907, 
    0.3573059, 0.3535002, 0.356099, 0.34616, 0.3755622, 0.3641561, 0.4532107, 
    0.4526657, 0.4501303, 0.4613133, 0.4620009, 0.472342, 0.463137, 
    0.4592363, 0.4493895, 0.4436007, 0.4381236, 0.4261696, 0.4129646, 
    0.394767, 0.3818905, 0.3733525, 0.3785792, 0.3739632, 0.3791246, 
    0.3815536, 0.3549239, 0.3697818, 0.3475825, 0.3487964, 0.3587877, 
    0.3486596, 0.4522832, 0.4554217, 0.4663767, 0.4577955, 0.4734731, 
    0.4646737, 0.4596403, 0.4404078, 0.4362237, 0.4323555, 0.4247545, 
    0.4150731, 0.3982946, 0.3839145, 0.3709691, 0.3719117, 0.3715797, 
    0.3687094, 0.3758347, 0.3675449, 0.3661604, 0.3697841, 0.3489591, 
    0.3548589, 0.3488223, 0.3526586, 0.4544007, 0.4491289, 0.4519747, 
    0.4466284, 0.4503921, 0.4337436, 0.4287971, 0.4059364, 0.4152626, 
    0.4004593, 0.41375, 0.4113826, 0.3999778, 0.4130279, 0.3847011, 
    0.4038194, 0.3685981, 0.3873762, 0.3674335, 0.3710247, 0.365087, 
    0.3598013, 0.3531967, 0.3411402, 0.3439169, 0.333934, 0.4413117, 
    0.4345505, 0.4351453, 0.4281081, 0.422931, 0.4117924, 0.3941636, 
    0.4007583, 0.388685, 0.3862783, 0.4046337, 0.3933237, 0.4300479, 
    0.4240299, 0.4276099, 0.4407764, 0.3992336, 0.42036, 0.3816789, 
    0.3928778, 0.3605529, 0.3764908, 0.3454492, 0.3325107, 0.3205261, 
    0.3067524, 0.4308778, 0.4354534, 0.4272743, 0.4160521, 0.4057435, 
    0.392191, 0.3908149, 0.388299, 0.3818128, 0.3763918, 0.3875039, 
    0.3750378, 0.4226368, 0.3974199, 0.4371869, 0.4250612, 0.4167109, 
    0.4203673, 0.401515, 0.3971196, 0.3794519, 0.3885465, 0.3356843, 
    0.3586875, 0.2964422, 0.3133321, 0.437056, 0.430894, 0.4097027, 
    0.4197356, 0.3912931, 0.3844101, 0.3788507, 0.3717889, 0.3710304, 
    0.3668748, 0.3736941, 0.3671436, 0.3921623, 0.3809021, 0.4121057, 
    0.4044234, 0.407951, 0.4118332, 0.3998968, 0.3873277, 0.3870624, 
    0.3830661, 0.3718895, 0.3911795, 0.3327586, 0.3683881, 0.4242118, 
    0.4125021, 0.4108415, 0.4153557, 0.3850979, 0.3959593, 0.3669761, 
    0.374724, 0.3620635, 0.3683329, 0.3692588, 0.3773822, 0.3824745, 
    0.3954584, 0.4061465, 0.4147, 0.4127052, 0.4033304, 0.3865643, 0.370961, 
    0.3743571, 0.3630196, 0.3933295, 0.3805029, 0.3854402, 0.372619, 
    0.4009338, 0.3767662, 0.4072036, 0.4044989, 0.396176, 0.3796379, 
    0.3760185, 0.3721664, 0.3745418, 0.3861426, 0.388057, 0.3963779, 
    0.3986866, 0.4050873, 0.4104152, 0.4055458, 0.4004558, 0.3861383, 
    0.3734096, 0.359726, 0.3564093, 0.3407404, 0.3534718, 0.332564, 
    0.3503032, 0.3198406, 0.375386, 0.3508336, 0.3957994, 0.3908533, 
    0.381967, 0.3618942, 0.3726789, 0.3600795, 0.3881322, 0.4030077, 
    0.4068934, 0.4141778, 0.4067274, 0.4073315, 0.4002466, 0.4025182, 
    0.3856664, 0.3946838, 0.3692817, 0.3601787, 0.3349741, 0.3198979, 
    0.3048561, 0.2983138, 0.2963348, 0.2955092,
  0.2132781, 0.2051227, 0.2066971, 0.2002013, 0.2037933, 0.1995565, 
    0.2116135, 0.2048016, 0.2091388, 0.2125385, 0.1878664, 0.1999138, 
    0.175726, 0.1831363, 0.1647988, 0.1768692, 0.1624146, 0.1651421, 
    0.1570015, 0.1593132, 0.1491191, 0.1559402, 0.1439669, 0.1507348, 
    0.1496656, 0.1561676, 0.1974624, 0.1893471, 0.1979479, 0.1967798, 
    0.1973038, 0.2037185, 0.206986, 0.2139079, 0.2126438, 0.2075638, 
    0.1962556, 0.2000624, 0.1905347, 0.1907475, 0.1803888, 0.1850258, 
    0.1680244, 0.1727774, 0.1592164, 0.1625765, 0.1593734, 0.1603415, 
    0.1593608, 0.1643026, 0.1621763, 0.1665579, 0.184153, 0.1788948, 
    0.194787, 0.2046423, 0.2113124, 0.2161034, 0.2154231, 0.2141289, 
    0.2075343, 0.2014199, 0.1968162, 0.1937639, 0.1907781, 0.1818698, 
    0.1772376, 0.1670705, 0.1688849, 0.1658172, 0.1629127, 0.1580914, 
    0.1588802, 0.1567732, 0.1658983, 0.1598055, 0.1699223, 0.1671257, 
    0.1899672, 0.1990322, 0.2029415, 0.2063939, 0.2149007, 0.2090094, 
    0.211323, 0.2058384, 0.2023869, 0.2040908, 0.1936807, 0.1976981, 
    0.1769648, 0.1857639, 0.1632502, 0.1685118, 0.1620011, 0.1653081, 
    0.1596614, 0.1647391, 0.1559928, 0.1541189, 0.1553982, 0.1505132, 
    0.1650227, 0.1593731, 0.2041385, 0.2038601, 0.2025658, 0.208283, 
    0.2086352, 0.2139424, 0.2092174, 0.2072195, 0.2021879, 0.1992378, 
    0.1964519, 0.1903905, 0.1837249, 0.1745923, 0.1681683, 0.1639262, 
    0.1665214, 0.1642292, 0.1667925, 0.1680007, 0.1548196, 0.1621563, 
    0.1512111, 0.151807, 0.1567232, 0.1517398, 0.2036648, 0.2052683, 
    0.2108787, 0.2064822, 0.214524, 0.2100052, 0.2074263, 0.1976131, 
    0.1954869, 0.1935239, 0.1896747, 0.1847871, 0.1763577, 0.169176, 
    0.1627446, 0.1632118, 0.1630472, 0.1616254, 0.165158, 0.161049, 0.160364, 
    0.1621575, 0.1518869, 0.1547876, 0.1518197, 0.1537049, 0.2047465, 
    0.2020549, 0.2035073, 0.20078, 0.2026994, 0.194228, 0.1917205, 0.1801903, 
    0.1848826, 0.1774423, 0.1841204, 0.1829285, 0.1772009, 0.1837568, 
    0.1695677, 0.1791275, 0.1615702, 0.1709011, 0.1609938, 0.1627721, 
    0.1598333, 0.1572231, 0.1539696, 0.1480537, 0.1494135, 0.1445325, 
    0.1980729, 0.1946375, 0.1949394, 0.1913717, 0.1887527, 0.1831347, 
    0.1742906, 0.1775922, 0.1715541, 0.1703538, 0.1795362, 0.1738707, 
    0.1923542, 0.1893082, 0.1911194, 0.1978006, 0.1768281, 0.187454, 
    0.168063, 0.1736478, 0.1575939, 0.1654838, 0.1501646, 0.1438382, 
    0.1380105, 0.1313518, 0.1927748, 0.1950958, 0.1909496, 0.1852805, 
    0.1800935, 0.1733046, 0.1726173, 0.1713615, 0.1681297, 0.1654347, 
    0.1709648, 0.1647624, 0.188604, 0.1759198, 0.1959761, 0.1898297, 
    0.1856127, 0.1874577, 0.1779716, 0.1757695, 0.1669552, 0.171485, 
    0.1453867, 0.1566737, 0.1263956, 0.1345273, 0.1959096, 0.192783, 
    0.1820833, 0.1871388, 0.1728561, 0.1694228, 0.1666564, 0.1631509, 
    0.162775, 0.1607174, 0.1640957, 0.1608504, 0.1732903, 0.1676766, 
    0.1832925, 0.1794307, 0.1812026, 0.1831553, 0.1771604, 0.170877, 
    0.1707447, 0.1687535, 0.1632006, 0.1727993, 0.143959, 0.1614661, 
    0.1894002, 0.1834919, 0.1826562, 0.1849295, 0.1697655, 0.1751887, 
    0.1607675, 0.1646067, 0.1583395, 0.1614389, 0.1618974, 0.1659266, 
    0.168459, 0.1749381, 0.1802959, 0.1845991, 0.1835943, 0.1788822, 
    0.1704963, 0.1627406, 0.1644246, 0.1588117, 0.1738736, 0.1674779, 
    0.169936, 0.1635624, 0.1776802, 0.1656205, 0.180827, 0.1794686, 
    0.1752972, 0.1670477, 0.1652493, 0.163338, 0.1645163, 0.1702861, 
    0.1712407, 0.1753982, 0.1765541, 0.179764, 0.1824417, 0.1799942, 
    0.1774406, 0.170284, 0.1639545, 0.1571859, 0.155551, 0.147858, 0.1541049, 
    0.1438641, 0.1525469, 0.137678, 0.1649352, 0.1528076, 0.1751088, 
    0.1726364, 0.1682064, 0.1582559, 0.1635921, 0.1573603, 0.1712783, 
    0.1787202, 0.1806711, 0.1843359, 0.1805877, 0.1808913, 0.1773357, 
    0.1784747, 0.1700488, 0.1745507, 0.1619087, 0.1574093, 0.14504, 
    0.1377058, 0.1304384, 0.1272935, 0.1263441, 0.1259483,
  0.05204878, 0.04963026, 0.0500953, 0.04818233, 0.04923828, 0.04799328, 
    0.05155321, 0.04953552, 0.05081828, 0.05182849, 0.04459244, 0.04809802, 
    0.0411155, 0.043231, 0.03803579, 0.04144046, 0.03737032, 0.0381318, 
    0.03586819, 0.03650819, 0.03370298, 0.0355751, 0.0323023, 0.03414462, 
    0.03385223, 0.03563787, 0.04738035, 0.04502038, 0.04752232, 0.04718091, 
    0.04733398, 0.04921624, 0.05018074, 0.05223652, 0.05185982, 0.05035171, 
    0.04702786, 0.04814159, 0.04536419, 0.04542585, 0.04244415, 0.04377382, 
    0.03893982, 0.04027974, 0.03648135, 0.03741544, 0.03652487, 0.03679358, 
    0.03652138, 0.03789709, 0.03730392, 0.03852829, 0.04352291, 0.04201751, 
    0.04659963, 0.04948852, 0.0514637, 0.05289211, 0.05268881, 0.05230245, 
    0.05034295, 0.04854005, 0.04719154, 0.04630176, 0.04543472, 0.04286793, 
    0.0415453, 0.03867203, 0.03918172, 0.03832075, 0.03750915, 0.03616965, 
    0.03638814, 0.03580511, 0.03834346, 0.03664477, 0.03947377, 0.0386875, 
    0.04519984, 0.04783968, 0.04898744, 0.05000569, 0.05253279, 0.05077992, 
    0.05146682, 0.04984154, 0.04882429, 0.04932592, 0.04627756, 0.04744924, 
    0.04146768, 0.04398623, 0.03760328, 0.0390768, 0.03725514, 0.03817824, 
    0.03660478, 0.03801909, 0.03558962, 0.03507328, 0.03542562, 0.03408398, 
    0.03809841, 0.03652481, 0.04933998, 0.04925795, 0.0488769, 0.05056464, 
    0.05066901, 0.05224683, 0.0508416, 0.05024981, 0.04876576, 0.04789989, 
    0.04708517, 0.04532242, 0.04339995, 0.04079375, 0.03898025, 0.03779197, 
    0.03851805, 0.03787659, 0.03859407, 0.03893315, 0.03526617, 0.03729837, 
    0.03427503, 0.03443832, 0.03579128, 0.0344199, 0.04920041, 0.04967322, 
    0.05133478, 0.05003178, 0.05242034, 0.05107534, 0.050311, 0.0474244, 
    0.04680361, 0.04623196, 0.04511517, 0.04370517, 0.04129502, 0.03926362, 
    0.03746228, 0.03759256, 0.03754666, 0.03715054, 0.03813626, 0.0369902, 
    0.03679984, 0.0372987, 0.03446022, 0.03525736, 0.0344418, 0.03495942, 
    0.04951926, 0.04872666, 0.04915402, 0.04835214, 0.04891621, 0.04643682, 
    0.04570804, 0.04238742, 0.04373263, 0.04160357, 0.04351356, 0.04317139, 
    0.04153485, 0.04340911, 0.03937389, 0.0420839, 0.0371352, 0.0397497, 
    0.03697488, 0.03746996, 0.03665248, 0.03592942, 0.03503222, 0.03341239, 
    0.03378338, 0.03245548, 0.04755887, 0.04655606, 0.04664401, 0.04560684, 
    0.0448485, 0.04323056, 0.0407082, 0.04164626, 0.03993401, 0.03959535, 
    0.04220059, 0.04058921, 0.04589199, 0.04500913, 0.04553369, 0.04747922, 
    0.04142877, 0.04447339, 0.03895067, 0.04052609, 0.03603197, 0.03822741, 
    0.03398864, 0.03226746, 0.03069767, 0.028923, 0.04601418, 0.04668959, 
    0.04548445, 0.0438471, 0.04235975, 0.04042891, 0.04023444, 0.03987962, 
    0.0389694, 0.03821366, 0.03976768, 0.03802561, 0.0448055, 0.04117056, 
    0.04694629, 0.04516004, 0.0439427, 0.04447447, 0.04175431, 0.04112785, 
    0.0386397, 0.03991449, 0.0326871, 0.03577762, 0.02761557, 0.02976679, 
    0.04692689, 0.04601657, 0.04292909, 0.04438246, 0.04030199, 0.03933309, 
    0.03855588, 0.03757559, 0.03747075, 0.03689804, 0.03783929, 0.03693499, 
    0.04042485, 0.03884212, 0.04327582, 0.04217045, 0.04267691, 0.04323646, 
    0.04152334, 0.03974289, 0.03970559, 0.03914475, 0.03758944, 0.04028593, 
    0.03230014, 0.03710623, 0.04503575, 0.04333307, 0.04309331, 0.04374613, 
    0.03942959, 0.04096296, 0.03691196, 0.03798208, 0.03623835, 0.03709867, 
    0.03722626, 0.03835139, 0.03906195, 0.04089185, 0.0424176, 0.04365112, 
    0.04336246, 0.04201391, 0.03963554, 0.03746117, 0.03793119, 0.03636914, 
    0.04059004, 0.03878636, 0.03947763, 0.0376904, 0.0416713, 0.03826566, 
    0.04256945, 0.04218126, 0.04099375, 0.03866562, 0.03816179, 0.03762778, 
    0.03795681, 0.03957628, 0.03984554, 0.04102243, 0.04135085, 0.04226562, 
    0.04303181, 0.04233139, 0.04160307, 0.03957568, 0.03779987, 0.03591916, 
    0.03546777, 0.03335906, 0.03506942, 0.03227446, 0.03464128, 0.03060855, 
    0.03807392, 0.03471285, 0.04094027, 0.04023986, 0.03899094, 0.03621517, 
    0.0376987, 0.03596736, 0.03985613, 0.04196771, 0.04252487, 0.04357549, 
    0.04250103, 0.04258784, 0.04157323, 0.04189771, 0.0395094, 0.04078197, 
    0.03722941, 0.0359809, 0.03259306, 0.03061602, 0.02868119, 0.02785156, 
    0.02760206, 0.02749815,
  0.004543171, 0.00427812, 0.004328803, 0.004121187, 0.004235503, 
    0.004100795, 0.004488567, 0.00426781, 0.004407865, 0.004518881, 
    0.003737931, 0.00411209, 0.003374959, 0.003594819, 0.003060545, 
    0.003408529, 0.002993513, 0.003070243, 0.002843425, 0.002907164, 
    0.002630129, 0.002814341, 0.002494121, 0.002673338, 0.002644715, 
    0.002820564, 0.00403484, 0.003783173, 0.004050096, 0.004013431, 
    0.00402986, 0.004233111, 0.004338129, 0.004563898, 0.004522334, 
    0.004356805, 0.003997019, 0.00411679, 0.003819609, 0.003826152, 
    0.003512682, 0.003651729, 0.003152128, 0.003288961, 0.002904484, 
    0.002998048, 0.002908829, 0.002935686, 0.00290848, 0.003046547, 
    0.002986843, 0.003110363, 0.003625399, 0.003468324, 0.003951181, 
    0.004262698, 0.00447872, 0.00463644, 0.004613916, 0.004571181, 
    0.004355848, 0.004159835, 0.004014571, 0.003919366, 0.003827093, 
    0.003556867, 0.003419376, 0.003124937, 0.003176735, 0.003089348, 
    0.00300747, 0.002873409, 0.002895184, 0.002837159, 0.003091646, 
    0.002920806, 0.003206501, 0.003126506, 0.003802182, 0.004084244, 
    0.004208284, 0.004319025, 0.004596648, 0.004403663, 0.004479064, 
    0.004301129, 0.004190601, 0.004245024, 0.003916785, 0.004042241, 
    0.003411344, 0.003674053, 0.003016941, 0.003166057, 0.002981945, 
    0.003074935, 0.00291681, 0.003058858, 0.00281578, 0.002764696, 
    0.002799532, 0.002667397, 0.003066869, 0.002908823, 0.004246552, 
    0.00423764, 0.004196302, 0.004380091, 0.004391515, 0.004565036, 
    0.004410421, 0.004345672, 0.004184261, 0.00409073, 0.004003163, 
    0.003815178, 0.003612511, 0.003341793, 0.003156238, 0.003035947, 
    0.003109326, 0.003044478, 0.00311703, 0.00315145, 0.002783755, 
    0.002986286, 0.002686126, 0.002702159, 0.002835787, 0.002700349, 
    0.004231391, 0.004282795, 0.004464547, 0.004321872, 0.004584211, 
    0.004436055, 0.004352356, 0.004039572, 0.003973, 0.00391192, 0.00379321, 
    0.003644521, 0.003393495, 0.003185076, 0.003002757, 0.003015863, 
    0.003011244, 0.002971448, 0.003070693, 0.002955372, 0.002936312, 
    0.002986319, 0.00270431, 0.002782884, 0.0027025, 0.002753458, 
    0.004266042, 0.004180028, 0.004226356, 0.004139523, 0.004200561, 
    0.003933785, 0.003856128, 0.003506776, 0.003647404, 0.003425407, 
    0.003624419, 0.003588582, 0.003418294, 0.00361347, 0.003196314, 
    0.003475219, 0.002969909, 0.003234679, 0.002953837, 0.003003529, 
    0.002921576, 0.00284951, 0.002760641, 0.002601784, 0.002637985, 
    0.002508919, 0.004054025, 0.003946524, 0.003955926, 0.003845371, 
    0.003764988, 0.003594773, 0.003332988, 0.003429827, 0.003253531, 
    0.00321891, 0.003487343, 0.003320748, 0.003875696, 0.003781982, 
    0.003837601, 0.004045463, 0.00340732, 0.003725368, 0.00315323, 
    0.003314259, 0.002859707, 0.003079907, 0.00265806, 0.002490758, 
    0.002340276, 0.002172651, 0.003888706, 0.0039608, 0.003832372, 
    0.003659427, 0.003503897, 0.003304274, 0.003284314, 0.003247966, 
    0.003155134, 0.003078517, 0.003236517, 0.003059517, 0.003760441, 
    0.003380641, 0.003988279, 0.003797964, 0.003669476, 0.003725481, 
    0.003441022, 0.003376234, 0.003121658, 0.003251534, 0.002531328, 
    0.00283443, 0.00205091, 0.002252014, 0.0039862, 0.003888961, 0.003563254, 
    0.003715777, 0.003291244, 0.003192155, 0.00311316, 0.003014154, 
    0.003003609, 0.002946141, 0.003040718, 0.002949842, 0.003303858, 
    0.003142201, 0.003599511, 0.00348421, 0.003536935, 0.00359539, 
    0.003417103, 0.003233983, 0.003230171, 0.003172972, 0.003015548, 
    0.003289597, 0.002493912, 0.002967003, 0.0037848, 0.003605505, 
    0.003580415, 0.003648821, 0.003201994, 0.003359227, 0.002947535, 
    0.003055122, 0.002880252, 0.002966245, 0.002979046, 0.003092449, 
    0.003164546, 0.003351897, 0.003509918, 0.003638847, 0.003608583, 
    0.00346795, 0.003223014, 0.003002645, 0.003049986, 0.00289329, 
    0.003320833, 0.003136539, 0.003206894, 0.003025714, 0.003432421, 
    0.003083775, 0.003525733, 0.003485335, 0.003362401, 0.003124287, 
    0.003073273, 0.003019408, 0.003052572, 0.003216962, 0.00324448, 
    0.003365358, 0.003399264, 0.003494105, 0.003573986, 0.003500946, 
    0.003425356, 0.003216901, 0.003036743, 0.00284849, 0.002803706, 
    0.002596589, 0.002764314, 0.002491433, 0.002722113, 0.002331794, 
    0.003064395, 0.002729158, 0.003356888, 0.00328487, 0.003157325, 
    0.002877943, 0.003026549, 0.002853282, 0.003245563, 0.003463154, 
    0.003521088, 0.003630912, 0.003518605, 0.003527649, 0.003422267, 
    0.003455892, 0.003210136, 0.00334058, 0.002979362, 0.002854628, 
    0.002522224, 0.002332505, 0.002150021, 0.002072772, 0.00204966, 
    0.002040051,
  0.0001251994, 0.0001159854, 0.0001177354, 0.0001106029, 0.0001145183, 
    0.0001099076, 0.0001232887, 0.0001156301, 0.0001204767, 0.0001243486, 
    9.769691e-05, 0.0001102927, 8.580387e-05, 9.29681e-05, 7.578008e-05, 
    8.68897e-05, 7.367827e-05, 7.608521e-05, 6.901897e-05, 7.098968e-05, 
    6.25126e-05, 6.81237e-05, 5.843752e-05, 6.381943e-05, 6.295308e-05, 
    6.831506e-05, 0.0001076652, 9.920227e-05, 0.000108183, 0.0001069395, 
    0.0001074963, 0.000114436, 0.0001180581, 0.0001259263, 0.0001244695, 
    0.0001187048, 0.0001063839, 0.000110453, 0.0001004182, 0.0001006369, 
    9.027719e-05, 9.484249e-05, 7.867203e-05, 8.303572e-05, 7.090659e-05, 
    7.382006e-05, 7.104132e-05, 7.187538e-05, 7.10305e-05, 7.534013e-05, 
    7.346983e-05, 7.735032e-05, 9.397427e-05, 8.883108e-05, 0.0001048354, 
    0.000115454, 0.0001229449, 0.0001284775, 0.0001276842, 0.0001261819, 
    0.0001186716, 0.0001119233, 0.0001069781, 0.0001037636, 0.0001006684, 
    9.172262e-05, 8.724119e-05, 7.781101e-05, 7.945303e-05, 7.668711e-05, 
    7.411486e-05, 6.994454e-05, 7.061836e-05, 6.882589e-05, 7.675956e-05, 
    7.141302e-05, 8.039994e-05, 7.786063e-05, 9.983624e-05, 0.000109344, 
    0.0001135834, 0.0001173974, 0.0001270767, 0.0001203306, 0.0001229569, 
    0.0001167792, 0.0001129769, 0.0001148457, 0.0001036767, 0.0001079164, 
    8.698091e-05, 9.557995e-05, 7.441143e-05, 7.911392e-05, 7.331685e-05, 
    7.623295e-05, 7.128895e-05, 7.572705e-05, 6.816793e-05, 6.660136e-05, 
    6.766883e-05, 6.363939e-05, 7.597905e-05, 7.104112e-05, 0.0001148982, 
    0.0001145917, 0.0001131723, 0.0001195121, 0.0001199087, 0.0001259662, 
    0.0001205655, 0.0001183192, 0.0001127596, 0.0001095648, 0.0001065918, 
    0.0001002702, 9.354993e-05, 8.473398e-05, 7.880237e-05, 7.500733e-05, 
    7.731757e-05, 7.527516e-05, 7.7561e-05, 7.865056e-05, 6.718493e-05, 
    7.345243e-05, 6.42073e-05, 6.469429e-05, 6.878361e-05, 6.463927e-05, 
    0.0001143769, 0.0001161466, 0.0001224503, 0.0001174958, 0.0001266396, 
    0.0001214574, 0.0001185507, 0.0001078258, 0.0001055719, 0.000103513, 
    9.953689e-05, 9.460464e-05, 8.640307e-05, 7.971811e-05, 7.396737e-05, 
    7.437765e-05, 7.4233e-05, 7.298921e-05, 7.609939e-05, 7.248807e-05, 
    7.189486e-05, 7.345346e-05, 6.475971e-05, 6.715824e-05, 6.470467e-05, 
    6.625779e-05, 0.0001155692, 0.0001126146, 0.0001142039, 0.0001112289, 
    0.0001133184, 0.000104249, 0.0001016401, 9.008435e-05, 9.469975e-05, 
    8.743677e-05, 9.394198e-05, 9.276318e-05, 8.720613e-05, 9.35815e-05, 
    8.007561e-05, 8.905551e-05, 7.29412e-05, 8.129858e-05, 7.244026e-05, 
    7.399153e-05, 7.143693e-05, 6.92066e-05, 6.647737e-05, 6.165847e-05, 
    6.274974e-05, 5.887801e-05, 0.0001083165, 0.0001046784, 0.0001049955, 
    0.0001012799, 9.859656e-05, 9.296659e-05, 8.445042e-05, 8.758014e-05, 
    8.190099e-05, 8.079541e-05, 8.945049e-05, 8.40566e-05, 0.0001022962, 
    9.916256e-05, 0.0001010198, 0.0001080257, 8.685055e-05, 9.727974e-05, 
    7.870699e-05, 8.384799e-05, 6.952124e-05, 7.638954e-05, 6.335669e-05, 
    5.83375e-05, 5.390045e-05, 4.904858e-05, 0.0001027329, 0.00010516, 
    0.0001008449, 9.509665e-05, 8.999037e-05, 8.352719e-05, 8.28867e-05, 
    8.172305e-05, 7.876736e-05, 7.634576e-05, 8.135727e-05, 7.574777e-05, 
    9.844526e-05, 8.598745e-05, 0.0001060883, 9.969548e-05, 9.542866e-05, 
    9.72835e-05, 8.794352e-05, 8.584504e-05, 7.770728e-05, 8.183712e-05, 
    5.954645e-05, 6.874183e-05, 4.558753e-05, 5.133351e-05, 0.000106018, 
    0.0001027414, 9.193197e-05, 9.696157e-05, 8.310895e-05, 7.994327e-05, 
    7.743869e-05, 7.432413e-05, 7.399402e-05, 7.220062e-05, 7.515708e-05, 
    7.231584e-05, 8.351381e-05, 7.835747e-05, 9.312232e-05, 8.93484e-05, 
    9.106998e-05, 9.298688e-05, 8.71675e-05, 8.127636e-05, 8.115466e-05, 
    7.933348e-05, 7.43678e-05, 8.30561e-05, 5.843129e-05, 7.285056e-05, 
    9.925648e-05, 9.331945e-05, 9.249499e-05, 9.474652e-05, 8.02564e-05, 
    8.5296e-05, 7.224402e-05, 7.560958e-05, 7.015614e-05, 7.282694e-05, 
    7.322633e-05, 7.678488e-05, 7.906597e-05, 8.505963e-05, 9.018691e-05, 
    9.441753e-05, 9.342069e-05, 8.88189e-05, 8.092631e-05, 7.396386e-05, 
    7.544817e-05, 7.05597e-05, 8.405935e-05, 7.817813e-05, 8.041248e-05, 
    7.468636e-05, 8.766432e-05, 7.651141e-05, 9.070362e-05, 8.938504e-05, 
    8.539842e-05, 7.779044e-05, 7.618062e-05, 7.448871e-05, 7.552943e-05, 
    8.073331e-05, 8.161163e-05, 8.549387e-05, 8.658974e-05, 8.967093e-05, 
    9.228398e-05, 8.989409e-05, 8.743508e-05, 8.073137e-05, 7.503232e-05, 
    6.917513e-05, 6.779696e-05, 6.15022e-05, 6.658968e-05, 5.835757e-05, 
    6.530149e-05, 5.365259e-05, 7.59012e-05, 6.551618e-05, 8.522056e-05, 
    8.290451e-05, 7.883684e-05, 7.008472e-05, 7.471255e-05, 6.932294e-05, 
    8.164624e-05, 8.866286e-05, 9.05518e-05, 9.415594e-05, 9.047065e-05, 
    9.076625e-05, 8.733491e-05, 8.842666e-05, 8.051575e-05, 8.469492e-05, 
    7.32362e-05, 6.936448e-05, 5.92747e-05, 5.367335e-05, 4.840114e-05, 
    4.620507e-05, 4.555227e-05, 4.528147e-05,
  9.624799e-07, 8.692003e-07, 8.867518e-07, 8.157223e-07, 8.545479e-07, 
    8.088703e-07, 9.429625e-07, 8.656469e-07, 9.144015e-07, 9.537783e-07, 
    6.9074e-07, 8.126629e-07, 5.79961e-07, 6.461634e-07, 4.902151e-07, 
    5.898884e-07, 4.718508e-07, 4.928947e-07, 4.317359e-07, 4.486012e-07, 
    3.771623e-07, 4.241246e-07, 3.438939e-07, 3.879831e-07, 3.808015e-07, 
    4.257488e-07, 7.868621e-07, 7.050716e-07, 7.919318e-07, 7.797693e-07, 
    7.852102e-07, 8.537281e-07, 8.899964e-07, 9.699286e-07, 9.550135e-07, 
    8.965072e-07, 7.743489e-07, 8.142431e-07, 7.166963e-07, 7.187919e-07, 
    6.211052e-07, 6.637511e-07, 5.157465e-07, 5.548305e-07, 4.47887e-07, 
    4.730845e-07, 4.490452e-07, 4.562299e-07, 4.489521e-07, 4.863575e-07, 
    4.700386e-07, 5.040405e-07, 6.55591e-07, 6.077336e-07, 7.592872e-07, 
    8.638871e-07, 9.394593e-07, 9.961738e-07, 9.879959e-07, 9.725512e-07, 
    8.961733e-07, 8.287699e-07, 7.801463e-07, 7.48901e-07, 7.190935e-07, 
    6.345371e-07, 5.931102e-07, 5.081135e-07, 5.226928e-07, 4.981902e-07, 
    4.75652e-07, 4.396381e-07, 4.454119e-07, 4.300917e-07, 4.988286e-07, 
    4.522437e-07, 5.311435e-07, 5.085528e-07, 7.111273e-07, 8.033253e-07, 
    8.4524e-07, 8.833553e-07, 9.817437e-07, 9.129236e-07, 9.395816e-07, 
    8.771516e-07, 8.392141e-07, 8.578129e-07, 7.480608e-07, 7.893202e-07, 
    5.90724e-07, 6.707002e-07, 4.782381e-07, 5.196741e-07, 4.687095e-07, 
    4.941933e-07, 4.511754e-07, 4.897498e-07, 4.244999e-07, 4.112556e-07, 
    4.202697e-07, 3.864881e-07, 4.91962e-07, 4.490434e-07, 8.583373e-07, 
    8.552802e-07, 8.411549e-07, 9.04651e-07, 9.086565e-07, 9.703383e-07, 
    9.153009e-07, 8.926235e-07, 8.370579e-07, 8.054964e-07, 7.763762e-07, 
    7.152788e-07, 6.516112e-07, 5.702177e-07, 5.169042e-07, 4.834444e-07, 
    5.037512e-07, 4.857886e-07, 5.059023e-07, 5.155558e-07, 4.161778e-07, 
    4.698873e-07, 3.912087e-07, 3.952674e-07, 4.297318e-07, 3.948084e-07, 
    8.531393e-07, 8.708137e-07, 9.344261e-07, 8.843435e-07, 9.772506e-07, 
    9.243395e-07, 8.949547e-07, 7.884333e-07, 7.664421e-07, 7.464782e-07, 
    7.082664e-07, 6.615133e-07, 5.854344e-07, 5.250554e-07, 4.743671e-07, 
    4.779434e-07, 4.766818e-07, 4.658661e-07, 4.930192e-07, 4.615247e-07, 
    4.56398e-07, 4.698963e-07, 3.958134e-07, 4.159523e-07, 3.95354e-07, 
    4.083643e-07, 8.650379e-07, 8.356192e-07, 8.514155e-07, 8.219024e-07, 
    8.426063e-07, 7.536011e-07, 7.284219e-07, 6.193183e-07, 6.624079e-07, 
    5.949046e-07, 6.55288e-07, 6.442472e-07, 5.927886e-07, 6.519071e-07, 
    5.282456e-07, 6.098045e-07, 4.654497e-07, 5.391925e-07, 4.61111e-07, 
    4.745775e-07, 4.524497e-07, 4.333351e-07, 4.102116e-07, 3.701293e-07, 
    3.791206e-07, 3.474546e-07, 7.932398e-07, 7.577634e-07, 7.608408e-07, 
    7.249605e-07, 6.992969e-07, 6.461493e-07, 5.676417e-07, 5.962209e-07, 
    5.446037e-07, 5.346823e-07, 6.134529e-07, 5.640686e-07, 7.347353e-07, 
    7.046926e-07, 7.224639e-07, 7.903911e-07, 5.895298e-07, 6.867803e-07, 
    5.16057e-07, 5.621779e-07, 4.360199e-07, 4.955705e-07, 3.841433e-07, 
    3.430865e-07, 3.077373e-07, 2.701712e-07, 7.389445e-07, 7.624382e-07, 
    7.207859e-07, 6.661442e-07, 6.184478e-07, 5.592734e-07, 5.534849e-07, 
    5.43004e-07, 5.165933e-07, 4.951854e-07, 5.397191e-07, 4.899316e-07, 
    6.978561e-07, 5.816367e-07, 7.714679e-07, 7.097816e-07, 6.692732e-07, 
    6.86816e-07, 5.995599e-07, 5.803367e-07, 5.071958e-07, 5.440294e-07, 
    3.528746e-07, 4.293763e-07, 2.441161e-07, 2.877159e-07, 7.707834e-07, 
    7.390271e-07, 6.364879e-07, 6.837638e-07, 5.55492e-07, 5.270641e-07, 
    5.048212e-07, 4.774766e-07, 4.745992e-07, 4.590388e-07, 4.847547e-07, 
    4.600349e-07, 5.591525e-07, 5.129548e-07, 6.476063e-07, 6.125093e-07, 
    6.284641e-07, 6.46339e-07, 5.924344e-07, 5.389931e-07, 5.379014e-07, 
    5.216282e-07, 4.778575e-07, 5.550145e-07, 3.438435e-07, 4.64664e-07, 
    7.055889e-07, 6.494519e-07, 6.417412e-07, 6.628479e-07, 5.298605e-07, 
    5.753311e-07, 4.59414e-07, 4.887193e-07, 4.414493e-07, 4.644593e-07, 
    4.679235e-07, 4.990517e-07, 5.192475e-07, 5.731793e-07, 6.202685e-07, 
    6.59754e-07, 6.504002e-07, 6.076212e-07, 5.358547e-07, 4.743365e-07, 
    4.873042e-07, 4.449085e-07, 5.640935e-07, 5.113649e-07, 5.312556e-07, 
    4.806384e-07, 5.96994e-07, 4.966431e-07, 6.250611e-07, 6.128479e-07, 
    5.762641e-07, 5.079315e-07, 4.937332e-07, 4.789126e-07, 4.880165e-07, 
    5.341262e-07, 5.420029e-07, 5.77134e-07, 5.87142e-07, 6.154913e-07, 
    6.397713e-07, 6.175563e-07, 5.948891e-07, 5.341088e-07, 4.836629e-07, 
    4.330668e-07, 4.213547e-07, 3.688459e-07, 4.111573e-07, 3.432484e-07, 
    4.003417e-07, 3.0579e-07, 4.912783e-07, 4.021395e-07, 5.746441e-07, 
    5.536457e-07, 5.172105e-07, 4.408378e-07, 4.808672e-07, 4.343274e-07, 
    5.423139e-07, 6.061825e-07, 6.236519e-07, 6.572965e-07, 6.228991e-07, 
    6.256425e-07, 5.939699e-07, 6.040061e-07, 5.321792e-07, 5.698626e-07, 
    4.680092e-07, 4.346817e-07, 3.506687e-07, 3.05953e-07, 2.652489e-07, 
    2.487178e-07, 2.43854e-07, 2.418433e-07,
  1.162747e-09, 9.63801e-10, 1.000341e-09, 8.551568e-10, 9.336257e-10, 
    8.415381e-10, 1.120171e-09, 9.564554e-10, 1.058759e-09, 1.143705e-09, 
    6.183029e-10, 8.490674e-10, 4.309834e-10, 5.401683e-10, 2.974938e-10, 
    4.468073e-10, 2.724508e-10, 3.012158e-10, 2.206866e-10, 2.419447e-10, 
    1.572559e-10, 2.113404e-10, 1.229216e-10, 1.691538e-10, 1.612185e-10, 
    2.133217e-10, 7.982728e-10, 6.441664e-10, 8.081739e-10, 7.84487e-10, 
    7.950552e-10, 9.319466e-10, 1.007143e-09, 1.179124e-09, 1.146402e-09, 
    1.020834e-09, 7.740041e-10, 8.522108e-10, 6.65402e-10, 6.692543e-10, 
    4.978439e-10, 5.705703e-10, 3.33642e-10, 3.918339e-10, 2.410294e-10, 
    2.741074e-10, 2.425143e-10, 2.518035e-10, 2.42395e-10, 2.921656e-10, 
    2.700242e-10, 3.168798e-10, 5.563947e-10, 4.757486e-10, 7.451164e-10, 
    9.528244e-10, 1.112581e-09, 1.237381e-09, 1.219136e-09, 1.184907e-09, 
    1.02013e-09, 8.81282e-10, 7.852176e-10, 7.254057e-10, 6.698094e-10, 
    5.203842e-10, 4.519855e-10, 3.226763e-10, 3.437367e-10, 3.086216e-10, 
    2.77567e-10, 2.305538e-10, 2.378676e-10, 2.186544e-10, 3.095188e-10, 
    2.466334e-10, 3.56164e-10, 3.233036e-10, 6.552004e-10, 8.305681e-10, 
    9.146154e-10, 9.932366e-10, 1.205244e-09, 1.05561e-09, 1.112846e-09, 
    9.803016e-10, 9.023741e-10, 9.403236e-10, 7.238187e-10, 8.030684e-10, 
    4.481482e-10, 5.82737e-10, 2.81068e-10, 3.393363e-10, 2.682496e-10, 
    3.030257e-10, 2.452548e-10, 2.968492e-10, 2.117976e-10, 1.958976e-10, 
    2.066667e-10, 1.674894e-10, 2.999184e-10, 2.425121e-10, 9.414005e-10, 
    9.351268e-10, 9.063109e-10, 1.03804e-09, 1.046536e-09, 1.180027e-09, 
    1.060676e-09, 1.01266e-09, 8.980067e-10, 8.348578e-10, 7.779193e-10, 
    6.628003e-10, 5.49525e-10, 4.156486e-10, 3.353169e-10, 2.881655e-10, 
    3.164695e-10, 2.913828e-10, 3.195245e-10, 3.333664e-10, 2.017503e-10, 
    2.69822e-10, 1.727674e-10, 1.773574e-10, 2.182106e-10, 1.768359e-10, 
    9.307409e-10, 9.671419e-10, 1.101704e-09, 9.953021e-10, 1.19529e-09, 
    1.080006e-09, 1.017564e-09, 8.013373e-10, 7.587947e-10, 7.208327e-10, 
    6.499796e-10, 5.666709e-10, 4.396831e-10, 3.47195e-10, 2.758335e-10, 
    2.806683e-10, 2.789591e-10, 2.644681e-10, 3.013892e-10, 2.587334e-10, 
    2.520224e-10, 2.69834e-10, 1.779785e-10, 2.014808e-10, 1.774558e-10, 
    1.924913e-10, 9.55198e-10, 8.950963e-10, 9.272142e-10, 8.675e-10, 
    9.092586e-10, 7.343043e-10, 6.870517e-10, 4.948713e-10, 5.682287e-10, 
    4.548786e-10, 5.558706e-10, 5.368902e-10, 4.514677e-10, 5.500348e-10, 
    3.518844e-10, 4.791478e-10, 2.63916e-10, 3.681478e-10, 2.581893e-10, 
    2.761172e-10, 2.468996e-10, 2.2267e-10, 1.94665e-10, 1.497113e-10, 
    1.593833e-10, 1.264293e-10, 8.107348e-10, 7.422138e-10, 7.480796e-10, 
    6.806368e-10, 6.337024e-10, 5.401442e-10, 4.116271e-10, 4.570049e-10, 
    3.762841e-10, 3.614152e-10, 4.851567e-10, 4.06072e-10, 6.988027e-10, 
    6.434778e-10, 6.760225e-10, 8.051608e-10, 4.462322e-10, 6.112194e-10, 
    3.340908e-10, 4.031434e-10, 2.260153e-10, 3.049496e-10, 1.64892e-10, 
    1.221319e-10, 8.969955e-11, 6.010963e-11, 7.066736e-10, 7.511304e-10, 
    6.729268e-10, 5.747504e-10, 4.934252e-10, 3.986589e-10, 3.897752e-10, 
    3.738722e-10, 3.348667e-10, 3.044112e-10, 3.689369e-10, 2.97101e-10, 
    6.311008e-10, 4.336403e-10, 7.684508e-10, 6.52743e-10, 5.802315e-10, 
    6.112829e-10, 4.62414e-10, 4.315786e-10, 3.213668e-10, 3.754176e-10, 
    1.31847e-10, 2.177725e-10, 4.279315e-11, 7.327448e-11, 7.671334e-10, 
    7.068282e-10, 5.236862e-10, 6.058415e-10, 3.928474e-10, 3.501451e-10, 
    3.179878e-10, 2.800353e-10, 2.761464e-10, 2.554709e-10, 2.899622e-10, 
    2.567763e-10, 3.984726e-10, 3.296159e-10, 5.426413e-10, 4.836002e-10, 
    5.101506e-10, 5.404691e-10, 4.508976e-10, 3.678493e-10, 3.662161e-10, 
    3.421825e-10, 2.805516e-10, 3.921158e-10, 1.228722e-10, 2.628754e-10, 
    6.451064e-10, 5.458098e-10, 5.326136e-10, 5.689955e-10, 3.542671e-10, 
    4.236721e-10, 2.559623e-10, 2.954235e-10, 2.328388e-10, 2.626047e-10, 
    2.672023e-10, 3.098326e-10, 3.387163e-10, 4.202891e-10, 4.964513e-10, 
    5.636116e-10, 5.474403e-10, 4.755644e-10, 3.631611e-10, 2.757923e-10, 
    2.9347e-10, 2.372264e-10, 4.061106e-10, 3.273309e-10, 3.5633e-10, 
    2.843322e-10, 4.582554e-10, 3.06451e-10, 5.044467e-10, 4.841586e-10, 
    4.251419e-10, 3.224164e-10, 3.023841e-10, 2.819838e-10, 2.944527e-10, 
    3.605883e-10, 3.723656e-10, 4.265138e-10, 4.424097e-10, 4.885252e-10, 
    5.292599e-10, 4.91946e-10, 4.548536e-10, 3.605624e-10, 2.884649e-10, 
    2.223369e-10, 2.079781e-10, 1.483507e-10, 1.957813e-10, 1.222901e-10, 
    1.831627e-10, 8.803826e-11, 2.989685e-10, 1.852373e-10, 4.22591e-10, 
    3.900209e-10, 3.357605e-10, 2.320663e-10, 2.846439e-10, 2.239042e-10, 
    3.728334e-10, 4.732081e-10, 5.020913e-10, 5.593475e-10, 5.008345e-10, 
    5.054197e-10, 4.533708e-10, 4.696513e-10, 3.576981e-10, 4.150934e-10, 
    2.673164e-10, 2.243456e-10, 1.296308e-10, 8.817689e-11, 5.662976e-11, 
    4.565089e-11, 4.263306e-11, 4.141423e-11,
  4.053973e-13, 4.046147e-13, 4.047585e-13, 4.041867e-13, 4.044959e-13, 
    4.041331e-13, 4.052299e-13, 4.045858e-13, 4.049884e-13, 4.053224e-13, 
    4.032521e-13, 4.041627e-13, 4.025111e-13, 4.029432e-13, 4.019818e-13, 
    4.025738e-13, 4.018823e-13, 4.019965e-13, 4.016765e-13, 4.017611e-13, 
    4.01424e-13, 4.016394e-13, 4.012872e-13, 4.014714e-13, 4.014398e-13, 
    4.016472e-13, 4.039625e-13, 4.033543e-13, 4.040015e-13, 4.039081e-13, 
    4.039498e-13, 4.044892e-13, 4.047853e-13, 4.054617e-13, 4.05333e-13, 
    4.048392e-13, 4.038668e-13, 4.041751e-13, 4.034382e-13, 4.034534e-13, 
    4.027758e-13, 4.030635e-13, 4.021252e-13, 4.023559e-13, 4.017574e-13, 
    4.018889e-13, 4.017633e-13, 4.018003e-13, 4.017629e-13, 4.019606e-13, 
    4.018727e-13, 4.020587e-13, 4.030074e-13, 4.026883e-13, 4.037528e-13, 
    4.045715e-13, 4.052001e-13, 4.056906e-13, 4.056189e-13, 4.054844e-13, 
    4.048364e-13, 4.042897e-13, 4.03911e-13, 4.03675e-13, 4.034556e-13, 
    4.02865e-13, 4.025942e-13, 4.020817e-13, 4.021653e-13, 4.020259e-13, 
    4.019026e-13, 4.017158e-13, 4.017449e-13, 4.016684e-13, 4.020295e-13, 
    4.017797e-13, 4.022145e-13, 4.020842e-13, 4.033979e-13, 4.040898e-13, 
    4.04421e-13, 4.047306e-13, 4.055643e-13, 4.04976e-13, 4.052011e-13, 
    4.046797e-13, 4.043728e-13, 4.045222e-13, 4.036688e-13, 4.039814e-13, 
    4.025791e-13, 4.031115e-13, 4.019165e-13, 4.021478e-13, 4.018656e-13, 
    4.020037e-13, 4.017742e-13, 4.019792e-13, 4.016412e-13, 4.015779e-13, 
    4.016208e-13, 4.014648e-13, 4.019914e-13, 4.017633e-13, 4.045265e-13, 
    4.045018e-13, 4.043883e-13, 4.049069e-13, 4.049403e-13, 4.054652e-13, 
    4.049959e-13, 4.04807e-13, 4.043556e-13, 4.041067e-13, 4.038822e-13, 
    4.034279e-13, 4.029802e-13, 4.024503e-13, 4.021319e-13, 4.019447e-13, 
    4.020571e-13, 4.019575e-13, 4.020692e-13, 4.021241e-13, 4.016012e-13, 
    4.018718e-13, 4.014858e-13, 4.015041e-13, 4.016667e-13, 4.01502e-13, 
    4.044845e-13, 4.046278e-13, 4.051573e-13, 4.047387e-13, 4.055252e-13, 
    4.05072e-13, 4.048263e-13, 4.039746e-13, 4.038068e-13, 4.03657e-13, 
    4.033773e-13, 4.03048e-13, 4.025455e-13, 4.02179e-13, 4.018957e-13, 
    4.019149e-13, 4.019081e-13, 4.018506e-13, 4.019972e-13, 4.018278e-13, 
    4.018011e-13, 4.018719e-13, 4.015066e-13, 4.016001e-13, 4.015045e-13, 
    4.015644e-13, 4.045808e-13, 4.043441e-13, 4.044706e-13, 4.042354e-13, 
    4.043999e-13, 4.037101e-13, 4.035237e-13, 4.02764e-13, 4.030542e-13, 
    4.026057e-13, 4.030053e-13, 4.029303e-13, 4.025922e-13, 4.029823e-13, 
    4.021976e-13, 4.027018e-13, 4.018484e-13, 4.02262e-13, 4.018256e-13, 
    4.018969e-13, 4.017808e-13, 4.016844e-13, 4.01573e-13, 4.01394e-13, 
    4.014325e-13, 4.013011e-13, 4.040116e-13, 4.037414e-13, 4.037645e-13, 
    4.034983e-13, 4.03313e-13, 4.029431e-13, 4.024344e-13, 4.026141e-13, 
    4.022943e-13, 4.022354e-13, 4.027256e-13, 4.024124e-13, 4.0357e-13, 
    4.033516e-13, 4.034801e-13, 4.039896e-13, 4.025715e-13, 4.032241e-13, 
    4.02127e-13, 4.024008e-13, 4.016977e-13, 4.020114e-13, 4.014545e-13, 
    4.01284e-13, 4.011546e-13, 4.010364e-13, 4.036011e-13, 4.037765e-13, 
    4.034679e-13, 4.0308e-13, 4.027583e-13, 4.02383e-13, 4.023478e-13, 
    4.022848e-13, 4.021301e-13, 4.020092e-13, 4.022652e-13, 4.019802e-13, 
    4.033027e-13, 4.025216e-13, 4.038449e-13, 4.033882e-13, 4.031017e-13, 
    4.032244e-13, 4.026356e-13, 4.025134e-13, 4.020765e-13, 4.022909e-13, 
    4.013228e-13, 4.016649e-13, 4.009671e-13, 4.01089e-13, 4.038397e-13, 
    4.036017e-13, 4.02878e-13, 4.032029e-13, 4.023599e-13, 4.021907e-13, 
    4.020631e-13, 4.019124e-13, 4.01897e-13, 4.018148e-13, 4.019518e-13, 
    4.0182e-13, 4.023823e-13, 4.021092e-13, 4.02953e-13, 4.027194e-13, 
    4.028245e-13, 4.029444e-13, 4.025899e-13, 4.022609e-13, 4.022544e-13, 
    4.021591e-13, 4.019145e-13, 4.023571e-13, 4.01287e-13, 4.018442e-13, 
    4.03358e-13, 4.029656e-13, 4.029134e-13, 4.030572e-13, 4.02207e-13, 
    4.024821e-13, 4.018168e-13, 4.019735e-13, 4.017249e-13, 4.018432e-13, 
    4.018614e-13, 4.020307e-13, 4.021453e-13, 4.024687e-13, 4.027703e-13, 
    4.030359e-13, 4.02972e-13, 4.026876e-13, 4.022423e-13, 4.018956e-13, 
    4.019658e-13, 4.017423e-13, 4.024125e-13, 4.021002e-13, 4.022152e-13, 
    4.019295e-13, 4.026191e-13, 4.020173e-13, 4.028019e-13, 4.027216e-13, 
    4.024879e-13, 4.020807e-13, 4.020012e-13, 4.019201e-13, 4.019697e-13, 
    4.022321e-13, 4.022788e-13, 4.024934e-13, 4.025563e-13, 4.027389e-13, 
    4.029001e-13, 4.027525e-13, 4.026056e-13, 4.02232e-13, 4.019459e-13, 
    4.016831e-13, 4.01626e-13, 4.013886e-13, 4.015775e-13, 4.012846e-13, 
    4.015272e-13, 4.011479e-13, 4.019876e-13, 4.015355e-13, 4.024778e-13, 
    4.023488e-13, 4.021336e-13, 4.017218e-13, 4.019307e-13, 4.016893e-13, 
    4.022806e-13, 4.026783e-13, 4.027926e-13, 4.030191e-13, 4.027876e-13, 
    4.028058e-13, 4.025997e-13, 4.026642e-13, 4.022206e-13, 4.024481e-13, 
    4.018619e-13, 4.016911e-13, 4.013139e-13, 4.011485e-13, 4.010224e-13, 
    4.009785e-13, 4.009665e-13, 4.009616e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949659e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 
    8.949657e-07, 8.949658e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949658e-07, 8.949657e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949658e-07, 
    8.949658e-07, 8.949659e-07, 8.949659e-07, 8.949659e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949657e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949656e-07, 8.949657e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 
    8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949659e-07, 
    8.949659e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949657e-07, 8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 
    8.949657e-07, 8.949657e-07, 8.949658e-07, 8.949656e-07, 8.949657e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949657e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949657e-07, 8.949656e-07, 8.949658e-07, 8.949657e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 
    8.949654e-07, 8.949655e-07, 8.949652e-07, 8.949653e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949654e-07, 8.949655e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949655e-07, 8.949654e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.708882e-16, 6.727296e-16, 6.723719e-16, 6.73856e-16, 6.730331e-16, 
    6.740046e-16, 6.712619e-16, 6.728025e-16, 6.718193e-16, 6.710544e-16, 
    6.767327e-16, 6.739223e-16, 6.796512e-16, 6.77861e-16, 6.823563e-16, 
    6.793724e-16, 6.829576e-16, 6.82271e-16, 6.843386e-16, 6.837465e-16, 
    6.863875e-16, 6.846118e-16, 6.877564e-16, 6.85964e-16, 6.862442e-16, 
    6.845531e-16, 6.744888e-16, 6.763828e-16, 6.743763e-16, 6.746465e-16, 
    6.745255e-16, 6.730499e-16, 6.723055e-16, 6.707478e-16, 6.710308e-16, 
    6.721751e-16, 6.747681e-16, 6.738886e-16, 6.761058e-16, 6.760557e-16, 
    6.785212e-16, 6.774099e-16, 6.815503e-16, 6.803745e-16, 6.837713e-16, 
    6.829174e-16, 6.83731e-16, 6.834844e-16, 6.837343e-16, 6.824819e-16, 
    6.830185e-16, 6.819164e-16, 6.776179e-16, 6.788819e-16, 6.751099e-16, 
    6.728379e-16, 6.713294e-16, 6.702579e-16, 6.704094e-16, 6.70698e-16, 
    6.721817e-16, 6.735765e-16, 6.746388e-16, 6.753489e-16, 6.760485e-16, 
    6.781632e-16, 6.792832e-16, 6.817877e-16, 6.813365e-16, 6.821013e-16, 
    6.828325e-16, 6.840587e-16, 6.83857e-16, 6.84397e-16, 6.820815e-16, 
    6.836204e-16, 6.810793e-16, 6.817745e-16, 6.762364e-16, 6.74126e-16, 
    6.732265e-16, 6.724406e-16, 6.705258e-16, 6.718481e-16, 6.713269e-16, 
    6.725673e-16, 6.733548e-16, 6.729654e-16, 6.753683e-16, 6.744343e-16, 
    6.793495e-16, 6.772337e-16, 6.827472e-16, 6.814292e-16, 6.830631e-16, 
    6.822296e-16, 6.836573e-16, 6.823724e-16, 6.845981e-16, 6.850822e-16, 
    6.847513e-16, 6.860226e-16, 6.823011e-16, 6.837308e-16, 6.729544e-16, 
    6.730179e-16, 6.73314e-16, 6.720123e-16, 6.719328e-16, 6.707399e-16, 
    6.718015e-16, 6.722533e-16, 6.734006e-16, 6.740786e-16, 6.74723e-16, 
    6.761394e-16, 6.777198e-16, 6.799287e-16, 6.815146e-16, 6.825769e-16, 
    6.819257e-16, 6.825007e-16, 6.818579e-16, 6.815566e-16, 6.849006e-16, 
    6.830234e-16, 6.858398e-16, 6.856841e-16, 6.844097e-16, 6.857017e-16, 
    6.730625e-16, 6.72697e-16, 6.71427e-16, 6.72421e-16, 6.706101e-16, 
    6.716236e-16, 6.72206e-16, 6.744534e-16, 6.749474e-16, 6.754047e-16, 
    6.763081e-16, 6.774668e-16, 6.794978e-16, 6.812638e-16, 6.828751e-16, 
    6.827571e-16, 6.827986e-16, 6.831582e-16, 6.822671e-16, 6.833044e-16, 
    6.834783e-16, 6.830234e-16, 6.856633e-16, 6.849095e-16, 6.856808e-16, 
    6.851901e-16, 6.728159e-16, 6.734309e-16, 6.730985e-16, 6.737233e-16, 
    6.73283e-16, 6.752397e-16, 6.75826e-16, 6.785683e-16, 6.774438e-16, 
    6.792339e-16, 6.776259e-16, 6.779108e-16, 6.792913e-16, 6.77713e-16, 
    6.811661e-16, 6.788247e-16, 6.831721e-16, 6.808353e-16, 6.833185e-16, 
    6.828681e-16, 6.836139e-16, 6.842814e-16, 6.851213e-16, 6.866694e-16, 
    6.863111e-16, 6.876055e-16, 6.743477e-16, 6.751446e-16, 6.750749e-16, 
    6.759089e-16, 6.765255e-16, 6.778618e-16, 6.800029e-16, 6.791981e-16, 
    6.806758e-16, 6.809722e-16, 6.787274e-16, 6.801055e-16, 6.756781e-16, 
    6.763936e-16, 6.759679e-16, 6.744103e-16, 6.79383e-16, 6.768321e-16, 
    6.815407e-16, 6.801606e-16, 6.841862e-16, 6.821847e-16, 6.861138e-16, 
    6.877901e-16, 6.893685e-16, 6.912091e-16, 6.755799e-16, 6.750385e-16, 
    6.760082e-16, 6.773484e-16, 6.785925e-16, 6.802447e-16, 6.804139e-16, 
    6.807231e-16, 6.815245e-16, 6.821978e-16, 6.808205e-16, 6.823666e-16, 
    6.765586e-16, 6.796045e-16, 6.748334e-16, 6.762705e-16, 6.772697e-16, 
    6.768318e-16, 6.791062e-16, 6.796418e-16, 6.818167e-16, 6.806929e-16, 
    6.873761e-16, 6.844218e-16, 6.926108e-16, 6.903254e-16, 6.748491e-16, 
    6.755782e-16, 6.781132e-16, 6.769075e-16, 6.803552e-16, 6.812028e-16, 
    6.81892e-16, 6.82772e-16, 6.828673e-16, 6.833886e-16, 6.825343e-16, 
    6.83355e-16, 6.802482e-16, 6.816372e-16, 6.778241e-16, 6.787525e-16, 
    6.783256e-16, 6.77857e-16, 6.793031e-16, 6.808421e-16, 6.808756e-16, 
    6.813688e-16, 6.827565e-16, 6.803692e-16, 6.877558e-16, 6.831958e-16, 
    6.76373e-16, 6.777752e-16, 6.779762e-16, 6.774331e-16, 6.811178e-16, 
    6.797833e-16, 6.83376e-16, 6.824057e-16, 6.839954e-16, 6.832056e-16, 
    6.830893e-16, 6.820745e-16, 6.814423e-16, 6.798444e-16, 6.785436e-16, 
    6.77512e-16, 6.777519e-16, 6.78885e-16, 6.809364e-16, 6.828756e-16, 
    6.824509e-16, 6.838747e-16, 6.801054e-16, 6.816863e-16, 6.810752e-16, 
    6.826685e-16, 6.791766e-16, 6.821483e-16, 6.784161e-16, 6.787437e-16, 
    6.797568e-16, 6.81793e-16, 6.822443e-16, 6.827248e-16, 6.824285e-16, 
    6.809885e-16, 6.807528e-16, 6.797323e-16, 6.794502e-16, 6.786724e-16, 
    6.78028e-16, 6.786166e-16, 6.792345e-16, 6.809894e-16, 6.825693e-16, 
    6.842908e-16, 6.847122e-16, 6.867196e-16, 6.850846e-16, 6.87781e-16, 
    6.854874e-16, 6.894569e-16, 6.823215e-16, 6.854213e-16, 6.798031e-16, 
    6.804092e-16, 6.815044e-16, 6.840156e-16, 6.82661e-16, 6.842454e-16, 
    6.807437e-16, 6.789238e-16, 6.784535e-16, 6.775745e-16, 6.784737e-16, 
    6.784005e-16, 6.792605e-16, 6.789843e-16, 6.810477e-16, 6.799396e-16, 
    6.830862e-16, 6.842331e-16, 6.874697e-16, 6.894508e-16, 6.914665e-16, 
    6.923554e-16, 6.926259e-16, 6.92739e-16 ;

 CWDC_TO_LITR2C =
  5.09875e-16, 5.112745e-16, 5.110026e-16, 5.121306e-16, 5.115051e-16, 
    5.122434e-16, 5.101591e-16, 5.113299e-16, 5.105827e-16, 5.100013e-16, 
    5.143168e-16, 5.121809e-16, 5.165349e-16, 5.151744e-16, 5.185908e-16, 
    5.16323e-16, 5.190478e-16, 5.185259e-16, 5.200973e-16, 5.196474e-16, 
    5.216546e-16, 5.20305e-16, 5.226949e-16, 5.213326e-16, 5.215456e-16, 
    5.202604e-16, 5.126115e-16, 5.140509e-16, 5.12526e-16, 5.127314e-16, 
    5.126394e-16, 5.115179e-16, 5.109522e-16, 5.097684e-16, 5.099834e-16, 
    5.10853e-16, 5.128238e-16, 5.121553e-16, 5.138404e-16, 5.138024e-16, 
    5.156761e-16, 5.148315e-16, 5.179783e-16, 5.170846e-16, 5.196661e-16, 
    5.190172e-16, 5.196356e-16, 5.194482e-16, 5.19638e-16, 5.186862e-16, 
    5.190941e-16, 5.182565e-16, 5.149896e-16, 5.159502e-16, 5.130835e-16, 
    5.113568e-16, 5.102103e-16, 5.09396e-16, 5.095111e-16, 5.097305e-16, 
    5.108581e-16, 5.119182e-16, 5.127255e-16, 5.132652e-16, 5.137969e-16, 
    5.15404e-16, 5.162552e-16, 5.181586e-16, 5.178158e-16, 5.18397e-16, 
    5.189527e-16, 5.198846e-16, 5.197313e-16, 5.201417e-16, 5.183819e-16, 
    5.195515e-16, 5.176203e-16, 5.181487e-16, 5.139397e-16, 5.123358e-16, 
    5.116522e-16, 5.110548e-16, 5.095996e-16, 5.106046e-16, 5.102084e-16, 
    5.111511e-16, 5.117496e-16, 5.114537e-16, 5.132799e-16, 5.125701e-16, 
    5.163057e-16, 5.146976e-16, 5.188879e-16, 5.178862e-16, 5.191279e-16, 
    5.184945e-16, 5.195796e-16, 5.186031e-16, 5.202945e-16, 5.206624e-16, 
    5.20411e-16, 5.213772e-16, 5.185489e-16, 5.196354e-16, 5.114453e-16, 
    5.114936e-16, 5.117186e-16, 5.107293e-16, 5.106689e-16, 5.097624e-16, 
    5.105692e-16, 5.109125e-16, 5.117845e-16, 5.122997e-16, 5.127895e-16, 
    5.138659e-16, 5.150671e-16, 5.167458e-16, 5.179511e-16, 5.187585e-16, 
    5.182636e-16, 5.187005e-16, 5.18212e-16, 5.17983e-16, 5.205245e-16, 
    5.190978e-16, 5.212382e-16, 5.211199e-16, 5.201514e-16, 5.211333e-16, 
    5.115275e-16, 5.112498e-16, 5.102845e-16, 5.1104e-16, 5.096636e-16, 
    5.104339e-16, 5.108766e-16, 5.125846e-16, 5.1296e-16, 5.133076e-16, 
    5.139942e-16, 5.148747e-16, 5.164183e-16, 5.177605e-16, 5.189851e-16, 
    5.188954e-16, 5.18927e-16, 5.192002e-16, 5.18523e-16, 5.193114e-16, 
    5.194435e-16, 5.190978e-16, 5.211041e-16, 5.205312e-16, 5.211174e-16, 
    5.207445e-16, 5.113401e-16, 5.118075e-16, 5.115549e-16, 5.120297e-16, 
    5.116951e-16, 5.131822e-16, 5.136278e-16, 5.157119e-16, 5.148573e-16, 
    5.162177e-16, 5.149957e-16, 5.152122e-16, 5.162613e-16, 5.150619e-16, 
    5.176862e-16, 5.159068e-16, 5.192109e-16, 5.174348e-16, 5.19322e-16, 
    5.189798e-16, 5.195466e-16, 5.200539e-16, 5.206922e-16, 5.218688e-16, 
    5.215965e-16, 5.225802e-16, 5.125042e-16, 5.131099e-16, 5.130569e-16, 
    5.136908e-16, 5.141594e-16, 5.151749e-16, 5.168022e-16, 5.161906e-16, 
    5.173136e-16, 5.175389e-16, 5.158328e-16, 5.168802e-16, 5.135154e-16, 
    5.140591e-16, 5.137356e-16, 5.125518e-16, 5.163311e-16, 5.143924e-16, 
    5.17971e-16, 5.16922e-16, 5.199815e-16, 5.184603e-16, 5.214465e-16, 
    5.227204e-16, 5.2392e-16, 5.253189e-16, 5.134407e-16, 5.130292e-16, 
    5.137662e-16, 5.147848e-16, 5.157303e-16, 5.16986e-16, 5.171146e-16, 
    5.173496e-16, 5.179586e-16, 5.184703e-16, 5.174236e-16, 5.185986e-16, 
    5.141845e-16, 5.164994e-16, 5.128734e-16, 5.139656e-16, 5.147249e-16, 
    5.143922e-16, 5.161207e-16, 5.165277e-16, 5.181807e-16, 5.173266e-16, 
    5.224058e-16, 5.201606e-16, 5.263842e-16, 5.246473e-16, 5.128854e-16, 
    5.134395e-16, 5.153661e-16, 5.144497e-16, 5.170699e-16, 5.177141e-16, 
    5.182379e-16, 5.189067e-16, 5.189792e-16, 5.193753e-16, 5.18726e-16, 
    5.193498e-16, 5.169886e-16, 5.180442e-16, 5.151464e-16, 5.15852e-16, 
    5.155275e-16, 5.151713e-16, 5.162703e-16, 5.1744e-16, 5.174655e-16, 
    5.178403e-16, 5.188949e-16, 5.170805e-16, 5.226944e-16, 5.192288e-16, 
    5.140434e-16, 5.151092e-16, 5.152619e-16, 5.148491e-16, 5.176495e-16, 
    5.166353e-16, 5.193657e-16, 5.186284e-16, 5.198365e-16, 5.192362e-16, 
    5.191479e-16, 5.183766e-16, 5.178962e-16, 5.166817e-16, 5.156931e-16, 
    5.149091e-16, 5.150915e-16, 5.159526e-16, 5.175116e-16, 5.189855e-16, 
    5.186627e-16, 5.197447e-16, 5.1688e-16, 5.180816e-16, 5.176171e-16, 
    5.18828e-16, 5.161742e-16, 5.184328e-16, 5.155962e-16, 5.158452e-16, 
    5.166152e-16, 5.181627e-16, 5.185057e-16, 5.188708e-16, 5.186456e-16, 
    5.175513e-16, 5.173722e-16, 5.165966e-16, 5.163821e-16, 5.15791e-16, 
    5.153013e-16, 5.157486e-16, 5.162182e-16, 5.17552e-16, 5.187527e-16, 
    5.20061e-16, 5.203813e-16, 5.219069e-16, 5.206643e-16, 5.227136e-16, 
    5.209704e-16, 5.239872e-16, 5.185643e-16, 5.209202e-16, 5.166504e-16, 
    5.17111e-16, 5.179433e-16, 5.198519e-16, 5.188223e-16, 5.200266e-16, 
    5.173652e-16, 5.159821e-16, 5.156247e-16, 5.149566e-16, 5.1564e-16, 
    5.155844e-16, 5.16238e-16, 5.16028e-16, 5.175962e-16, 5.16754e-16, 
    5.191455e-16, 5.200172e-16, 5.224769e-16, 5.239826e-16, 5.255145e-16, 
    5.261901e-16, 5.263957e-16, 5.264816e-16 ;

 CWDC_TO_LITR3C =
  1.610132e-16, 1.614551e-16, 1.613693e-16, 1.617254e-16, 1.615279e-16, 
    1.617611e-16, 1.611029e-16, 1.614726e-16, 1.612366e-16, 1.610531e-16, 
    1.624158e-16, 1.617414e-16, 1.631163e-16, 1.626866e-16, 1.637655e-16, 
    1.630494e-16, 1.639098e-16, 1.63745e-16, 1.642413e-16, 1.640992e-16, 
    1.64733e-16, 1.643068e-16, 1.650615e-16, 1.646314e-16, 1.646986e-16, 
    1.642927e-16, 1.618773e-16, 1.623319e-16, 1.618503e-16, 1.619152e-16, 
    1.618861e-16, 1.61532e-16, 1.613533e-16, 1.609795e-16, 1.610474e-16, 
    1.61322e-16, 1.619443e-16, 1.617333e-16, 1.622654e-16, 1.622534e-16, 
    1.628451e-16, 1.625784e-16, 1.635721e-16, 1.632899e-16, 1.641051e-16, 
    1.639002e-16, 1.640954e-16, 1.640363e-16, 1.640962e-16, 1.637957e-16, 
    1.639244e-16, 1.636599e-16, 1.626283e-16, 1.629316e-16, 1.620264e-16, 
    1.614811e-16, 1.61119e-16, 1.608619e-16, 1.608982e-16, 1.609675e-16, 
    1.613236e-16, 1.616584e-16, 1.619133e-16, 1.620837e-16, 1.622516e-16, 
    1.627592e-16, 1.63028e-16, 1.636291e-16, 1.635208e-16, 1.637043e-16, 
    1.638798e-16, 1.641741e-16, 1.641257e-16, 1.642553e-16, 1.636996e-16, 
    1.640689e-16, 1.63459e-16, 1.636259e-16, 1.622967e-16, 1.617902e-16, 
    1.615744e-16, 1.613857e-16, 1.609262e-16, 1.612435e-16, 1.611185e-16, 
    1.614161e-16, 1.616052e-16, 1.615117e-16, 1.620884e-16, 1.618642e-16, 
    1.630439e-16, 1.625361e-16, 1.638593e-16, 1.63543e-16, 1.639351e-16, 
    1.637351e-16, 1.640778e-16, 1.637694e-16, 1.643035e-16, 1.644197e-16, 
    1.643403e-16, 1.646454e-16, 1.637523e-16, 1.640954e-16, 1.615091e-16, 
    1.615243e-16, 1.615953e-16, 1.612829e-16, 1.612639e-16, 1.609776e-16, 
    1.612324e-16, 1.613408e-16, 1.616161e-16, 1.617789e-16, 1.619335e-16, 
    1.622734e-16, 1.626528e-16, 1.631829e-16, 1.635635e-16, 1.638185e-16, 
    1.636622e-16, 1.638002e-16, 1.636459e-16, 1.635736e-16, 1.643762e-16, 
    1.639256e-16, 1.646016e-16, 1.645642e-16, 1.642583e-16, 1.645684e-16, 
    1.61535e-16, 1.614473e-16, 1.611425e-16, 1.61381e-16, 1.609464e-16, 
    1.611897e-16, 1.613295e-16, 1.618688e-16, 1.619874e-16, 1.620971e-16, 
    1.623139e-16, 1.62592e-16, 1.630795e-16, 1.635033e-16, 1.6389e-16, 
    1.638617e-16, 1.638717e-16, 1.63958e-16, 1.637441e-16, 1.639931e-16, 
    1.640348e-16, 1.639256e-16, 1.645592e-16, 1.643783e-16, 1.645634e-16, 
    1.644456e-16, 1.614758e-16, 1.616234e-16, 1.615437e-16, 1.616936e-16, 
    1.615879e-16, 1.620575e-16, 1.621982e-16, 1.628564e-16, 1.625865e-16, 
    1.630161e-16, 1.626302e-16, 1.626986e-16, 1.630299e-16, 1.626511e-16, 
    1.634798e-16, 1.629179e-16, 1.639613e-16, 1.634005e-16, 1.639964e-16, 
    1.638884e-16, 1.640673e-16, 1.642275e-16, 1.644291e-16, 1.648007e-16, 
    1.647147e-16, 1.650253e-16, 1.618434e-16, 1.620347e-16, 1.62018e-16, 
    1.622181e-16, 1.623661e-16, 1.626868e-16, 1.632007e-16, 1.630075e-16, 
    1.633622e-16, 1.634333e-16, 1.628946e-16, 1.632253e-16, 1.621628e-16, 
    1.623345e-16, 1.622323e-16, 1.618585e-16, 1.630519e-16, 1.624397e-16, 
    1.635698e-16, 1.632385e-16, 1.642047e-16, 1.637243e-16, 1.646673e-16, 
    1.650696e-16, 1.654484e-16, 1.658902e-16, 1.621392e-16, 1.620092e-16, 
    1.62242e-16, 1.625636e-16, 1.628622e-16, 1.632587e-16, 1.632993e-16, 
    1.633736e-16, 1.635659e-16, 1.637275e-16, 1.633969e-16, 1.63768e-16, 
    1.623741e-16, 1.631051e-16, 1.6196e-16, 1.623049e-16, 1.625447e-16, 
    1.624396e-16, 1.629855e-16, 1.63114e-16, 1.63636e-16, 1.633663e-16, 
    1.649703e-16, 1.642612e-16, 1.662266e-16, 1.656781e-16, 1.619638e-16, 
    1.621388e-16, 1.627472e-16, 1.624578e-16, 1.632852e-16, 1.634887e-16, 
    1.636541e-16, 1.638653e-16, 1.638882e-16, 1.640133e-16, 1.638082e-16, 
    1.640052e-16, 1.632596e-16, 1.635929e-16, 1.626778e-16, 1.629006e-16, 
    1.627982e-16, 1.626857e-16, 1.630327e-16, 1.634021e-16, 1.634102e-16, 
    1.635285e-16, 1.638616e-16, 1.632886e-16, 1.650614e-16, 1.63967e-16, 
    1.623295e-16, 1.62666e-16, 1.627143e-16, 1.625839e-16, 1.634683e-16, 
    1.63148e-16, 1.640102e-16, 1.637774e-16, 1.641589e-16, 1.639693e-16, 
    1.639414e-16, 1.636979e-16, 1.635462e-16, 1.631626e-16, 1.628505e-16, 
    1.626029e-16, 1.626605e-16, 1.629324e-16, 1.634247e-16, 1.638902e-16, 
    1.637882e-16, 1.641299e-16, 1.632253e-16, 1.636047e-16, 1.63458e-16, 
    1.638404e-16, 1.630024e-16, 1.637156e-16, 1.628199e-16, 1.628985e-16, 
    1.631416e-16, 1.636303e-16, 1.637386e-16, 1.638539e-16, 1.637828e-16, 
    1.634372e-16, 1.633807e-16, 1.631358e-16, 1.63068e-16, 1.628814e-16, 
    1.627267e-16, 1.62868e-16, 1.630163e-16, 1.634375e-16, 1.638166e-16, 
    1.642298e-16, 1.643309e-16, 1.648127e-16, 1.644203e-16, 1.650674e-16, 
    1.64517e-16, 1.654696e-16, 1.637572e-16, 1.645011e-16, 1.631527e-16, 
    1.632982e-16, 1.635611e-16, 1.641637e-16, 1.638386e-16, 1.642189e-16, 
    1.633785e-16, 1.629417e-16, 1.628288e-16, 1.626179e-16, 1.628337e-16, 
    1.628161e-16, 1.630225e-16, 1.629562e-16, 1.634514e-16, 1.631855e-16, 
    1.639407e-16, 1.642159e-16, 1.649927e-16, 1.654682e-16, 1.65952e-16, 
    1.661653e-16, 1.662302e-16, 1.662573e-16 ;

 CWDC_vr =
  5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110348e-05, 5.110348e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110348e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110348e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110347e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789932e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789932e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.01975e-18, 1.022549e-18, 1.022005e-18, 1.024261e-18, 1.02301e-18, 
    1.024487e-18, 1.020318e-18, 1.02266e-18, 1.021165e-18, 1.020003e-18, 
    1.028634e-18, 1.024362e-18, 1.03307e-18, 1.030349e-18, 1.037182e-18, 
    1.032646e-18, 1.038096e-18, 1.037052e-18, 1.040195e-18, 1.039295e-18, 
    1.043309e-18, 1.04061e-18, 1.04539e-18, 1.042665e-18, 1.043091e-18, 
    1.040521e-18, 1.025223e-18, 1.028102e-18, 1.025052e-18, 1.025463e-18, 
    1.025279e-18, 1.023036e-18, 1.021904e-18, 1.019537e-18, 1.019967e-18, 
    1.021706e-18, 1.025648e-18, 1.024311e-18, 1.027681e-18, 1.027605e-18, 
    1.031352e-18, 1.029663e-18, 1.035957e-18, 1.034169e-18, 1.039332e-18, 
    1.038034e-18, 1.039271e-18, 1.038896e-18, 1.039276e-18, 1.037372e-18, 
    1.038188e-18, 1.036513e-18, 1.029979e-18, 1.0319e-18, 1.026167e-18, 
    1.022714e-18, 1.020421e-18, 1.018792e-18, 1.019022e-18, 1.019461e-18, 
    1.021716e-18, 1.023836e-18, 1.025451e-18, 1.02653e-18, 1.027594e-18, 
    1.030808e-18, 1.03251e-18, 1.036317e-18, 1.035631e-18, 1.036794e-18, 
    1.037905e-18, 1.039769e-18, 1.039463e-18, 1.040283e-18, 1.036764e-18, 
    1.039103e-18, 1.035241e-18, 1.036297e-18, 1.027879e-18, 1.024672e-18, 
    1.023304e-18, 1.02211e-18, 1.019199e-18, 1.021209e-18, 1.020417e-18, 
    1.022302e-18, 1.023499e-18, 1.022907e-18, 1.02656e-18, 1.02514e-18, 
    1.032611e-18, 1.029395e-18, 1.037776e-18, 1.035772e-18, 1.038256e-18, 
    1.036989e-18, 1.039159e-18, 1.037206e-18, 1.040589e-18, 1.041325e-18, 
    1.040822e-18, 1.042754e-18, 1.037098e-18, 1.039271e-18, 1.022891e-18, 
    1.022987e-18, 1.023437e-18, 1.021459e-18, 1.021338e-18, 1.019525e-18, 
    1.021138e-18, 1.021825e-18, 1.023569e-18, 1.024599e-18, 1.025579e-18, 
    1.027732e-18, 1.030134e-18, 1.033492e-18, 1.035902e-18, 1.037517e-18, 
    1.036527e-18, 1.037401e-18, 1.036424e-18, 1.035966e-18, 1.041049e-18, 
    1.038196e-18, 1.042476e-18, 1.04224e-18, 1.040303e-18, 1.042267e-18, 
    1.023055e-18, 1.022499e-18, 1.020569e-18, 1.02208e-18, 1.019327e-18, 
    1.020868e-18, 1.021753e-18, 1.025169e-18, 1.02592e-18, 1.026615e-18, 
    1.027988e-18, 1.029749e-18, 1.032837e-18, 1.035521e-18, 1.03797e-18, 
    1.037791e-18, 1.037854e-18, 1.0384e-18, 1.037046e-18, 1.038623e-18, 
    1.038887e-18, 1.038196e-18, 1.042208e-18, 1.041062e-18, 1.042235e-18, 
    1.041489e-18, 1.02268e-18, 1.023615e-18, 1.02311e-18, 1.02406e-18, 
    1.02339e-18, 1.026364e-18, 1.027256e-18, 1.031424e-18, 1.029715e-18, 
    1.032435e-18, 1.029991e-18, 1.030424e-18, 1.032523e-18, 1.030124e-18, 
    1.035372e-18, 1.031814e-18, 1.038422e-18, 1.03487e-18, 1.038644e-18, 
    1.03796e-18, 1.039093e-18, 1.040108e-18, 1.041384e-18, 1.043738e-18, 
    1.043193e-18, 1.04516e-18, 1.025008e-18, 1.02622e-18, 1.026114e-18, 
    1.027382e-18, 1.028319e-18, 1.03035e-18, 1.033604e-18, 1.032381e-18, 
    1.034627e-18, 1.035078e-18, 1.031666e-18, 1.03376e-18, 1.027031e-18, 
    1.028118e-18, 1.027471e-18, 1.025104e-18, 1.032662e-18, 1.028785e-18, 
    1.035942e-18, 1.033844e-18, 1.039963e-18, 1.036921e-18, 1.042893e-18, 
    1.045441e-18, 1.04784e-18, 1.050638e-18, 1.026881e-18, 1.026059e-18, 
    1.027532e-18, 1.02957e-18, 1.031461e-18, 1.033972e-18, 1.034229e-18, 
    1.034699e-18, 1.035917e-18, 1.036941e-18, 1.034847e-18, 1.037197e-18, 
    1.028369e-18, 1.032999e-18, 1.025747e-18, 1.027931e-18, 1.02945e-18, 
    1.028784e-18, 1.032241e-18, 1.033056e-18, 1.036361e-18, 1.034653e-18, 
    1.044812e-18, 1.040321e-18, 1.052768e-18, 1.049295e-18, 1.025771e-18, 
    1.026879e-18, 1.030732e-18, 1.028899e-18, 1.03414e-18, 1.035428e-18, 
    1.036476e-18, 1.037813e-18, 1.037958e-18, 1.038751e-18, 1.037452e-18, 
    1.0387e-18, 1.033977e-18, 1.036088e-18, 1.030293e-18, 1.031704e-18, 
    1.031055e-18, 1.030343e-18, 1.032541e-18, 1.03488e-18, 1.034931e-18, 
    1.03568e-18, 1.03779e-18, 1.034161e-18, 1.045389e-18, 1.038458e-18, 
    1.028087e-18, 1.030218e-18, 1.030524e-18, 1.029698e-18, 1.035299e-18, 
    1.033271e-18, 1.038731e-18, 1.037257e-18, 1.039673e-18, 1.038472e-18, 
    1.038296e-18, 1.036753e-18, 1.035792e-18, 1.033363e-18, 1.031386e-18, 
    1.029818e-18, 1.030183e-18, 1.031905e-18, 1.035023e-18, 1.037971e-18, 
    1.037325e-18, 1.039489e-18, 1.03376e-18, 1.036163e-18, 1.035234e-18, 
    1.037656e-18, 1.032348e-18, 1.036866e-18, 1.031192e-18, 1.03169e-18, 
    1.03323e-18, 1.036325e-18, 1.037011e-18, 1.037742e-18, 1.037291e-18, 
    1.035103e-18, 1.034744e-18, 1.033193e-18, 1.032764e-18, 1.031582e-18, 
    1.030603e-18, 1.031497e-18, 1.032436e-18, 1.035104e-18, 1.037505e-18, 
    1.040122e-18, 1.040762e-18, 1.043814e-18, 1.041329e-18, 1.045427e-18, 
    1.041941e-18, 1.047974e-18, 1.037129e-18, 1.04184e-18, 1.033301e-18, 
    1.034222e-18, 1.035887e-18, 1.039704e-18, 1.037645e-18, 1.040053e-18, 
    1.03473e-18, 1.031964e-18, 1.031249e-18, 1.029913e-18, 1.03128e-18, 
    1.031169e-18, 1.032476e-18, 1.032056e-18, 1.035192e-18, 1.033508e-18, 
    1.038291e-18, 1.040034e-18, 1.044954e-18, 1.047965e-18, 1.051029e-18, 
    1.05238e-18, 1.052791e-18, 1.052963e-18 ;

 CWDN_TO_LITR3N =
  3.220263e-19, 3.229102e-19, 3.227385e-19, 3.234509e-19, 3.230559e-19, 
    3.235222e-19, 3.222057e-19, 3.229452e-19, 3.224733e-19, 3.221061e-19, 
    3.248317e-19, 3.234827e-19, 3.262326e-19, 3.253733e-19, 3.27531e-19, 
    3.260987e-19, 3.278197e-19, 3.274901e-19, 3.284825e-19, 3.281983e-19, 
    3.29466e-19, 3.286137e-19, 3.301231e-19, 3.292627e-19, 3.293972e-19, 
    3.285855e-19, 3.237546e-19, 3.246637e-19, 3.237006e-19, 3.238304e-19, 
    3.237722e-19, 3.230639e-19, 3.227066e-19, 3.21959e-19, 3.220948e-19, 
    3.22644e-19, 3.238887e-19, 3.234665e-19, 3.245308e-19, 3.245068e-19, 
    3.256902e-19, 3.251567e-19, 3.271442e-19, 3.265797e-19, 3.282102e-19, 
    3.278004e-19, 3.281909e-19, 3.280725e-19, 3.281924e-19, 3.275913e-19, 
    3.278489e-19, 3.273199e-19, 3.252566e-19, 3.258633e-19, 3.240527e-19, 
    3.229622e-19, 3.222381e-19, 3.217238e-19, 3.217965e-19, 3.21935e-19, 
    3.226473e-19, 3.233168e-19, 3.238266e-19, 3.241675e-19, 3.245033e-19, 
    3.255183e-19, 3.260559e-19, 3.272581e-19, 3.270415e-19, 3.274086e-19, 
    3.277596e-19, 3.283482e-19, 3.282514e-19, 3.285105e-19, 3.273991e-19, 
    3.281378e-19, 3.269181e-19, 3.272518e-19, 3.245935e-19, 3.235805e-19, 
    3.231487e-19, 3.227715e-19, 3.218524e-19, 3.224871e-19, 3.222369e-19, 
    3.228323e-19, 3.232103e-19, 3.230234e-19, 3.241768e-19, 3.237285e-19, 
    3.260878e-19, 3.250722e-19, 3.277186e-19, 3.27086e-19, 3.278703e-19, 
    3.274702e-19, 3.281555e-19, 3.275388e-19, 3.286071e-19, 3.288394e-19, 
    3.286806e-19, 3.292909e-19, 3.275045e-19, 3.281908e-19, 3.230181e-19, 
    3.230486e-19, 3.231907e-19, 3.225659e-19, 3.225277e-19, 3.219552e-19, 
    3.224647e-19, 3.226816e-19, 3.232323e-19, 3.235577e-19, 3.238671e-19, 
    3.245469e-19, 3.253055e-19, 3.263658e-19, 3.27127e-19, 3.276369e-19, 
    3.273244e-19, 3.276003e-19, 3.272918e-19, 3.271472e-19, 3.287523e-19, 
    3.278512e-19, 3.292031e-19, 3.291284e-19, 3.285167e-19, 3.291368e-19, 
    3.2307e-19, 3.228946e-19, 3.22285e-19, 3.227621e-19, 3.218928e-19, 
    3.223793e-19, 3.226589e-19, 3.237376e-19, 3.239747e-19, 3.241943e-19, 
    3.246279e-19, 3.251841e-19, 3.261589e-19, 3.270066e-19, 3.2778e-19, 
    3.277234e-19, 3.277433e-19, 3.279159e-19, 3.274882e-19, 3.279861e-19, 
    3.280696e-19, 3.278513e-19, 3.291184e-19, 3.287565e-19, 3.291268e-19, 
    3.288913e-19, 3.229516e-19, 3.232468e-19, 3.230873e-19, 3.233872e-19, 
    3.231758e-19, 3.241151e-19, 3.243965e-19, 3.257128e-19, 3.25173e-19, 
    3.260323e-19, 3.252604e-19, 3.253972e-19, 3.260598e-19, 3.253022e-19, 
    3.269597e-19, 3.258359e-19, 3.279226e-19, 3.268009e-19, 3.279929e-19, 
    3.277767e-19, 3.281347e-19, 3.284551e-19, 3.288582e-19, 3.296013e-19, 
    3.294293e-19, 3.300506e-19, 3.236869e-19, 3.240694e-19, 3.240359e-19, 
    3.244363e-19, 3.247322e-19, 3.253736e-19, 3.264014e-19, 3.260151e-19, 
    3.267244e-19, 3.268666e-19, 3.257891e-19, 3.264507e-19, 3.243255e-19, 
    3.246689e-19, 3.244646e-19, 3.23717e-19, 3.261038e-19, 3.248794e-19, 
    3.271395e-19, 3.264771e-19, 3.284094e-19, 3.274486e-19, 3.293346e-19, 
    3.301392e-19, 3.308969e-19, 3.317803e-19, 3.242783e-19, 3.240185e-19, 
    3.244839e-19, 3.251272e-19, 3.257244e-19, 3.265174e-19, 3.265987e-19, 
    3.267471e-19, 3.271318e-19, 3.274549e-19, 3.267938e-19, 3.27536e-19, 
    3.247481e-19, 3.262102e-19, 3.2392e-19, 3.246098e-19, 3.250894e-19, 
    3.248793e-19, 3.25971e-19, 3.262281e-19, 3.27272e-19, 3.267326e-19, 
    3.299405e-19, 3.285225e-19, 3.324532e-19, 3.313562e-19, 3.239276e-19, 
    3.242775e-19, 3.254944e-19, 3.249156e-19, 3.265705e-19, 3.269773e-19, 
    3.273082e-19, 3.277306e-19, 3.277763e-19, 3.280265e-19, 3.276165e-19, 
    3.280104e-19, 3.265191e-19, 3.271858e-19, 3.253556e-19, 3.258012e-19, 
    3.255963e-19, 3.253713e-19, 3.260655e-19, 3.268042e-19, 3.268203e-19, 
    3.27057e-19, 3.277231e-19, 3.265772e-19, 3.301228e-19, 3.27934e-19, 
    3.24659e-19, 3.253321e-19, 3.254286e-19, 3.251679e-19, 3.269365e-19, 
    3.26296e-19, 3.280205e-19, 3.275547e-19, 3.283178e-19, 3.279386e-19, 
    3.278829e-19, 3.273958e-19, 3.270923e-19, 3.263253e-19, 3.257009e-19, 
    3.252057e-19, 3.253209e-19, 3.258648e-19, 3.268494e-19, 3.277803e-19, 
    3.275764e-19, 3.282598e-19, 3.264506e-19, 3.272094e-19, 3.269161e-19, 
    3.276809e-19, 3.260048e-19, 3.274312e-19, 3.256397e-19, 3.25797e-19, 
    3.262833e-19, 3.272606e-19, 3.274773e-19, 3.277079e-19, 3.275657e-19, 
    3.268745e-19, 3.267614e-19, 3.262715e-19, 3.261361e-19, 3.257628e-19, 
    3.254534e-19, 3.25736e-19, 3.260326e-19, 3.268749e-19, 3.276333e-19, 
    3.284596e-19, 3.286618e-19, 3.296254e-19, 3.288406e-19, 3.301349e-19, 
    3.29034e-19, 3.309393e-19, 3.275143e-19, 3.290022e-19, 3.263055e-19, 
    3.265964e-19, 3.271221e-19, 3.283275e-19, 3.276773e-19, 3.284378e-19, 
    3.267569e-19, 3.258834e-19, 3.256577e-19, 3.252358e-19, 3.256673e-19, 
    3.256323e-19, 3.260451e-19, 3.259124e-19, 3.269029e-19, 3.26371e-19, 
    3.278814e-19, 3.284319e-19, 3.299854e-19, 3.309364e-19, 3.319039e-19, 
    3.323306e-19, 3.324604e-19, 3.325147e-19 ;

 CWDN_vr =
  1.02207e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.02207e-07, 1.02207e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.02207e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.484155e-43, 0, 1.912772e-42, 
    3.629363e-43, 4.945042e-41, 1.242251e-41, 5.060599e-39, 9.290469e-41, 
    9.736725e-38, 1.98011e-39, 3.686572e-39, 8.117582e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.165713e-44, 2.802597e-45, 1.31652e-41, 
    1.734807e-42, 1.19825e-41, 6.695404e-42, 1.207219e-41, 6.067622e-43, 
    2.209848e-42, 1.527415e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.107026e-43, 3.643376e-44, 2.39622e-43, 1.41391e-42, 2.581612e-41, 
    1.610512e-41, 5.664469e-41, 2.284116e-43, 9.242965e-42, 1.961818e-44, 
    1.079e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.151867e-42, 
    4.624285e-44, 2.457878e-42, 3.279038e-43, 1.007954e-41, 4.652311e-43, 
    9.005024e-41, 2.726717e-40, 1.280843e-40, 2.25279e-39, 3.909623e-43, 
    1.19839e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    5.605194e-44, 7.637077e-43, 1.555441e-43, 6.347882e-43, 1.317221e-43, 
    6.305843e-44, 1.803401e-40, 2.237874e-42, 1.5001e-39, 1.059208e-39, 
    5.835567e-41, 1.101639e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.082857e-44, 1.566652e-42, 1.178492e-42, 1.303208e-42, 3.085659e-42, 
    3.601337e-43, 4.37065e-42, 6.605721e-42, 2.235071e-42, 1.01087e-39, 
    1.837845e-40, 1.051384e-39, 3.479578e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.382207e-44, 0, 3.190757e-42, 9.809089e-45, 4.519188e-42, 
    1.540027e-42, 9.090223e-42, 4.333936e-41, 2.977451e-40, 9.368527e-39, 
    4.266976e-39, 7.056501e-38, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 
    7.006492e-45, 1.401298e-44, 0, 1.401298e-45, 0, 0, 0, 0, 0, 0, 
    6.025583e-44, 1.401298e-45, 3.474379e-41, 2.942727e-43, 2.759103e-39, 
    1.047586e-37, 2.781373e-36, 1.085173e-34, 0, 0, 0, 0, 0, 2.802597e-45, 
    4.203895e-45, 8.407791e-45, 5.745324e-44, 3.040818e-43, 9.809089e-45, 
    4.582246e-43, 0, 0, 0, 0, 0, 0, 0, 0, 1.191104e-43, 7.006492e-45, 
    4.333622e-38, 6.009609e-41, 1.567935e-33, 1.911503e-35, 0, 0, 0, 0, 
    2.802597e-45, 2.662467e-44, 1.429324e-43, 1.223334e-42, 1.537224e-42, 
    5.338947e-42, 6.880375e-43, 4.926965e-42, 2.802597e-45, 7.707142e-44, 0, 
    0, 0, 0, 0, 9.809089e-45, 1.121039e-44, 3.923636e-44, 1.1869e-42, 
    2.802597e-45, 9.780159e-38, 3.396747e-42, 0, 0, 0, 0, 2.101948e-44, 0, 
    5.179199e-42, 5.044674e-43, 2.225822e-41, 3.454201e-42, 2.617626e-42, 
    2.242078e-43, 4.764415e-44, 1.401298e-45, 0, 0, 0, 0, 1.261169e-44, 
    1.569454e-42, 5.63322e-43, 1.677915e-41, 1.401298e-45, 8.68805e-44, 
    1.821688e-44, 9.52883e-43, 0, 2.704506e-43, 0, 0, 0, 1.121039e-43, 
    3.405155e-43, 1.091612e-42, 5.324934e-43, 1.541428e-44, 8.407791e-45, 0, 
    0, 0, 0, 0, 0, 1.541428e-44, 7.496947e-43, 4.430766e-41, 1.170028e-40, 
    1.048755e-38, 2.749264e-40, 1.032221e-37, 6.868086e-40, 3.346619e-36, 
    4.119817e-43, 5.894758e-40, 1.401298e-45, 2.802597e-45, 5.465064e-44, 
    2.339888e-41, 9.360674e-43, 3.99356e-41, 8.407791e-45, 0, 0, 0, 0, 0, 0, 
    0, 1.821688e-44, 1.401298e-45, 2.599409e-42, 3.878654e-41, 5.282891e-38, 
    3.295288e-36, 1.781647e-34, 9.699692e-34, 1.611632e-33, 1.990581e-33 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  23.61273, 23.67458, 23.66257, 23.71245, 23.68481, 23.71745, 23.6253, 
    23.677, 23.64402, 23.61835, 23.80925, 23.71469, 23.90811, 23.84758, 
    23.99988, 23.89862, 24.02034, 23.99706, 24.06741, 24.04725, 24.13711, 
    24.07672, 24.18391, 24.12274, 24.13227, 24.07471, 23.7338, 23.79743, 
    23.73001, 23.73908, 23.73503, 23.68535, 23.66026, 23.60807, 23.61756, 
    23.65593, 23.74316, 23.7136, 23.78833, 23.78665, 23.86992, 23.83236, 
    23.97259, 23.93272, 24.0481, 24.01904, 24.04671, 24.03834, 24.04682, 
    24.00422, 24.02247, 23.98503, 23.83937, 23.8821, 23.7547, 23.67812, 
    23.62755, 23.59163, 23.5967, 23.60636, 23.65616, 23.7031, 23.73887, 
    23.7628, 23.7864, 23.85766, 23.89564, 23.9806, 23.96535, 23.99126, 
    24.01616, 24.05786, 24.05101, 24.06936, 23.99064, 24.04292, 23.95664, 
    23.98021, 23.79248, 23.72159, 23.6912, 23.66487, 23.6006, 23.64495, 
    23.62746, 23.66917, 23.69564, 23.68256, 23.76345, 23.73198, 23.89789, 
    23.82636, 24.01325, 23.96848, 24.024, 23.99568, 24.04419, 24.00053, 
    24.07623, 24.09268, 24.08143, 24.12479, 23.9981, 24.04668, 23.68217, 
    23.68431, 23.69427, 23.65046, 23.6478, 23.60779, 23.64342, 23.65858, 
    23.6972, 23.71999, 23.74169, 23.78944, 23.84278, 23.91755, 23.97138, 
    24.00748, 23.98537, 24.00489, 23.98305, 23.97284, 24.08649, 24.02262, 
    24.11855, 24.11325, 24.06979, 24.11385, 23.68581, 23.67353, 23.63084, 
    23.66425, 23.60344, 23.63743, 23.65696, 23.73256, 23.74927, 23.76466, 
    23.79515, 23.83427, 23.90296, 23.96284, 24.01762, 24.01361, 24.01502, 
    24.02723, 23.99694, 24.0322, 24.03809, 24.02265, 24.11254, 24.08685, 
    24.11314, 24.09642, 23.67753, 23.6982, 23.68703, 23.70802, 23.6932, 
    23.75904, 23.77879, 23.87145, 23.83348, 23.89401, 23.83966, 23.84926, 
    23.89584, 23.84262, 23.95947, 23.88009, 24.0277, 23.94819, 24.03268, 
    24.01738, 24.04275, 24.06544, 24.09406, 24.14681, 24.1346, 24.1788, 
    23.72906, 23.75587, 23.75357, 23.78168, 23.80247, 23.84764, 23.92009, 
    23.89286, 23.94294, 23.95298, 23.87693, 23.92355, 23.77386, 23.79795, 
    23.78365, 23.73114, 23.89904, 23.81276, 23.97226, 23.92545, 24.06219, 
    23.99408, 24.12787, 24.18499, 24.23911, 24.30205, 23.77057, 23.75234, 
    23.78504, 23.83021, 23.87234, 23.92829, 23.93406, 23.94453, 23.97174, 
    23.9946, 23.94778, 24.00034, 23.80341, 23.90657, 23.74539, 23.79378, 
    23.82757, 23.81281, 23.88976, 23.90789, 23.9816, 23.94352, 24.17083, 
    24.07014, 24.35025, 24.27179, 23.74596, 23.77054, 23.85609, 23.81538, 
    23.93206, 23.9608, 23.98422, 24.01407, 24.01735, 24.03505, 24.00603, 
    24.03393, 23.92841, 23.97555, 23.84638, 23.87775, 23.86334, 23.84749, 
    23.89642, 23.9485, 23.94971, 23.9664, 24.01328, 23.93254, 24.18365, 
    24.02826, 23.79735, 23.84462, 23.8515, 23.83316, 23.95791, 23.91266, 
    24.03464, 24.00167, 24.05572, 24.02884, 24.02489, 23.99041, 23.96893, 
    23.91472, 23.87067, 23.83583, 23.84394, 23.88223, 23.95171, 24.0176, 
    24.00314, 24.05161, 23.92359, 23.97718, 23.95643, 24.01058, 23.89211, 
    23.99266, 23.8664, 23.87748, 23.91177, 23.98075, 23.99618, 24.01247, 
    24.00244, 23.95349, 23.94552, 23.91096, 23.90137, 23.87508, 23.85328, 
    23.87317, 23.89405, 23.95356, 24.00718, 24.06575, 24.08013, 24.14838, 
    24.09267, 24.18449, 24.1062, 24.24191, 23.99865, 24.10411, 23.91336, 
    23.9339, 23.97097, 24.0563, 24.01033, 24.06415, 23.94522, 23.88349, 
    23.86766, 23.83793, 23.86834, 23.86587, 23.89499, 23.88564, 23.95553, 
    23.91798, 24.02476, 24.06375, 24.17413, 24.24183, 24.311, 24.34151, 
    24.35081, 24.35468 ;

 EFLX_LH_TOT_R =
  23.61273, 23.67458, 23.66257, 23.71245, 23.68481, 23.71745, 23.6253, 
    23.677, 23.64402, 23.61835, 23.80925, 23.71469, 23.90811, 23.84758, 
    23.99988, 23.89862, 24.02034, 23.99706, 24.06741, 24.04725, 24.13711, 
    24.07672, 24.18391, 24.12274, 24.13227, 24.07471, 23.7338, 23.79743, 
    23.73001, 23.73908, 23.73503, 23.68535, 23.66026, 23.60807, 23.61756, 
    23.65593, 23.74316, 23.7136, 23.78833, 23.78665, 23.86992, 23.83236, 
    23.97259, 23.93272, 24.0481, 24.01904, 24.04671, 24.03834, 24.04682, 
    24.00422, 24.02247, 23.98503, 23.83937, 23.8821, 23.7547, 23.67812, 
    23.62755, 23.59163, 23.5967, 23.60636, 23.65616, 23.7031, 23.73887, 
    23.7628, 23.7864, 23.85766, 23.89564, 23.9806, 23.96535, 23.99126, 
    24.01616, 24.05786, 24.05101, 24.06936, 23.99064, 24.04292, 23.95664, 
    23.98021, 23.79248, 23.72159, 23.6912, 23.66487, 23.6006, 23.64495, 
    23.62746, 23.66917, 23.69564, 23.68256, 23.76345, 23.73198, 23.89789, 
    23.82636, 24.01325, 23.96848, 24.024, 23.99568, 24.04419, 24.00053, 
    24.07623, 24.09268, 24.08143, 24.12479, 23.9981, 24.04668, 23.68217, 
    23.68431, 23.69427, 23.65046, 23.6478, 23.60779, 23.64342, 23.65858, 
    23.6972, 23.71999, 23.74169, 23.78944, 23.84278, 23.91755, 23.97138, 
    24.00748, 23.98537, 24.00489, 23.98305, 23.97284, 24.08649, 24.02262, 
    24.11855, 24.11325, 24.06979, 24.11385, 23.68581, 23.67353, 23.63084, 
    23.66425, 23.60344, 23.63743, 23.65696, 23.73256, 23.74927, 23.76466, 
    23.79515, 23.83427, 23.90296, 23.96284, 24.01762, 24.01361, 24.01502, 
    24.02723, 23.99694, 24.0322, 24.03809, 24.02265, 24.11254, 24.08685, 
    24.11314, 24.09642, 23.67753, 23.6982, 23.68703, 23.70802, 23.6932, 
    23.75904, 23.77879, 23.87145, 23.83348, 23.89401, 23.83966, 23.84926, 
    23.89584, 23.84262, 23.95947, 23.88009, 24.0277, 23.94819, 24.03268, 
    24.01738, 24.04275, 24.06544, 24.09406, 24.14681, 24.1346, 24.1788, 
    23.72906, 23.75587, 23.75357, 23.78168, 23.80247, 23.84764, 23.92009, 
    23.89286, 23.94294, 23.95298, 23.87693, 23.92355, 23.77386, 23.79795, 
    23.78365, 23.73114, 23.89904, 23.81276, 23.97226, 23.92545, 24.06219, 
    23.99408, 24.12787, 24.18499, 24.23911, 24.30205, 23.77057, 23.75234, 
    23.78504, 23.83021, 23.87234, 23.92829, 23.93406, 23.94453, 23.97174, 
    23.9946, 23.94778, 24.00034, 23.80341, 23.90657, 23.74539, 23.79378, 
    23.82757, 23.81281, 23.88976, 23.90789, 23.9816, 23.94352, 24.17083, 
    24.07014, 24.35025, 24.27179, 23.74596, 23.77054, 23.85609, 23.81538, 
    23.93206, 23.9608, 23.98422, 24.01407, 24.01735, 24.03505, 24.00603, 
    24.03393, 23.92841, 23.97555, 23.84638, 23.87775, 23.86334, 23.84749, 
    23.89642, 23.9485, 23.94971, 23.9664, 24.01328, 23.93254, 24.18365, 
    24.02826, 23.79735, 23.84462, 23.8515, 23.83316, 23.95791, 23.91266, 
    24.03464, 24.00167, 24.05572, 24.02884, 24.02489, 23.99041, 23.96893, 
    23.91472, 23.87067, 23.83583, 23.84394, 23.88223, 23.95171, 24.0176, 
    24.00314, 24.05161, 23.92359, 23.97718, 23.95643, 24.01058, 23.89211, 
    23.99266, 23.8664, 23.87748, 23.91177, 23.98075, 23.99618, 24.01247, 
    24.00244, 23.95349, 23.94552, 23.91096, 23.90137, 23.87508, 23.85328, 
    23.87317, 23.89405, 23.95356, 24.00718, 24.06575, 24.08013, 24.14838, 
    24.09267, 24.18449, 24.1062, 24.24191, 23.99865, 24.10411, 23.91336, 
    23.9339, 23.97097, 24.0563, 24.01033, 24.06415, 23.94522, 23.88349, 
    23.86766, 23.83793, 23.86834, 23.86587, 23.89499, 23.88564, 23.95553, 
    23.91798, 24.02476, 24.06375, 24.17413, 24.24183, 24.311, 24.34151, 
    24.35081, 24.35468 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.191079e-08, 6.218382e-08, 6.213074e-08, 6.235096e-08, 6.22288e-08, 
    6.2373e-08, 6.196615e-08, 6.219464e-08, 6.204878e-08, 6.193537e-08, 
    6.277832e-08, 6.236078e-08, 6.321213e-08, 6.294581e-08, 6.361488e-08, 
    6.317068e-08, 6.370446e-08, 6.360209e-08, 6.391026e-08, 6.382197e-08, 
    6.421612e-08, 6.395101e-08, 6.442048e-08, 6.415281e-08, 6.419468e-08, 
    6.394226e-08, 6.244482e-08, 6.272633e-08, 6.242814e-08, 6.246828e-08, 
    6.245027e-08, 6.223132e-08, 6.212098e-08, 6.188993e-08, 6.193188e-08, 
    6.210158e-08, 6.248633e-08, 6.235573e-08, 6.268491e-08, 6.267748e-08, 
    6.304396e-08, 6.287872e-08, 6.349475e-08, 6.331966e-08, 6.382565e-08, 
    6.369839e-08, 6.381968e-08, 6.378291e-08, 6.382015e-08, 6.363351e-08, 
    6.371348e-08, 6.354926e-08, 6.290966e-08, 6.309762e-08, 6.253705e-08, 
    6.219999e-08, 6.197617e-08, 6.181733e-08, 6.183978e-08, 6.188259e-08, 
    6.210257e-08, 6.230942e-08, 6.246706e-08, 6.25725e-08, 6.267641e-08, 
    6.299089e-08, 6.315737e-08, 6.353015e-08, 6.346289e-08, 6.357685e-08, 
    6.368574e-08, 6.386854e-08, 6.383846e-08, 6.391899e-08, 6.357385e-08, 
    6.380323e-08, 6.342457e-08, 6.352813e-08, 6.270461e-08, 6.239097e-08, 
    6.225762e-08, 6.214094e-08, 6.185705e-08, 6.20531e-08, 6.197581e-08, 
    6.215969e-08, 6.227652e-08, 6.221874e-08, 6.257539e-08, 6.243673e-08, 
    6.316724e-08, 6.285257e-08, 6.367303e-08, 6.34767e-08, 6.37201e-08, 
    6.35959e-08, 6.380871e-08, 6.361718e-08, 6.394897e-08, 6.402121e-08, 
    6.397185e-08, 6.416151e-08, 6.360656e-08, 6.381967e-08, 6.221712e-08, 
    6.222654e-08, 6.227045e-08, 6.207744e-08, 6.206563e-08, 6.188878e-08, 
    6.204615e-08, 6.211316e-08, 6.22833e-08, 6.238393e-08, 6.247959e-08, 
    6.268994e-08, 6.292485e-08, 6.325337e-08, 6.348942e-08, 6.364765e-08, 
    6.355063e-08, 6.363629e-08, 6.354053e-08, 6.349565e-08, 6.399414e-08, 
    6.371423e-08, 6.413423e-08, 6.411099e-08, 6.392091e-08, 6.411361e-08, 
    6.223316e-08, 6.217893e-08, 6.199063e-08, 6.213799e-08, 6.186952e-08, 
    6.201979e-08, 6.210619e-08, 6.243962e-08, 6.251289e-08, 6.258082e-08, 
    6.271499e-08, 6.288717e-08, 6.318925e-08, 6.34521e-08, 6.369208e-08, 
    6.367449e-08, 6.368068e-08, 6.373428e-08, 6.36015e-08, 6.375608e-08, 
    6.378202e-08, 6.37142e-08, 6.410788e-08, 6.39954e-08, 6.411049e-08, 
    6.403727e-08, 6.219656e-08, 6.228781e-08, 6.22385e-08, 6.233122e-08, 
    6.22659e-08, 6.255637e-08, 6.264347e-08, 6.305104e-08, 6.288379e-08, 
    6.315e-08, 6.291083e-08, 6.295321e-08, 6.315866e-08, 6.292376e-08, 
    6.34376e-08, 6.30892e-08, 6.373637e-08, 6.338842e-08, 6.375817e-08, 
    6.369104e-08, 6.38022e-08, 6.390175e-08, 6.402701e-08, 6.425812e-08, 
    6.420461e-08, 6.43979e-08, 6.242386e-08, 6.254222e-08, 6.253181e-08, 
    6.265568e-08, 6.27473e-08, 6.294588e-08, 6.326439e-08, 6.314462e-08, 
    6.336451e-08, 6.340865e-08, 6.307459e-08, 6.327969e-08, 6.262145e-08, 
    6.272778e-08, 6.266447e-08, 6.243319e-08, 6.31722e-08, 6.279292e-08, 
    6.349332e-08, 6.328784e-08, 6.388755e-08, 6.358929e-08, 6.417515e-08, 
    6.442559e-08, 6.466136e-08, 6.493683e-08, 6.260683e-08, 6.25264e-08, 
    6.267042e-08, 6.286966e-08, 6.305456e-08, 6.330037e-08, 6.332552e-08, 
    6.337157e-08, 6.349087e-08, 6.359117e-08, 6.338612e-08, 6.361631e-08, 
    6.275242e-08, 6.320513e-08, 6.249599e-08, 6.27095e-08, 6.285792e-08, 
    6.279282e-08, 6.313093e-08, 6.321061e-08, 6.353445e-08, 6.336705e-08, 
    6.436377e-08, 6.392277e-08, 6.514664e-08, 6.480458e-08, 6.24983e-08, 
    6.260656e-08, 6.298333e-08, 6.280406e-08, 6.331678e-08, 6.3443e-08, 
    6.354561e-08, 6.367676e-08, 6.369093e-08, 6.376864e-08, 6.364129e-08, 
    6.376361e-08, 6.33009e-08, 6.350767e-08, 6.294027e-08, 6.307836e-08, 
    6.301484e-08, 6.294515e-08, 6.316022e-08, 6.338935e-08, 6.339426e-08, 
    6.346773e-08, 6.367474e-08, 6.331886e-08, 6.442066e-08, 6.374017e-08, 
    6.272461e-08, 6.293312e-08, 6.296292e-08, 6.288214e-08, 6.343034e-08, 
    6.32317e-08, 6.376674e-08, 6.362214e-08, 6.385908e-08, 6.374134e-08, 
    6.372401e-08, 6.35728e-08, 6.347865e-08, 6.32408e-08, 6.30473e-08, 
    6.289386e-08, 6.292954e-08, 6.309808e-08, 6.340337e-08, 6.36922e-08, 
    6.362893e-08, 6.384107e-08, 6.327961e-08, 6.351502e-08, 6.342403e-08, 
    6.36613e-08, 6.314143e-08, 6.358408e-08, 6.302828e-08, 6.307702e-08, 
    6.322776e-08, 6.353098e-08, 6.359809e-08, 6.366972e-08, 6.362552e-08, 
    6.341112e-08, 6.337601e-08, 6.322409e-08, 6.318215e-08, 6.306641e-08, 
    6.297058e-08, 6.305813e-08, 6.315008e-08, 6.341122e-08, 6.364657e-08, 
    6.390317e-08, 6.396598e-08, 6.426577e-08, 6.402171e-08, 6.442445e-08, 
    6.408201e-08, 6.467483e-08, 6.360975e-08, 6.407196e-08, 6.323462e-08, 
    6.332483e-08, 6.348797e-08, 6.386221e-08, 6.366019e-08, 6.389647e-08, 
    6.337463e-08, 6.310389e-08, 6.303387e-08, 6.290318e-08, 6.303685e-08, 
    6.302598e-08, 6.315389e-08, 6.311279e-08, 6.341989e-08, 6.325493e-08, 
    6.372358e-08, 6.38946e-08, 6.437764e-08, 6.467376e-08, 6.497525e-08, 
    6.510835e-08, 6.514885e-08, 6.516579e-08 ;

 ERRH2O =
  -22917.11, -22951.63, -22944.87, -22973.11, -22957.39, -22975.96, 
    -22924.05, -22953.02, -22934.47, -22920.19, -23029.13, -22974.38, 
    -23087.75, -23051.51, -23143.27, -23082.06, -23155.84, -23141.47, 
    -23185.1, -23172.48, -23229.54, -23190.95, -23259.93, -23220.24, 
    -23226.38, -23189.7, -22985.28, -23022.25, -22983.11, -22988.34, 
    -22985.99, -22957.71, -22943.63, -22914.49, -22919.75, -22941.16, 
    -22990.69, -22973.72, -23016.76, -23015.78, -23064.77, -23042.5, 
    -23126.55, -23102.5, -23173.01, -23154.98, -23172.16, -23166.93, 
    -23172.23, -23145.87, -23157.11, -23134.11, -23046.65, -23072.07, 
    -22997.33, -22953.71, -22925.31, -22905.41, -22908.21, -22913.57, 
    -22941.29, -22967.74, -22988.17, -23001.98, -23015.64, -23057.6, 
    -23080.23, -23131.46, -23122.14, -23137.96, -23153.2, -23179.13, 
    -23174.83, -23186.36, -23137.53, -23169.82, -23116.86, -23131.18, 
    -23019.38, -22978.28, -22961.09, -22946.16, -22910.37, -22935.02, 
    -22925.27, -22948.55, -22963.51, -22956.1, -23002.36, -22984.22, 
    -23081.59, -23039.01, -23151.41, -23124.05, -23158.04, -23140.61, 
    -23170.6, -23143.58, -23190.66, -23201.09, -23193.96, -23221.51, 
    -23142.1, -23172.16, -22955.89, -22957.1, -22962.73, -22938.1, -22936.6, 
    -22914.34, -22934.14, -22942.63, -22964.38, -22977.37, -22989.81, 
    -23017.42, -23048.69, -23093.43, -23125.81, -23147.85, -23134.3, 
    -23146.26, -23132.9, -23126.67, -23197.18, -23157.21, -23217.52, 
    -23214.12, -23186.63, -23214.5, -22957.95, -22951, -22927.13, -22945.79, 
    -22911.93, -22930.81, -22941.75, -22984.61, -22994.16, -23003.07, 
    -23020.73, -23043.63, -23084.6, -23120.66, -23154.09, -23151.62, 
    -23152.49, -23160.05, -23141.39, -23163.13, -23166.81, -23157.21, 
    -23213.67, -23197.35, -23214.05, -23203.4, -22953.26, -22964.96, 
    -22958.63, -22970.56, -22962.15, -22999.87, -23011.32, -23065.74, 
    -23043.18, -23079.22, -23046.81, -23052.5, -23080.42, -23048.54, 
    -23118.66, -23070.93, -23160.34, -23111.91, -23163.43, -23153.95, 
    -23169.67, -23183.88, -23201.92, -23235.73, -23227.84, -23256.54, 
    -22982.55, -22998.01, -22996.64, -23012.91, -23025.01, -23051.52, 
    -23094.95, -23078.48, -23108.62, -23114.68, -23068.93, -23097.06, 
    -23008.42, -23022.43, -23014.07, -22983.77, -23082.27, -23031.06, 
    -23126.35, -23098.16, -23181.85, -23139.69, -23223.51, -23260.7, 
    -23296.52, -23339.05, -23006.5, -22995.93, -23014.85, -23041.29, 
    -23066.21, -23099.87, -23103.3, -23109.59, -23126.01, -23139.95, 
    -23111.59, -23143.46, -23025.7, -23086.79, -22991.95, -23020.01, 
    -23039.72, -23031.04, -23076.61, -23087.54, -23132.05, -23108.97, 
    -23251.44, -23186.9, -23371.76, -23318.66, -22992.25, -23006.46, 
    -23056.57, -23032.54, -23102.1, -23119.4, -23133.6, -23151.94, -23153.93, 
    -23164.91, -23146.96, -23164.2, -23099.94, -23128.34, -23050.76, 
    -23069.44, -23060.82, -23051.42, -23080.62, -23112.03, -23112.7, 
    -23122.82, -23151.68, -23102.39, -23259.97, -23160.9, -23022, -23049.81, 
    -23053.81, -23042.96, -23117.66, -23090.44, -23164.64, -23144.28, 
    -23177.78, -23161.04, -23158.6, -23137.38, -23124.32, -23091.7, 
    -23065.22, -23044.53, -23049.32, -23072.13, -23113.96, -23154.11, 
    -23145.23, -23175.21, -23097.04, -23129.36, -23116.79, -23149.77, 
    -23078.05, -23138.98, -23062.64, -23069.26, -23089.9, -23131.58, 
    -23140.91, -23150.95, -23144.75, -23115.02, -23110.2, -23089.39, 
    -23083.62, -23067.81, -23054.84, -23066.69, -23079.23, -23115.03, 
    -23147.7, -23184.09, -23193.11, -23236.88, -23201.17, -23260.54, 
    -23209.93, -23298.61, -23142.55, -23208.46, -23090.84, -23103.2, 
    -23125.62, -23178.23, -23149.61, -23183.13, -23110.01, -23072.93, 
    -23063.4, -23045.78, -23063.8, -23062.33, -23079.75, -23074.13, 
    -23116.22, -23093.64, -23158.54, -23182.87, -23253.5, -23298.43, -23345, 
    -23365.74, -23372.1, -23374.77 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -1.391141e-14, -1.570146e-14, -1.126283e-14, -7.917224e-15, -1.209914e-14, 
    -2.302252e-14, -6.177798e-15, -5.781344e-15, -1.630007e-14, 
    -2.495912e-14, -1.553075e-14, -6.488593e-15, -1.390573e-14, 
    -9.813985e-15, -1.421952e-14, -1.179e-14, -1.146756e-14, -6.143575e-15, 
    -1.265104e-14, -9.648389e-15, -1.656536e-14, -3.539731e-15, 
    -1.042794e-14, -1.439804e-14, -6.364243e-15, -3.247922e-15, 
    -1.374868e-14, -1.802247e-14, -1.199577e-14, -7.572756e-15, 
    -1.668098e-14, -1.436094e-14, -1.643472e-14, -1.981884e-14, 
    -1.620193e-14, -1.167657e-14, -7.357919e-15, -1.199333e-14, 
    -1.532354e-14, -6.912196e-15, -1.919204e-14, -1.926221e-14, 
    -1.150654e-14, -1.648021e-14, -1.058201e-14, -1.396022e-14, 
    -1.711105e-14, -1.232407e-14, -1.982997e-14, -9.78941e-15, -1.635528e-14, 
    -1.397102e-14, -1.158874e-14, -2.231852e-14, -1.619222e-14, 
    -2.958253e-15, -1.719422e-14, -1.19095e-14, -4.90194e-15, -1.542257e-14, 
    -5.674319e-15, -1.169466e-14, -1.079505e-14, -2.280947e-14, 
    -1.116903e-14, -1.212656e-14, -1.473404e-14, -5.009407e-15, 
    -1.095218e-14, -7.127751e-15, -1.476591e-14, -1.855698e-14, 
    -1.835963e-14, -1.095022e-14, -1.359158e-14, -1.506284e-14, 
    -1.757226e-16, -1.166995e-14, -1.660382e-14, -1.720861e-14, 
    -9.145998e-15, -1.242841e-14, -1.787334e-14, -9.322959e-15, 
    -1.681737e-14, -1.080511e-14, -1.942201e-14, -1.044943e-14, 
    -1.261301e-14, -7.303438e-15, -2.091508e-14, -1.525515e-14, 
    -1.725938e-14, -1.391725e-14, -9.561551e-15, -1.236555e-14, 
    -1.668984e-14, -1.033878e-14, -8.512132e-15, -8.834637e-15, 
    -2.069017e-14, -1.007789e-14, -9.327828e-15, -2.281002e-14, 
    -7.136039e-15, -1.250046e-14, -1.429242e-14, -1.201493e-14, 
    -1.581577e-14, -1.583106e-14, -7.892564e-15, -1.9326e-14, -8.583755e-15, 
    -1.133297e-14, -1.003208e-14, -6.423033e-15, -1.35445e-14, -1.361302e-14, 
    -1.266404e-14, -7.502326e-15, -1.922084e-14, -1.713099e-14, 
    -1.173016e-14, -4.532274e-15, -1.583672e-14, -1.230282e-14, 
    -1.311597e-14, -9.888612e-15, -1.036496e-14, -1.860786e-14, 
    -1.157154e-14, -2.137996e-14, -8.990806e-15, -4.911294e-15, 
    -9.854336e-15, -1.546852e-14, -1.466978e-14, -4.775967e-15, 
    -8.724388e-15, -1.580735e-14, -1.417445e-14, -8.922649e-15, 
    -1.307352e-14, -1.085229e-14, -1.51656e-14, -1.25766e-14, -1.463963e-14, 
    -1.186027e-14, -1.169386e-14, -5.985311e-15, -1.009561e-14, 
    -9.280076e-15, -8.271661e-15, -7.250444e-15, -1.006482e-14, 
    -1.263992e-14, -8.949996e-15, -1.271004e-14, -1.126639e-14, 
    -5.605795e-15, -1.148152e-14, -1.739421e-14, -1.203436e-14, 
    -1.255543e-14, -6.369944e-15, -9.504428e-15, -1.045897e-14, 
    -1.596529e-14, -1.950206e-14, -9.116657e-15, -9.53774e-15, -2.036699e-14, 
    -1.228291e-14, -8.779698e-15, -1.13576e-14, -1.374954e-14, -1.127385e-14, 
    -1.108214e-14, -2.77596e-15, -1.216381e-14, 1.555816e-15, -2.682886e-15, 
    -6.851363e-15, -1.80659e-14, -1.776454e-14, -1.187931e-14, -1.300295e-14, 
    -1.434136e-14, -1.466526e-14, -1.655267e-14, -2.158869e-14, 
    -1.414235e-14, -1.395773e-14, -1.083398e-14, -5.961931e-15, 
    -7.385797e-15, -1.121367e-14, -1.17807e-14, -6.811303e-15, -7.630665e-15, 
    -1.420365e-14, -4.567324e-15, -1.701614e-14, -1.043011e-14, 
    -2.004829e-14, -1.312145e-14, -2.136039e-14, -1.270696e-14, 
    -1.225836e-14, -1.410178e-15, -1.122309e-14, -1.055113e-14, 
    -1.467201e-14, -1.599217e-14, -1.421476e-14, -2.155474e-14, 
    -1.569113e-14, -5.9223e-15, -6.723629e-15, -1.21631e-14, -1.636952e-14, 
    -9.150355e-15, -1.443981e-14, -2.197916e-14, -8.931236e-15, 
    -1.118278e-14, -8.178992e-15, -1.587292e-14, -1.578597e-14, 
    -5.454387e-15, -1.797317e-14, -9.242564e-15, -1.248498e-14, 
    -1.452412e-14, -1.425794e-15, 1.907699e-15, -1.361483e-14, -1.827363e-14, 
    -2.196601e-14, -8.340204e-15, -6.441043e-15, -1.420467e-14, -1.49856e-14, 
    -8.980983e-15, -1.022532e-14, -1.528606e-14, -1.788478e-14, 
    -2.019705e-14, -4.223794e-15, -1.694965e-14, -1.303448e-14, 
    -1.066416e-14, -1.107509e-14, -1.23802e-14, -2.279187e-14, -1.754138e-14, 
    -1.33459e-14, -8.854113e-15, -1.121863e-14, -2.68215e-15, -1.78619e-14, 
    -9.323921e-15, -1.2673e-14, -1.145106e-14, -3.96501e-15, -1.076243e-14, 
    -1.737066e-14, -2.058942e-14, -8.816862e-15, -1.435651e-14, 
    -8.583012e-15, -1.958154e-14, -1.771297e-14, -1.635956e-14, 
    -1.698028e-14, -1.1009e-14, -1.52984e-14, -1.682025e-14, -7.864233e-15, 
    -6.143332e-15, -1.243327e-14, -1.226269e-14, -6.429246e-15, 
    -1.546479e-14, -1.899335e-14, -1.566122e-14, -8.724141e-15, 
    -1.579585e-14, -1.478904e-14, -4.416675e-15, -6.230938e-15, 
    -7.299029e-15, -1.314764e-14, -1.232922e-14, -1.618324e-14, 
    -1.491142e-14, -1.060629e-14, -1.119616e-14, -1.83433e-14, -2.179965e-14, 
    -1.050867e-14, -1.414443e-14, -1.53393e-14, -1.273398e-14, -1.629328e-14, 
    -1.937411e-14, -4.899542e-15, -1.191187e-14, -1.584327e-14, 
    -1.301605e-14, -1.262826e-15, -8.678742e-15, -1.163093e-14, 
    -1.321058e-14, -7.754646e-15, -1.385736e-14, -9.142768e-17, 
    -1.349506e-14, -1.254895e-14, -1.924067e-14, -6.947423e-15, -6.70815e-15, 
    -2.794965e-14, -1.516536e-14, -1.021617e-14, -5.174171e-15, 
    -1.050696e-14, -6.202647e-15, -1.162474e-14, -1.873371e-14, -3.62568e-15, 
    -1.452511e-14, -1.514318e-14, -1.53087e-14, -1.367095e-14, -1.872747e-14, 
    -1.252414e-14, -5.28902e-15 ;

 ERRSOI =
  -2.679635e-10, -2.914086e-10, -3.361442e-10, -4.074025e-10, -3.561985e-10, 
    -4.10075e-10, -4.877573e-10, -2.512739e-10, -3.354465e-10, -4.597309e-10, 
    -2.077554e-10, -4.234575e-10, -4.400583e-10, -4.14928e-10, -8.925779e-11, 
    -2.622515e-10, -5.46077e-10, -3.225623e-10, -5.00241e-10, -2.862025e-10, 
    -2.757815e-10, -3.636293e-10, -4.491896e-10, -1.619652e-10, -2.41464e-10, 
    -4.364058e-10, -3.79787e-10, -2.737034e-10, -4.831806e-10, -2.473732e-10, 
    -6.680314e-10, -3.96623e-10, -3.111149e-10, -3.527134e-10, -2.275502e-10, 
    -4.238651e-10, -4.238372e-10, -4.257125e-10, -2.822862e-10, 
    -3.062466e-10, -1.493668e-10, -5.207458e-10, -2.291384e-10, 
    -3.470213e-10, -4.497254e-10, -3.89888e-10, -1.071405e-10, -3.504692e-10, 
    -1.274127e-10, -2.949308e-10, -3.286343e-10, -4.636837e-10, 
    -3.970938e-10, -3.635082e-10, -3.187569e-10, -4.519713e-10, 
    -2.602159e-10, -5.422919e-10, -2.890276e-10, -3.248208e-10, 
    -2.596713e-10, -3.304994e-10, -4.269066e-10, -3.242039e-10, 
    -3.819834e-10, -4.311789e-10, -3.224023e-10, -2.222365e-10, 
    -2.774969e-10, -3.051426e-10, -4.360152e-10, -5.054094e-10, 
    -2.951249e-10, -2.938544e-10, -1.952754e-10, -3.145183e-10, 
    -2.263311e-10, -1.752899e-10, -2.037214e-10, -5.955132e-10, 
    -4.205686e-10, -3.80871e-10, -3.808623e-10, -3.093601e-10, -3.338894e-10, 
    -3.476961e-10, -3.029003e-10, -5.838067e-10, -2.416276e-10, 
    -3.646096e-10, -3.218414e-10, -3.881331e-10, -4.318302e-10, 
    -4.040998e-10, -5.212606e-10, -3.056674e-10, -2.312184e-10, -2.27672e-10, 
    -3.727248e-10, -4.339655e-10, -2.998869e-10, -3.400986e-10, -3.11286e-10, 
    -3.923221e-10, -4.75605e-10, -4.161751e-10, -3.887031e-10, -4.07798e-10, 
    -2.092682e-10, -2.957119e-10, -3.699219e-10, -4.028385e-10, 
    -3.340543e-10, -4.327266e-10, -3.583224e-10, -4.672568e-10, 
    -1.165585e-10, -1.699862e-10, -2.331557e-10, -3.860033e-10, 
    -2.043377e-10, -3.300536e-10, -2.202532e-10, -3.759272e-10, 
    -2.630893e-10, -3.73158e-10, -2.44844e-10, -3.570985e-10, -3.285157e-10, 
    -3.727192e-10, -3.4024e-10, -1.802368e-10, -4.576224e-10, -2.851215e-10, 
    -1.846197e-10, -4.168052e-10, -4.506023e-10, -1.542811e-10, 
    -2.213304e-10, -2.695022e-10, -3.627426e-10, -3.480275e-10, 
    -4.473348e-10, -3.893925e-10, -3.169457e-10, -3.023087e-10, -3.66764e-10, 
    -2.141298e-10, -1.671617e-10, -1.672575e-10, -2.767867e-10, 
    -3.313685e-10, -3.039081e-10, -3.386581e-10, -2.180727e-10, -2.38583e-10, 
    -3.356785e-10, -3.170186e-10, -3.91183e-10, -3.496449e-10, -2.543479e-10, 
    -3.892768e-10, -4.228686e-10, -2.12153e-10, -2.488499e-10, -4.561686e-10, 
    -4.777643e-10, -4.401481e-10, -3.303394e-10, -4.476501e-10, 
    -3.568577e-10, -2.420122e-10, -4.018038e-10, -2.461547e-10, 
    -4.244326e-10, -3.208262e-10, -4.288472e-10, -3.387818e-10, -3.17869e-10, 
    -2.065804e-10, -5.2428e-10, -3.136875e-10, -4.0338e-10, -2.164403e-10, 
    -3.507523e-10, -3.136446e-10, -2.916511e-10, -1.78732e-10, -4.215365e-10, 
    -2.394427e-10, -5.425744e-10, -2.266272e-10, -3.773827e-10, 
    -4.063842e-10, -1.345799e-10, -4.080159e-10, -4.382694e-10, -3.37428e-10, 
    -5.758179e-10, -3.454529e-10, -2.863051e-10, -4.482787e-10, 
    -4.619027e-10, -1.782703e-10, -3.210581e-10, -4.031184e-10, 
    -5.546082e-10, -2.796433e-10, -3.648342e-10, -2.324861e-10, 
    -2.506498e-10, -3.138256e-10, -3.151116e-10, -1.419421e-10, 
    -5.145245e-10, -2.031632e-10, -3.693027e-10, -2.810608e-10, 
    -2.346769e-10, -1.622973e-10, -3.989336e-10, -4.232488e-10, 
    -4.357856e-10, -2.194806e-10, -3.944323e-10, -2.786974e-10, 
    -4.901172e-10, -3.910227e-10, -2.780066e-10, -2.113183e-10, 
    -2.413659e-10, -4.190494e-10, -4.130927e-10, -2.67014e-10, -3.27977e-10, 
    -2.471707e-10, -4.181598e-10, -4.440394e-10, -2.339539e-10, 
    -3.767676e-10, -2.464134e-10, -3.28604e-10, -2.451861e-10, -3.72705e-10, 
    -3.326015e-10, -3.831358e-10, -2.011471e-10, -3.258586e-10, -4.29404e-10, 
    -1.204261e-10, -3.991341e-10, -3.395152e-10, -4.551261e-10, -5.16171e-10, 
    -3.060446e-10, -4.400143e-10, -4.543085e-10, -2.656505e-10, 
    -1.582156e-10, -3.610339e-10, -2.576117e-10, -3.540091e-10, 
    -3.217533e-10, -3.979809e-10, -3.906603e-10, -4.750623e-10, 
    -1.655943e-10, -4.330003e-10, -1.927588e-10, -3.851929e-10, 
    -1.949533e-10, -2.954856e-10, -3.677322e-10, -5.310872e-10, 
    -3.583153e-10, -4.224367e-10, -3.630541e-10, -3.892885e-10, 
    -3.112057e-10, -2.45088e-10, -2.984173e-10, -4.232201e-10, -2.514166e-10, 
    -2.891791e-10, -3.120201e-10, -4.963495e-10, -3.704411e-10, 
    -2.009126e-10, -5.646567e-10, -2.129796e-10, -5.488628e-10, 
    -2.122215e-10, -2.655829e-10, -3.048611e-10, -3.999213e-10, -3.50376e-10, 
    -2.852637e-10, -4.787329e-10, -4.434904e-10, -3.191341e-10, 
    -2.851294e-10, -1.402986e-10, -4.878166e-10, -2.77126e-10, -4.051051e-10, 
    -3.13473e-10, -2.019586e-10, -1.697614e-10, -4.483171e-10, -3.044696e-10, 
    -3.825088e-10, -1.672014e-10, -2.1518e-10, -2.790084e-10, -4.145181e-10, 
    -3.399813e-10, -2.841289e-10, -3.121922e-10, -3.751709e-10, 
    -4.999566e-10, -2.140913e-10, -2.800739e-10, -2.997562e-10, 
    -4.253354e-10, -3.506783e-10, -3.473713e-10, -5.57707e-10, -3.597539e-10, 
    -2.548677e-10, -3.33828e-10, -3.061482e-10, -3.125953e-10, -4.092405e-10, 
    -4.035629e-10, -2.034844e-10, -2.411257e-10, -4.51481e-10, -3.665725e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  1.984312e-16, 1.934074e-16, 1.943843e-16, 1.903312e-16, 1.925798e-16, 
    1.899256e-16, 1.974129e-16, 1.932078e-16, 1.958925e-16, 1.979792e-16, 
    1.824624e-16, 1.901504e-16, 1.744736e-16, 1.793796e-16, 1.670525e-16, 
    1.75237e-16, 1.654016e-16, 1.67289e-16, 1.616083e-16, 1.63236e-16, 
    1.559667e-16, 1.60857e-16, 1.521973e-16, 1.571349e-16, 1.563625e-16, 
    1.610182e-16, 1.886038e-16, 1.834197e-16, 1.889109e-16, 1.881717e-16, 
    1.885035e-16, 1.925332e-16, 1.945634e-16, 1.988153e-16, 1.980435e-16, 
    1.949207e-16, 1.878394e-16, 1.902437e-16, 1.841841e-16, 1.843209e-16, 
    1.775718e-16, 1.806152e-16, 1.692671e-16, 1.724934e-16, 1.63168e-16, 
    1.655139e-16, 1.632782e-16, 1.639562e-16, 1.632694e-16, 1.667097e-16, 
    1.652357e-16, 1.682627e-16, 1.800452e-16, 1.765834e-16, 1.869059e-16, 
    1.93109e-16, 1.972285e-16, 2.001509e-16, 1.997378e-16, 1.989502e-16, 
    1.949024e-16, 1.91096e-16, 1.881946e-16, 1.862535e-16, 1.843406e-16, 
    1.785484e-16, 1.754824e-16, 1.686144e-16, 1.698544e-16, 1.677539e-16, 
    1.657472e-16, 1.623772e-16, 1.62932e-16, 1.61447e-16, 1.678095e-16, 
    1.635812e-16, 1.705606e-16, 1.686521e-16, 1.838195e-16, 1.895951e-16, 
    1.920485e-16, 1.941965e-16, 1.994201e-16, 1.958129e-16, 1.97235e-16, 
    1.938518e-16, 1.917015e-16, 1.927651e-16, 1.862004e-16, 1.887528e-16, 
    1.753006e-16, 1.810964e-16, 1.659813e-16, 1.696e-16, 1.651139e-16, 
    1.674033e-16, 1.634802e-16, 1.67011e-16, 1.608943e-16, 1.59562e-16, 
    1.604725e-16, 1.569749e-16, 1.672067e-16, 1.632781e-16, 1.927948e-16, 
    1.926214e-16, 1.918134e-16, 1.953649e-16, 1.955822e-16, 1.988364e-16, 
    1.959409e-16, 1.947077e-16, 1.91577e-16, 1.897247e-16, 1.879638e-16, 
    1.840914e-16, 1.797653e-16, 1.737141e-16, 1.693654e-16, 1.664494e-16, 
    1.682376e-16, 1.666589e-16, 1.684237e-16, 1.692508e-16, 1.600611e-16, 
    1.65222e-16, 1.57478e-16, 1.579067e-16, 1.614116e-16, 1.578584e-16, 
    1.924996e-16, 1.934977e-16, 1.969624e-16, 1.94251e-16, 1.991908e-16, 
    1.964258e-16, 1.948357e-16, 1.886993e-16, 1.87351e-16, 1.861003e-16, 
    1.836302e-16, 1.804595e-16, 1.748955e-16, 1.700529e-16, 1.656305e-16, 
    1.659546e-16, 1.658405e-16, 1.648523e-16, 1.672999e-16, 1.644504e-16, 
    1.639721e-16, 1.652227e-16, 1.579641e-16, 1.600382e-16, 1.579158e-16, 
    1.592663e-16, 1.931733e-16, 1.914938e-16, 1.924014e-16, 1.906946e-16, 
    1.91897e-16, 1.865498e-16, 1.849462e-16, 1.774409e-16, 1.805218e-16, 
    1.756185e-16, 1.800239e-16, 1.792433e-16, 1.754581e-16, 1.797859e-16, 
    1.703198e-16, 1.767378e-16, 1.648139e-16, 1.712255e-16, 1.64412e-16, 
    1.656497e-16, 1.636005e-16, 1.617649e-16, 1.594553e-16, 1.551926e-16, 
    1.561798e-16, 1.526143e-16, 1.889898e-16, 1.868106e-16, 1.870027e-16, 
    1.847221e-16, 1.830352e-16, 1.793785e-16, 1.735116e-16, 1.757181e-16, 
    1.716672e-16, 1.708537e-16, 1.770081e-16, 1.732296e-16, 1.853522e-16, 
    1.833941e-16, 1.845601e-16, 1.888178e-16, 1.752094e-16, 1.821947e-16, 
    1.692935e-16, 1.730796e-16, 1.620266e-16, 1.675245e-16, 1.567232e-16, 
    1.521025e-16, 1.47753e-16, 1.42667e-16, 1.856214e-16, 1.871022e-16, 
    1.844509e-16, 1.807816e-16, 1.773767e-16, 1.728487e-16, 1.723854e-16, 
    1.715369e-16, 1.69339e-16, 1.674905e-16, 1.712684e-16, 1.670271e-16, 
    1.829396e-16, 1.74603e-16, 1.876619e-16, 1.837305e-16, 1.80998e-16, 
    1.821969e-16, 1.759703e-16, 1.745024e-16, 1.685354e-16, 1.716204e-16, 
    1.532429e-16, 1.613768e-16, 1.387937e-16, 1.451088e-16, 1.876195e-16, 
    1.856266e-16, 1.786884e-16, 1.8199e-16, 1.725464e-16, 1.702209e-16, 
    1.683302e-16, 1.659126e-16, 1.656517e-16, 1.64219e-16, 1.665666e-16, 
    1.643118e-16, 1.72839e-16, 1.690292e-16, 1.794818e-16, 1.769383e-16, 
    1.781085e-16, 1.793919e-16, 1.754306e-16, 1.712089e-16, 1.71119e-16, 
    1.697649e-16, 1.659478e-16, 1.725082e-16, 1.521921e-16, 1.647421e-16, 
    1.834532e-16, 1.796128e-16, 1.790646e-16, 1.805524e-16, 1.704541e-16, 
    1.741138e-16, 1.64254e-16, 1.669196e-16, 1.625518e-16, 1.647224e-16, 
    1.650417e-16, 1.67829e-16, 1.695639e-16, 1.73946e-16, 1.775105e-16, 
    1.803366e-16, 1.796796e-16, 1.765749e-16, 1.709507e-16, 1.656279e-16, 
    1.66794e-16, 1.628838e-16, 1.732314e-16, 1.688934e-16, 1.705701e-16, 
    1.661976e-16, 1.757767e-16, 1.676191e-16, 1.778609e-16, 1.769633e-16, 
    1.741864e-16, 1.685989e-16, 1.673628e-16, 1.660423e-16, 1.668572e-16, 
    1.708079e-16, 1.714552e-16, 1.74254e-16, 1.750265e-16, 1.771588e-16, 
    1.789237e-16, 1.773111e-16, 1.756173e-16, 1.708064e-16, 1.664691e-16, 
    1.617387e-16, 1.605809e-16, 1.550505e-16, 1.595522e-16, 1.521222e-16, 
    1.584387e-16, 1.475027e-16, 1.671467e-16, 1.586251e-16, 1.740602e-16, 
    1.723983e-16, 1.693916e-16, 1.624933e-16, 1.662182e-16, 1.618619e-16, 
    1.714805e-16, 1.764677e-16, 1.777581e-16, 1.801648e-16, 1.777031e-16, 
    1.779033e-16, 1.755474e-16, 1.763045e-16, 1.706466e-16, 1.736861e-16, 
    1.650496e-16, 1.618964e-16, 1.529879e-16, 1.475233e-16, 1.419587e-16, 
    1.395011e-16, 1.387529e-16, 1.384402e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  23.61273, 23.67458, 23.66257, 23.71245, 23.68481, 23.71745, 23.6253, 
    23.677, 23.64402, 23.61835, 23.80925, 23.71469, 23.90811, 23.84758, 
    23.99988, 23.89862, 24.02034, 23.99706, 24.06741, 24.04725, 24.13711, 
    24.07672, 24.18391, 24.12274, 24.13227, 24.07471, 23.7338, 23.79743, 
    23.73001, 23.73908, 23.73503, 23.68535, 23.66026, 23.60807, 23.61756, 
    23.65593, 23.74316, 23.7136, 23.78833, 23.78665, 23.86992, 23.83236, 
    23.97259, 23.93272, 24.0481, 24.01904, 24.04671, 24.03834, 24.04682, 
    24.00422, 24.02247, 23.98503, 23.83937, 23.8821, 23.7547, 23.67812, 
    23.62755, 23.59163, 23.5967, 23.60636, 23.65616, 23.7031, 23.73887, 
    23.7628, 23.7864, 23.85766, 23.89564, 23.9806, 23.96535, 23.99126, 
    24.01616, 24.05786, 24.05101, 24.06936, 23.99064, 24.04292, 23.95664, 
    23.98021, 23.79248, 23.72159, 23.6912, 23.66487, 23.6006, 23.64495, 
    23.62746, 23.66917, 23.69564, 23.68256, 23.76345, 23.73198, 23.89789, 
    23.82636, 24.01325, 23.96848, 24.024, 23.99568, 24.04419, 24.00053, 
    24.07623, 24.09268, 24.08143, 24.12479, 23.9981, 24.04668, 23.68217, 
    23.68431, 23.69427, 23.65046, 23.6478, 23.60779, 23.64342, 23.65858, 
    23.6972, 23.71999, 23.74169, 23.78944, 23.84278, 23.91755, 23.97138, 
    24.00748, 23.98537, 24.00489, 23.98305, 23.97284, 24.08649, 24.02262, 
    24.11855, 24.11325, 24.06979, 24.11385, 23.68581, 23.67353, 23.63084, 
    23.66425, 23.60344, 23.63743, 23.65696, 23.73256, 23.74927, 23.76466, 
    23.79515, 23.83427, 23.90296, 23.96284, 24.01762, 24.01361, 24.01502, 
    24.02723, 23.99694, 24.0322, 24.03809, 24.02265, 24.11254, 24.08685, 
    24.11314, 24.09642, 23.67753, 23.6982, 23.68703, 23.70802, 23.6932, 
    23.75904, 23.77879, 23.87145, 23.83348, 23.89401, 23.83966, 23.84926, 
    23.89584, 23.84262, 23.95947, 23.88009, 24.0277, 23.94819, 24.03268, 
    24.01738, 24.04275, 24.06544, 24.09406, 24.14681, 24.1346, 24.1788, 
    23.72906, 23.75587, 23.75357, 23.78168, 23.80247, 23.84764, 23.92009, 
    23.89286, 23.94294, 23.95298, 23.87693, 23.92355, 23.77386, 23.79795, 
    23.78365, 23.73114, 23.89904, 23.81276, 23.97226, 23.92545, 24.06219, 
    23.99408, 24.12787, 24.18499, 24.23911, 24.30205, 23.77057, 23.75234, 
    23.78504, 23.83021, 23.87234, 23.92829, 23.93406, 23.94453, 23.97174, 
    23.9946, 23.94778, 24.00034, 23.80341, 23.90657, 23.74539, 23.79378, 
    23.82757, 23.81281, 23.88976, 23.90789, 23.9816, 23.94352, 24.17083, 
    24.07014, 24.35025, 24.27179, 23.74596, 23.77054, 23.85609, 23.81538, 
    23.93206, 23.9608, 23.98422, 24.01407, 24.01735, 24.03505, 24.00603, 
    24.03393, 23.92841, 23.97555, 23.84638, 23.87775, 23.86334, 23.84749, 
    23.89642, 23.9485, 23.94971, 23.9664, 24.01328, 23.93254, 24.18365, 
    24.02826, 23.79735, 23.84462, 23.8515, 23.83316, 23.95791, 23.91266, 
    24.03464, 24.00167, 24.05572, 24.02884, 24.02489, 23.99041, 23.96893, 
    23.91472, 23.87067, 23.83583, 23.84394, 23.88223, 23.95171, 24.0176, 
    24.00314, 24.05161, 23.92359, 23.97718, 23.95643, 24.01058, 23.89211, 
    23.99266, 23.8664, 23.87748, 23.91177, 23.98075, 23.99618, 24.01247, 
    24.00244, 23.95349, 23.94552, 23.91096, 23.90137, 23.87508, 23.85328, 
    23.87317, 23.89405, 23.95356, 24.00718, 24.06575, 24.08013, 24.14838, 
    24.09267, 24.18449, 24.1062, 24.24191, 23.99865, 24.10411, 23.91336, 
    23.9339, 23.97097, 24.0563, 24.01033, 24.06415, 23.94522, 23.88349, 
    23.86766, 23.83793, 23.86834, 23.86587, 23.89499, 23.88564, 23.95553, 
    23.91798, 24.02476, 24.06375, 24.17413, 24.24183, 24.311, 24.34151, 
    24.35081, 24.35468 ;

 FGR =
  -424.0618, -425.0807, -424.8828, -425.7042, -425.2488, -425.7865, 
    -424.2686, -425.1208, -424.577, -424.1539, -427.298, -425.7409, 
    -428.9189, -427.9251, -430.423, -428.7639, -430.7577, -430.3759, 
    -431.527, -431.1973, -432.6681, -431.6792, -433.4318, -432.4323, 
    -432.5884, -431.6465, -426.0549, -427.1039, -425.9926, -426.1422, 
    -426.0753, -425.258, -424.8456, -423.9844, -424.1409, -424.7737, 
    -426.2095, -425.7225, -426.9514, -426.9237, -428.2916, -427.6748, 
    -429.975, -429.3214, -431.211, -430.7357, -431.1886, -431.0513, 
    -431.1904, -430.4932, -430.7918, -430.1787, -427.7902, -428.4918, 
    -426.399, -425.1401, -424.3059, -423.7135, -423.7972, -423.9567, 
    -424.7774, -425.5497, -426.1382, -426.5317, -426.9197, -428.0922, 
    -428.7145, -430.1068, -429.8562, -430.2813, -430.6884, -431.371, 
    -431.2587, -431.5593, -430.2706, -431.1268, -429.7133, -430.0998, 
    -427.0226, -425.854, -425.3553, -424.9207, -423.8615, -424.5928, 
    -424.3045, -424.991, -425.4269, -425.2114, -426.5425, -426.0248, 
    -428.7513, -427.5768, -430.6409, -429.9077, -430.8167, -430.353, 
    -431.1474, -430.4325, -431.6714, -431.9409, -431.7567, -432.4652, 
    -430.3928, -431.1883, -425.2053, -425.2404, -425.4044, -424.6836, 
    -424.6396, -423.98, -424.5672, -424.817, -425.4524, -425.8277, -426.1848, 
    -426.9699, -427.8466, -429.0733, -429.9552, -430.5462, -430.184, 
    -430.5038, -430.1462, -429.9787, -431.8398, -430.7945, -432.3633, 
    -432.2766, -431.5664, -432.2864, -425.2651, -425.0629, -424.36, -424.91, 
    -423.9082, -424.4686, -424.7907, -426.0351, -426.3092, -426.5626, 
    -427.0636, -427.7064, -428.834, -429.8156, -430.7122, -430.6465, 
    -430.6696, -430.8697, -430.3738, -430.9511, -431.0477, -430.7947, 
    -432.265, -431.8449, -432.2747, -432.0013, -425.1287, -425.4691, 
    -425.2851, -425.6309, -425.3871, -426.4708, -426.7958, -428.3175, 
    -427.6936, -428.6873, -427.7947, -427.9527, -428.7186, -427.8431, 
    -429.761, -428.4597, -430.8774, -429.5768, -430.9589, -430.7083, 
    -431.1234, -431.495, -431.963, -432.8256, -432.6259, -433.3478, 
    -425.9768, -426.4183, -426.3799, -426.8422, -427.1841, -427.9256, 
    -429.1147, -428.6677, -429.4889, -429.6536, -428.4063, -429.1716, 
    -426.7141, -427.1106, -426.8748, -426.0114, -428.77, -427.3538, 
    -429.9697, -429.2024, -431.442, -430.3276, -432.5159, -433.4502, 
    -434.3318, -435.3595, -426.6597, -426.3597, -426.8973, -427.6404, 
    -428.3312, -429.2491, -429.3433, -429.5151, -429.9608, -430.3353, 
    -429.569, -430.4292, -427.2016, -428.8932, -426.2458, -427.0422, 
    -427.5968, -427.354, -428.6167, -428.9142, -430.123, -429.4984, 
    -433.2192, -431.5728, -436.1436, -434.8659, -426.2548, -426.6589, 
    -428.065, -427.396, -429.3106, -429.7818, -430.1652, -430.6546, 
    -430.7078, -430.9978, -430.5225, -430.9792, -429.251, -430.0234, 
    -427.9048, -428.4201, -428.1832, -427.923, -428.7261, -429.5809, 
    -429.5999, -429.8739, -430.6447, -429.3184, -433.4303, -430.8894, 
    -427.0996, -427.8771, -427.9891, -427.6877, -429.7345, -428.9927, 
    -430.9909, -430.451, -431.3358, -430.8961, -430.8313, -430.2667, 
    -429.915, -429.0266, -428.304, -427.7316, -427.8647, -428.4937, 
    -429.6334, -430.7123, -430.4758, -431.2686, -429.1718, -430.0505, 
    -429.7106, -430.5971, -428.6557, -430.3065, -428.2335, -428.4153, 
    -428.978, -430.1096, -430.3611, -430.6283, -430.4636, -429.6625, 
    -429.5316, -428.9645, -428.8076, -428.3758, -428.018, -428.3447, 
    -428.6877, -429.6631, -430.5418, -431.5002, -431.735, -432.8529, 
    -431.9419, -433.4443, -432.1654, -434.3801, -430.4034, -432.1293, 
    -429.0039, -429.3407, -429.9492, -431.3466, -430.593, -431.4747, 
    -429.5265, -428.515, -428.2542, -427.7662, -428.2654, -428.2248, 
    -428.7025, -428.549, -429.6955, -429.0797, -430.8295, -431.4679, 
    -433.2719, -434.3774, -435.504, -436.0009, -436.1523, -436.2155 ;

 FGR12 =
  -127.4189, -127.4744, -127.4637, -127.5084, -127.4837, -127.513, -127.4302, 
    -127.4766, -127.447, -127.424, -127.596, -127.5105, -127.6865, -127.6312, 
    -127.7708, -127.6778, -127.7898, -127.7684, -127.8334, -127.8147, 
    -127.8979, -127.842, -127.9415, -127.8847, -127.8934, -127.8402, 
    -127.5278, -127.5853, -127.5244, -127.5326, -127.5289, -127.4842, 
    -127.4615, -127.4148, -127.4233, -127.4577, -127.5362, -127.5096, 
    -127.5773, -127.5758, -127.6516, -127.6174, -127.7458, -127.7092, 
    -127.8155, -127.7886, -127.8142, -127.8065, -127.8143, -127.775, 
    -127.7918, -127.7573, -127.6237, -127.6627, -127.5467, -127.4775, 
    -127.4322, -127.4001, -127.4046, -127.4132, -127.4579, -127.5001, 
    -127.5324, -127.5541, -127.5756, -127.6403, -127.6751, -127.7531, 
    -127.7392, -127.763, -127.786, -127.8245, -127.8182, -127.8352, 
    -127.7625, -127.8107, -127.7312, -127.7528, -127.5808, -127.5168, 
    -127.4893, -127.4657, -127.4081, -127.4478, -127.4321, -127.4696, 
    -127.4934, -127.4817, -127.5547, -127.5262, -127.6771, -127.6119, 
    -127.7833, -127.742, -127.7932, -127.7671, -127.8119, -127.7716, 
    -127.8416, -127.8568, -127.8464, -127.8866, -127.7693, -127.8142, 
    -127.4813, -127.4832, -127.4922, -127.4528, -127.4504, -127.4146, 
    -127.4465, -127.4601, -127.4948, -127.5153, -127.535, -127.5783, 
    -127.6268, -127.6952, -127.7447, -127.778, -127.7576, -127.7756, 
    -127.7555, -127.7461, -127.851, -127.7919, -127.8808, -127.8759, 
    -127.8356, -127.8764, -127.4846, -127.4736, -127.4352, -127.4652, 
    -127.4107, -127.4411, -127.4586, -127.5266, -127.5418, -127.5558, 
    -127.5835, -127.6191, -127.6818, -127.7368, -127.7873, -127.7836, 
    -127.7849, -127.7962, -127.7683, -127.8008, -127.8062, -127.792, 
    -127.8752, -127.8514, -127.8758, -127.8603, -127.4772, -127.4957, 
    -127.4857, -127.5045, -127.4912, -127.5506, -127.5686, -127.6529, 
    -127.6184, -127.6736, -127.624, -127.6328, -127.6752, -127.6267, 
    -127.7336, -127.6608, -127.7966, -127.7233, -127.8012, -127.7871, 
    -127.8106, -127.8315, -127.8581, -127.907, -127.8957, -127.9368, 
    -127.5235, -127.5478, -127.5457, -127.5712, -127.5901, -127.6313, 
    -127.6975, -127.6726, -127.7186, -127.7278, -127.6581, -127.7007, 
    -127.5641, -127.5859, -127.573, -127.5254, -127.6782, -127.5995, 
    -127.7455, -127.7025, -127.8285, -127.7656, -127.8895, -127.9425, 
    -127.9932, -128.0521, -127.5611, -127.5446, -127.5743, -127.6153, 
    -127.6538, -127.7051, -127.7104, -127.72, -127.745, -127.7661, -127.7229, 
    -127.7714, -127.5908, -127.6851, -127.5383, -127.5821, -127.613, 
    -127.5995, -127.6698, -127.6864, -127.7541, -127.7191, -127.9293, 
    -127.8358, -128.0975, -128.0237, -127.5389, -127.5611, -127.639, 
    -127.6019, -127.7086, -127.7349, -127.7565, -127.784, -127.7871, 
    -127.8034, -127.7766, -127.8024, -127.7052, -127.7485, -127.6302, 
    -127.6588, -127.6456, -127.6312, -127.6759, -127.7236, -127.7248, 
    -127.7401, -127.783, -127.709, -127.941, -127.797, -127.5855, -127.6284, 
    -127.6348, -127.6181, -127.7323, -127.6908, -127.803, -127.7726, 
    -127.8225, -127.7977, -127.794, -127.7622, -127.7424, -127.6926, 
    -127.6523, -127.6206, -127.628, -127.6629, -127.7266, -127.7873, 
    -127.7739, -127.8187, -127.7008, -127.75, -127.7309, -127.7808, -127.672, 
    -127.764, -127.6485, -127.6586, -127.6899, -127.7532, -127.7676, 
    -127.7825, -127.7733, -127.7282, -127.7209, -127.6892, -127.6804, 
    -127.6564, -127.6365, -127.6546, -127.6737, -127.7283, -127.7777, 
    -127.8318, -127.8452, -127.9083, -127.8567, -127.9418, -127.8691, 
    -127.9956, -127.7697, -127.8672, -127.6914, -127.7103, -127.7443, 
    -127.823, -127.7806, -127.8303, -127.7206, -127.664, -127.6496, 
    -127.6225, -127.6502, -127.648, -127.6746, -127.666, -127.7301, 
    -127.6957, -127.7939, -127.8299, -127.9325, -127.9956, -128.0606, 
    -128.0894, -128.0981, -128.1018 ;

 FGR_R =
  -424.0618, -425.0807, -424.8828, -425.7042, -425.2488, -425.7865, 
    -424.2686, -425.1208, -424.577, -424.1539, -427.298, -425.7409, 
    -428.9189, -427.9251, -430.423, -428.7639, -430.7577, -430.3759, 
    -431.527, -431.1973, -432.6681, -431.6792, -433.4318, -432.4323, 
    -432.5884, -431.6465, -426.0549, -427.1039, -425.9926, -426.1422, 
    -426.0753, -425.258, -424.8456, -423.9844, -424.1409, -424.7737, 
    -426.2095, -425.7225, -426.9514, -426.9237, -428.2916, -427.6748, 
    -429.975, -429.3214, -431.211, -430.7357, -431.1886, -431.0513, 
    -431.1904, -430.4932, -430.7918, -430.1787, -427.7902, -428.4918, 
    -426.399, -425.1401, -424.3059, -423.7135, -423.7972, -423.9567, 
    -424.7774, -425.5497, -426.1382, -426.5317, -426.9197, -428.0922, 
    -428.7145, -430.1068, -429.8562, -430.2813, -430.6884, -431.371, 
    -431.2587, -431.5593, -430.2706, -431.1268, -429.7133, -430.0998, 
    -427.0226, -425.854, -425.3553, -424.9207, -423.8615, -424.5928, 
    -424.3045, -424.991, -425.4269, -425.2114, -426.5425, -426.0248, 
    -428.7513, -427.5768, -430.6409, -429.9077, -430.8167, -430.353, 
    -431.1474, -430.4325, -431.6714, -431.9409, -431.7567, -432.4652, 
    -430.3928, -431.1883, -425.2053, -425.2404, -425.4044, -424.6836, 
    -424.6396, -423.98, -424.5672, -424.817, -425.4524, -425.8277, -426.1848, 
    -426.9699, -427.8466, -429.0733, -429.9552, -430.5462, -430.184, 
    -430.5038, -430.1462, -429.9787, -431.8398, -430.7945, -432.3633, 
    -432.2766, -431.5664, -432.2864, -425.2651, -425.0629, -424.36, -424.91, 
    -423.9082, -424.4686, -424.7907, -426.0351, -426.3092, -426.5626, 
    -427.0636, -427.7064, -428.834, -429.8156, -430.7122, -430.6465, 
    -430.6696, -430.8697, -430.3738, -430.9511, -431.0477, -430.7947, 
    -432.265, -431.8449, -432.2747, -432.0013, -425.1287, -425.4691, 
    -425.2851, -425.6309, -425.3871, -426.4708, -426.7958, -428.3175, 
    -427.6936, -428.6873, -427.7947, -427.9527, -428.7186, -427.8431, 
    -429.761, -428.4597, -430.8774, -429.5768, -430.9589, -430.7083, 
    -431.1234, -431.495, -431.963, -432.8256, -432.6259, -433.3478, 
    -425.9768, -426.4183, -426.3799, -426.8422, -427.1841, -427.9256, 
    -429.1147, -428.6677, -429.4889, -429.6536, -428.4063, -429.1716, 
    -426.7141, -427.1106, -426.8748, -426.0114, -428.77, -427.3538, 
    -429.9697, -429.2024, -431.442, -430.3276, -432.5159, -433.4502, 
    -434.3318, -435.3595, -426.6597, -426.3597, -426.8973, -427.6404, 
    -428.3312, -429.2491, -429.3433, -429.5151, -429.9608, -430.3353, 
    -429.569, -430.4292, -427.2016, -428.8932, -426.2458, -427.0422, 
    -427.5968, -427.354, -428.6167, -428.9142, -430.123, -429.4984, 
    -433.2192, -431.5728, -436.1436, -434.8659, -426.2548, -426.6589, 
    -428.065, -427.396, -429.3106, -429.7818, -430.1652, -430.6546, 
    -430.7078, -430.9978, -430.5225, -430.9792, -429.251, -430.0234, 
    -427.9048, -428.4201, -428.1832, -427.923, -428.7261, -429.5809, 
    -429.5999, -429.8739, -430.6447, -429.3184, -433.4303, -430.8894, 
    -427.0996, -427.8771, -427.9891, -427.6877, -429.7345, -428.9927, 
    -430.9909, -430.451, -431.3358, -430.8961, -430.8313, -430.2667, 
    -429.915, -429.0266, -428.304, -427.7316, -427.8647, -428.4937, 
    -429.6334, -430.7123, -430.4758, -431.2686, -429.1718, -430.0505, 
    -429.7106, -430.5971, -428.6557, -430.3065, -428.2335, -428.4153, 
    -428.978, -430.1096, -430.3611, -430.6283, -430.4636, -429.6625, 
    -429.5316, -428.9645, -428.8076, -428.3758, -428.018, -428.3447, 
    -428.6877, -429.6631, -430.5418, -431.5002, -431.735, -432.8529, 
    -431.9419, -433.4443, -432.1654, -434.3801, -430.4034, -432.1293, 
    -429.0039, -429.3407, -429.9492, -431.3466, -430.593, -431.4747, 
    -429.5265, -428.515, -428.2542, -427.7662, -428.2654, -428.2248, 
    -428.7025, -428.549, -429.6955, -429.0797, -430.8295, -431.4679, 
    -433.2719, -434.3774, -435.504, -436.0009, -436.1523, -436.2155 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  48.80871, 48.87994, 48.86611, 48.92353, 48.8917, 48.92929, 48.82317, 
    48.88275, 48.84473, 48.81516, 49.03493, 48.92611, 49.14824, 49.07878, 
    49.25336, 49.1374, 49.27675, 49.25007, 49.33052, 49.30748, 49.41026, 
    49.34116, 49.46364, 49.39379, 49.4047, 49.33887, 48.94806, 49.02137, 
    48.9437, 48.95416, 48.94948, 48.89234, 48.86351, 48.8033, 48.81424, 
    48.85848, 48.95886, 48.92482, 49.01073, 49.00879, 49.1044, 49.06129, 
    49.22205, 49.17637, 49.30844, 49.27522, 49.30687, 49.29728, 49.307, 
    49.25827, 49.27914, 49.23629, 49.06935, 49.11839, 48.97211, 48.88409, 
    48.82578, 48.78436, 48.79021, 48.80136, 48.85874, 48.91274, 48.95388, 
    48.98139, 49.00851, 49.09045, 49.13395, 49.23127, 49.21375, 49.24346, 
    49.27192, 49.31962, 49.31178, 49.33278, 49.24271, 49.30256, 49.20376, 
    49.23077, 49.01569, 48.93401, 48.89914, 48.86876, 48.79471, 48.84583, 
    48.82568, 48.87368, 48.90415, 48.88909, 48.98214, 48.94596, 49.13652, 
    49.05444, 49.26859, 49.21735, 49.28088, 49.24847, 49.30399, 49.25403, 
    49.34062, 49.35945, 49.34658, 49.3961, 49.25125, 49.30685, 48.88866, 
    48.89111, 48.90258, 48.85218, 48.84911, 48.80299, 48.84405, 48.86152, 
    48.90593, 48.93217, 48.95713, 49.01202, 49.07329, 49.15903, 49.22067, 
    49.26198, 49.23666, 49.25901, 49.23402, 49.22231, 49.35238, 49.27933, 
    49.38897, 49.38291, 49.33327, 49.38359, 48.89284, 48.8787, 48.82956, 
    48.86802, 48.79797, 48.83715, 48.85967, 48.94667, 48.96584, 48.98354, 
    49.01857, 49.06349, 49.1423, 49.21091, 49.27358, 49.26899, 49.2706, 
    49.28458, 49.24993, 49.29027, 49.29703, 49.27934, 49.3821, 49.35275, 
    49.38278, 49.36367, 48.8833, 48.9071, 48.89424, 48.91842, 48.90137, 
    48.97713, 48.99984, 49.1062, 49.0626, 49.13205, 49.06967, 49.08071, 
    49.13423, 49.07305, 49.20709, 49.11614, 49.28513, 49.19421, 49.29082, 
    49.27331, 49.30232, 49.32829, 49.36099, 49.42128, 49.40733, 49.45778, 
    48.9426, 48.97345, 48.97078, 49.00309, 49.02699, 49.07882, 49.16193, 
    49.13068, 49.18808, 49.19959, 49.11242, 49.1659, 48.99413, 49.02184, 
    49.00537, 48.94501, 49.13783, 49.03885, 49.22168, 49.16806, 49.32458, 
    49.2467, 49.39964, 49.46492, 49.52654, 49.59835, 48.99033, 48.96936, 
    49.00695, 49.05888, 49.10717, 49.17132, 49.1779, 49.18991, 49.22106, 
    49.24723, 49.19367, 49.2538, 49.0282, 49.14644, 48.9614, 49.01707, 
    49.05583, 49.03886, 49.12712, 49.14791, 49.2324, 49.18874, 49.44878, 
    49.33372, 49.65315, 49.56386, 48.96203, 48.99028, 49.08856, 49.0418, 
    49.17562, 49.20855, 49.23535, 49.26955, 49.27327, 49.29354, 49.26032, 
    49.29224, 49.17146, 49.22544, 49.07737, 49.11338, 49.09682, 49.07864, 
    49.13477, 49.19451, 49.19584, 49.21499, 49.26884, 49.17617, 49.46352, 
    49.28595, 49.02108, 49.07542, 49.08326, 49.06219, 49.20525, 49.1534, 
    49.29306, 49.25532, 49.31716, 49.28643, 49.2819, 49.24244, 49.21786, 
    49.15577, 49.10527, 49.06526, 49.07457, 49.11852, 49.19817, 49.27358, 
    49.25705, 49.31247, 49.16592, 49.22733, 49.20358, 49.26553, 49.12984, 
    49.24521, 49.10033, 49.11305, 49.15237, 49.23146, 49.24904, 49.26772, 
    49.25621, 49.20021, 49.19106, 49.15143, 49.14046, 49.11029, 49.08528, 
    49.10811, 49.13208, 49.20026, 49.26167, 49.32865, 49.34507, 49.42318, 
    49.35951, 49.4645, 49.37512, 49.5299, 49.25198, 49.3726, 49.15418, 
    49.17772, 49.22025, 49.31791, 49.26524, 49.32686, 49.19071, 49.12001, 
    49.10179, 49.06768, 49.10257, 49.09973, 49.13311, 49.12239, 49.20252, 
    49.15948, 49.28177, 49.32639, 49.45247, 49.52972, 49.60846, 49.64318, 
    49.65376, 49.65818 ;

 FIRA_R =
  48.80871, 48.87994, 48.86611, 48.92353, 48.8917, 48.92929, 48.82317, 
    48.88275, 48.84473, 48.81516, 49.03493, 48.92611, 49.14824, 49.07878, 
    49.25336, 49.1374, 49.27675, 49.25007, 49.33052, 49.30748, 49.41026, 
    49.34116, 49.46364, 49.39379, 49.4047, 49.33887, 48.94806, 49.02137, 
    48.9437, 48.95416, 48.94948, 48.89234, 48.86351, 48.8033, 48.81424, 
    48.85848, 48.95886, 48.92482, 49.01073, 49.00879, 49.1044, 49.06129, 
    49.22205, 49.17637, 49.30844, 49.27522, 49.30687, 49.29728, 49.307, 
    49.25827, 49.27914, 49.23629, 49.06935, 49.11839, 48.97211, 48.88409, 
    48.82578, 48.78436, 48.79021, 48.80136, 48.85874, 48.91274, 48.95388, 
    48.98139, 49.00851, 49.09045, 49.13395, 49.23127, 49.21375, 49.24346, 
    49.27192, 49.31962, 49.31178, 49.33278, 49.24271, 49.30256, 49.20376, 
    49.23077, 49.01569, 48.93401, 48.89914, 48.86876, 48.79471, 48.84583, 
    48.82568, 48.87368, 48.90415, 48.88909, 48.98214, 48.94596, 49.13652, 
    49.05444, 49.26859, 49.21735, 49.28088, 49.24847, 49.30399, 49.25403, 
    49.34062, 49.35945, 49.34658, 49.3961, 49.25125, 49.30685, 48.88866, 
    48.89111, 48.90258, 48.85218, 48.84911, 48.80299, 48.84405, 48.86152, 
    48.90593, 48.93217, 48.95713, 49.01202, 49.07329, 49.15903, 49.22067, 
    49.26198, 49.23666, 49.25901, 49.23402, 49.22231, 49.35238, 49.27933, 
    49.38897, 49.38291, 49.33327, 49.38359, 48.89284, 48.8787, 48.82956, 
    48.86802, 48.79797, 48.83715, 48.85967, 48.94667, 48.96584, 48.98354, 
    49.01857, 49.06349, 49.1423, 49.21091, 49.27358, 49.26899, 49.2706, 
    49.28458, 49.24993, 49.29027, 49.29703, 49.27934, 49.3821, 49.35275, 
    49.38278, 49.36367, 48.8833, 48.9071, 48.89424, 48.91842, 48.90137, 
    48.97713, 48.99984, 49.1062, 49.0626, 49.13205, 49.06967, 49.08071, 
    49.13423, 49.07305, 49.20709, 49.11614, 49.28513, 49.19421, 49.29082, 
    49.27331, 49.30232, 49.32829, 49.36099, 49.42128, 49.40733, 49.45778, 
    48.9426, 48.97345, 48.97078, 49.00309, 49.02699, 49.07882, 49.16193, 
    49.13068, 49.18808, 49.19959, 49.11242, 49.1659, 48.99413, 49.02184, 
    49.00537, 48.94501, 49.13783, 49.03885, 49.22168, 49.16806, 49.32458, 
    49.2467, 49.39964, 49.46492, 49.52654, 49.59835, 48.99033, 48.96936, 
    49.00695, 49.05888, 49.10717, 49.17132, 49.1779, 49.18991, 49.22106, 
    49.24723, 49.19367, 49.2538, 49.0282, 49.14644, 48.9614, 49.01707, 
    49.05583, 49.03886, 49.12712, 49.14791, 49.2324, 49.18874, 49.44878, 
    49.33372, 49.65315, 49.56386, 48.96203, 48.99028, 49.08856, 49.0418, 
    49.17562, 49.20855, 49.23535, 49.26955, 49.27327, 49.29354, 49.26032, 
    49.29224, 49.17146, 49.22544, 49.07737, 49.11338, 49.09682, 49.07864, 
    49.13477, 49.19451, 49.19584, 49.21499, 49.26884, 49.17617, 49.46352, 
    49.28595, 49.02108, 49.07542, 49.08326, 49.06219, 49.20525, 49.1534, 
    49.29306, 49.25532, 49.31716, 49.28643, 49.2819, 49.24244, 49.21786, 
    49.15577, 49.10527, 49.06526, 49.07457, 49.11852, 49.19817, 49.27358, 
    49.25705, 49.31247, 49.16592, 49.22733, 49.20358, 49.26553, 49.12984, 
    49.24521, 49.10033, 49.11305, 49.15237, 49.23146, 49.24904, 49.26772, 
    49.25621, 49.20021, 49.19106, 49.15143, 49.14046, 49.11029, 49.08528, 
    49.10811, 49.13208, 49.20026, 49.26167, 49.32865, 49.34507, 49.42318, 
    49.35951, 49.4645, 49.37512, 49.5299, 49.25198, 49.3726, 49.15418, 
    49.17772, 49.22025, 49.31791, 49.26524, 49.32686, 49.19071, 49.12001, 
    49.10179, 49.06768, 49.10257, 49.09973, 49.13311, 49.12239, 49.20252, 
    49.15948, 49.28177, 49.32639, 49.45247, 49.52972, 49.60846, 49.64318, 
    49.65376, 49.65818 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.1548, 263.2261, 263.2122, 263.2697, 263.2379, 263.2754, 263.1693, 
    263.2289, 263.1909, 263.1613, 263.3811, 263.2722, 263.4944, 263.4249, 
    263.5995, 263.4836, 263.6229, 263.5962, 263.6767, 263.6536, 263.7564, 
    263.6873, 263.8098, 263.7399, 263.7509, 263.685, 263.2942, 263.3675, 
    263.2899, 263.3003, 263.2956, 263.2385, 263.2097, 263.1494, 263.1604, 
    263.2046, 263.305, 263.271, 263.3569, 263.3549, 263.4505, 263.4074, 
    263.5682, 263.5225, 263.6546, 263.6214, 263.653, 263.6434, 263.6531, 
    263.6044, 263.6253, 263.5824, 263.4155, 263.4645, 263.3183, 263.2302, 
    263.1719, 263.1305, 263.1364, 263.1475, 263.2049, 263.2589, 263.3, 
    263.3275, 263.3546, 263.4366, 263.4801, 263.5774, 263.5599, 263.5896, 
    263.6181, 263.6658, 263.6579, 263.6789, 263.5889, 263.6487, 263.5499, 
    263.5769, 263.3618, 263.2802, 263.2453, 263.2149, 263.1409, 263.192, 
    263.1718, 263.2198, 263.2503, 263.2352, 263.3283, 263.2921, 263.4827, 
    263.4006, 263.6147, 263.5635, 263.627, 263.5946, 263.6501, 263.6002, 
    263.6868, 263.7056, 263.6927, 263.7422, 263.5974, 263.653, 263.2348, 
    263.2372, 263.2487, 263.1983, 263.1953, 263.1491, 263.1902, 263.2077, 
    263.2521, 263.2783, 263.3033, 263.3582, 263.4194, 263.5052, 263.5668, 
    263.6081, 263.5828, 263.6052, 263.5802, 263.5685, 263.6985, 263.6255, 
    263.7351, 263.7291, 263.6794, 263.7297, 263.239, 263.2249, 263.1757, 
    263.2142, 263.1441, 263.1833, 263.2058, 263.2928, 263.312, 263.3297, 
    263.3647, 263.4096, 263.4884, 263.5571, 263.6197, 263.6151, 263.6168, 
    263.6307, 263.5961, 263.6364, 263.6432, 263.6255, 263.7282, 263.6989, 
    263.7289, 263.7098, 263.2295, 263.2532, 263.2404, 263.2646, 263.2475, 
    263.3233, 263.346, 263.4523, 263.4088, 263.4782, 263.4158, 263.4268, 
    263.4804, 263.4192, 263.5532, 263.4623, 263.6313, 263.5403, 263.637, 
    263.6194, 263.6485, 263.6744, 263.7071, 263.7674, 263.7535, 263.8039, 
    263.2888, 263.3196, 263.3169, 263.3492, 263.3731, 263.425, 263.5081, 
    263.4768, 263.5342, 263.5457, 263.4586, 263.5121, 263.3403, 263.368, 
    263.3515, 263.2912, 263.484, 263.385, 263.5678, 263.5142, 263.6707, 
    263.5928, 263.7458, 263.8111, 263.8727, 263.9445, 263.3365, 263.3155, 
    263.3531, 263.405, 263.4533, 263.5175, 263.524, 263.536, 263.5672, 
    263.5934, 263.5398, 263.5999, 263.3743, 263.4926, 263.3076, 263.3632, 
    263.402, 263.385, 263.4733, 263.494, 263.5786, 263.5349, 263.7949, 
    263.6799, 263.9993, 263.91, 263.3082, 263.3364, 263.4347, 263.3879, 
    263.5218, 263.5547, 263.5815, 263.6157, 263.6194, 263.6397, 263.6065, 
    263.6384, 263.5176, 263.5716, 263.4235, 263.4595, 263.443, 263.4248, 
    263.4809, 263.5406, 263.542, 263.5611, 263.615, 263.5223, 263.8097, 
    263.6321, 263.3672, 263.4216, 263.4294, 263.4083, 263.5514, 263.4995, 
    263.6392, 263.6015, 263.6633, 263.6326, 263.6281, 263.5886, 263.564, 
    263.5019, 263.4514, 263.4114, 263.4207, 263.4647, 263.5443, 263.6197, 
    263.6032, 263.6586, 263.5121, 263.5735, 263.5497, 263.6117, 263.476, 
    263.5913, 263.4465, 263.4592, 263.4985, 263.5776, 263.5952, 263.6139, 
    263.6024, 263.5464, 263.5372, 263.4976, 263.4866, 263.4564, 263.4314, 
    263.4543, 263.4782, 263.5464, 263.6078, 263.6748, 263.6912, 263.7693, 
    263.7057, 263.8106, 263.7213, 263.876, 263.5981, 263.7188, 263.5003, 
    263.5239, 263.5664, 263.6641, 263.6114, 263.673, 263.5369, 263.4662, 
    263.4479, 263.4138, 263.4487, 263.4459, 263.4792, 263.4685, 263.5487, 
    263.5056, 263.6279, 263.6725, 263.7986, 263.8759, 263.9546, 263.9893, 
    263.9999, 264.0043 ;

 FIRE_R =
  263.1548, 263.2261, 263.2122, 263.2697, 263.2379, 263.2754, 263.1693, 
    263.2289, 263.1909, 263.1613, 263.3811, 263.2722, 263.4944, 263.4249, 
    263.5995, 263.4836, 263.6229, 263.5962, 263.6767, 263.6536, 263.7564, 
    263.6873, 263.8098, 263.7399, 263.7509, 263.685, 263.2942, 263.3675, 
    263.2899, 263.3003, 263.2956, 263.2385, 263.2097, 263.1494, 263.1604, 
    263.2046, 263.305, 263.271, 263.3569, 263.3549, 263.4505, 263.4074, 
    263.5682, 263.5225, 263.6546, 263.6214, 263.653, 263.6434, 263.6531, 
    263.6044, 263.6253, 263.5824, 263.4155, 263.4645, 263.3183, 263.2302, 
    263.1719, 263.1305, 263.1364, 263.1475, 263.2049, 263.2589, 263.3, 
    263.3275, 263.3546, 263.4366, 263.4801, 263.5774, 263.5599, 263.5896, 
    263.6181, 263.6658, 263.6579, 263.6789, 263.5889, 263.6487, 263.5499, 
    263.5769, 263.3618, 263.2802, 263.2453, 263.2149, 263.1409, 263.192, 
    263.1718, 263.2198, 263.2503, 263.2352, 263.3283, 263.2921, 263.4827, 
    263.4006, 263.6147, 263.5635, 263.627, 263.5946, 263.6501, 263.6002, 
    263.6868, 263.7056, 263.6927, 263.7422, 263.5974, 263.653, 263.2348, 
    263.2372, 263.2487, 263.1983, 263.1953, 263.1491, 263.1902, 263.2077, 
    263.2521, 263.2783, 263.3033, 263.3582, 263.4194, 263.5052, 263.5668, 
    263.6081, 263.5828, 263.6052, 263.5802, 263.5685, 263.6985, 263.6255, 
    263.7351, 263.7291, 263.6794, 263.7297, 263.239, 263.2249, 263.1757, 
    263.2142, 263.1441, 263.1833, 263.2058, 263.2928, 263.312, 263.3297, 
    263.3647, 263.4096, 263.4884, 263.5571, 263.6197, 263.6151, 263.6168, 
    263.6307, 263.5961, 263.6364, 263.6432, 263.6255, 263.7282, 263.6989, 
    263.7289, 263.7098, 263.2295, 263.2532, 263.2404, 263.2646, 263.2475, 
    263.3233, 263.346, 263.4523, 263.4088, 263.4782, 263.4158, 263.4268, 
    263.4804, 263.4192, 263.5532, 263.4623, 263.6313, 263.5403, 263.637, 
    263.6194, 263.6485, 263.6744, 263.7071, 263.7674, 263.7535, 263.8039, 
    263.2888, 263.3196, 263.3169, 263.3492, 263.3731, 263.425, 263.5081, 
    263.4768, 263.5342, 263.5457, 263.4586, 263.5121, 263.3403, 263.368, 
    263.3515, 263.2912, 263.484, 263.385, 263.5678, 263.5142, 263.6707, 
    263.5928, 263.7458, 263.8111, 263.8727, 263.9445, 263.3365, 263.3155, 
    263.3531, 263.405, 263.4533, 263.5175, 263.524, 263.536, 263.5672, 
    263.5934, 263.5398, 263.5999, 263.3743, 263.4926, 263.3076, 263.3632, 
    263.402, 263.385, 263.4733, 263.494, 263.5786, 263.5349, 263.7949, 
    263.6799, 263.9993, 263.91, 263.3082, 263.3364, 263.4347, 263.3879, 
    263.5218, 263.5547, 263.5815, 263.6157, 263.6194, 263.6397, 263.6065, 
    263.6384, 263.5176, 263.5716, 263.4235, 263.4595, 263.443, 263.4248, 
    263.4809, 263.5406, 263.542, 263.5611, 263.615, 263.5223, 263.8097, 
    263.6321, 263.3672, 263.4216, 263.4294, 263.4083, 263.5514, 263.4995, 
    263.6392, 263.6015, 263.6633, 263.6326, 263.6281, 263.5886, 263.564, 
    263.5019, 263.4514, 263.4114, 263.4207, 263.4647, 263.5443, 263.6197, 
    263.6032, 263.6586, 263.5121, 263.5735, 263.5497, 263.6117, 263.476, 
    263.5913, 263.4465, 263.4592, 263.4985, 263.5776, 263.5952, 263.6139, 
    263.6024, 263.5464, 263.5372, 263.4976, 263.4866, 263.4564, 263.4314, 
    263.4543, 263.4782, 263.5464, 263.6078, 263.6748, 263.6912, 263.7693, 
    263.7057, 263.8106, 263.7213, 263.876, 263.5981, 263.7188, 263.5003, 
    263.5239, 263.5664, 263.6641, 263.6114, 263.673, 263.5369, 263.4662, 
    263.4479, 263.4138, 263.4487, 263.4459, 263.4792, 263.4685, 263.5487, 
    263.5056, 263.6279, 263.6725, 263.7986, 263.8759, 263.9546, 263.9893, 
    263.9999, 264.0043 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  351.6926, 352.5784, 352.4064, 353.1205, 352.7246, 353.192, 351.8725, 
    352.6134, 352.1405, 351.7727, 354.5061, 353.1524, 355.9149, 355.051, 
    357.222, 355.7801, 357.5129, 357.181, 358.1813, 357.8948, 359.173, 
    358.3136, 359.8365, 358.9681, 359.1037, 358.2852, 353.4254, 354.3373, 
    353.3712, 353.5013, 353.443, 352.7326, 352.3741, 351.6253, 351.7614, 
    352.3116, 353.5598, 353.1364, 354.2047, 354.1805, 355.3696, 354.8335, 
    356.8327, 356.2646, 357.9068, 357.4937, 357.8873, 357.768, 357.8888, 
    357.283, 357.5425, 357.0096, 354.9337, 355.5436, 353.7245, 352.6302, 
    351.9048, 351.3898, 351.4626, 351.6013, 352.3148, 352.9862, 353.4977, 
    353.8398, 354.1771, 355.1964, 355.7372, 356.9473, 356.7294, 357.0989, 
    357.4526, 358.0458, 357.9482, 358.2095, 357.0895, 357.8336, 356.6052, 
    356.9411, 354.2668, 353.2507, 352.8173, 352.4394, 351.5185, 352.1543, 
    351.9036, 352.5005, 352.8794, 352.6921, 353.8492, 353.3992, 355.7692, 
    354.7483, 357.4113, 356.7741, 357.5641, 357.1611, 357.8515, 357.2302, 
    358.3069, 358.5411, 358.381, 358.9966, 357.1957, 357.8871, 352.6867, 
    352.7173, 352.8598, 352.2332, 352.195, 351.6215, 352.132, 352.3492, 
    352.9016, 353.2278, 353.5382, 354.2208, 354.9828, 356.049, 356.8154, 
    357.3291, 357.0143, 357.2922, 356.9814, 356.8358, 358.4532, 357.5448, 
    358.9081, 358.8327, 358.2156, 358.8412, 352.7388, 352.5629, 351.9518, 
    352.4301, 351.5591, 352.0464, 352.3264, 353.4082, 353.6464, 353.8666, 
    354.3022, 354.8609, 355.841, 356.6941, 357.4733, 357.4162, 357.4363, 
    357.6101, 357.1792, 357.6809, 357.7649, 357.545, 358.8226, 358.4576, 
    358.8311, 358.5935, 352.6201, 352.9161, 352.7561, 353.0568, 352.8448, 
    353.7869, 354.0695, 355.3921, 354.8498, 355.7135, 354.9377, 355.075, 
    355.7408, 354.9797, 356.6467, 355.5157, 357.6169, 356.4867, 357.6877, 
    357.4699, 357.8307, 358.1536, 358.5602, 359.3098, 359.1363, 359.7635, 
    353.3575, 353.7412, 353.7078, 354.1097, 354.4069, 355.0515, 356.085, 
    355.6964, 356.4102, 356.5533, 355.4692, 356.1345, 353.9984, 354.343, 
    354.1381, 353.3875, 355.7855, 354.5545, 356.828, 356.1612, 358.1075, 
    357.1392, 359.0407, 359.8526, 360.6185, 361.5114, 353.9511, 353.6903, 
    354.1576, 354.8036, 355.404, 356.2018, 356.2836, 356.433, 356.8203, 
    357.1457, 356.4798, 357.2274, 354.4223, 355.8925, 353.5913, 354.2837, 
    354.7657, 354.5546, 355.6521, 355.9107, 356.9613, 356.4184, 359.6519, 
    358.2213, 362.1925, 361.0826, 353.5991, 353.9504, 355.1726, 354.5911, 
    356.2552, 356.6647, 356.9979, 357.4233, 357.4695, 357.7216, 357.3084, 
    357.7054, 356.2035, 356.8747, 355.0334, 355.4813, 355.2754, 355.0492, 
    355.7472, 356.4902, 356.5067, 356.7448, 357.4149, 356.262, 359.8354, 
    357.6275, 354.3334, 355.0094, 355.1067, 354.8447, 356.6236, 355.9789, 
    357.7155, 357.2463, 358.0152, 357.6331, 357.5768, 357.0861, 356.7805, 
    356.0084, 355.3804, 354.8828, 354.9985, 355.5452, 356.5358, 357.4734, 
    357.2679, 357.9568, 356.1346, 356.8983, 356.6029, 357.3733, 355.686, 
    357.1209, 355.319, 355.4771, 355.9662, 356.9497, 357.1682, 357.4005, 
    357.2573, 356.5611, 356.4473, 355.9544, 355.8181, 355.4427, 355.1317, 
    355.4157, 355.7139, 356.5616, 357.3253, 358.1581, 358.3622, 359.3337, 
    358.542, 359.8476, 358.7363, 360.6606, 357.205, 358.7048, 355.9886, 
    356.2814, 356.8103, 358.0246, 357.3697, 358.136, 356.4428, 355.5638, 
    355.3371, 354.9129, 355.3468, 355.3115, 355.7267, 355.5933, 356.5898, 
    356.0545, 357.5753, 358.1301, 359.6976, 360.6581, 361.6368, 362.0685, 
    362.2, 362.2549 ;

 FSH_G =
  358.3519, 359.2383, 359.0661, 359.7806, 359.3845, 359.8522, 358.5319, 
    359.2732, 358.8001, 358.4321, 361.1671, 359.8126, 362.5768, 361.7123, 
    363.8847, 362.4419, 364.1758, 363.8437, 364.8446, 364.5579, 365.8369, 
    364.977, 366.5009, 365.6319, 365.7676, 364.9485, 360.0857, 360.9982, 
    360.0315, 360.1617, 360.1034, 359.3925, 359.0338, 358.2846, 358.4207, 
    358.9712, 360.2202, 359.7966, 360.8655, 360.8414, 362.0312, 361.4947, 
    363.4951, 362.9267, 364.5699, 364.1566, 364.5504, 364.4311, 364.5519, 
    363.9457, 364.2054, 363.6722, 361.595, 362.2053, 360.385, 359.29, 
    358.5643, 358.0489, 358.1217, 358.2605, 358.9744, 359.6462, 360.1581, 
    360.5005, 360.8379, 361.8578, 362.399, 363.6098, 363.3918, 363.7615, 
    364.1154, 364.709, 364.6114, 364.8728, 363.7521, 364.4967, 363.2675, 
    363.6036, 360.9276, 359.9109, 359.4772, 359.0991, 358.1777, 358.8139, 
    358.563, 359.1602, 359.5394, 359.352, 360.5098, 360.0595, 362.431, 
    361.4095, 364.0742, 363.4366, 364.2271, 363.8238, 364.5146, 363.8929, 
    364.9702, 365.2046, 365.0444, 365.6605, 363.8584, 364.5502, 359.3466, 
    359.3772, 359.5198, 358.8929, 358.8546, 358.2807, 358.7916, 359.0089, 
    359.5616, 359.8881, 360.1986, 360.8816, 361.6441, 362.711, 363.4779, 
    363.9919, 363.6768, 363.9549, 363.644, 363.4983, 365.1166, 364.2077, 
    365.5718, 365.4964, 364.8789, 365.5049, 359.3987, 359.2227, 358.6113, 
    359.0898, 358.2183, 358.7058, 358.9861, 360.0685, 360.3069, 360.5273, 
    360.963, 361.5221, 362.5028, 363.3565, 364.1361, 364.079, 364.0991, 
    364.2731, 363.8419, 364.3439, 364.4279, 364.2079, 365.4863, 365.1211, 
    365.4948, 365.2571, 359.28, 359.5761, 359.4161, 359.7169, 359.5048, 
    360.4475, 360.7302, 362.0537, 361.511, 362.3752, 361.5989, 361.7364, 
    362.4026, 361.641, 363.309, 362.1774, 364.2798, 363.1489, 364.3507, 
    364.1328, 364.4938, 364.8169, 365.2237, 365.9738, 365.8002, 366.4278, 
    360.0178, 360.4018, 360.3683, 360.7705, 361.0678, 361.7128, 362.7469, 
    362.3582, 363.0724, 363.2156, 362.1309, 362.7965, 360.6591, 361.004, 
    360.7989, 360.0479, 362.4472, 361.2155, 363.4905, 362.8232, 364.7708, 
    363.8018, 365.7046, 366.5169, 367.2833, 368.1768, 360.6118, 360.3508, 
    360.8184, 361.4648, 362.0656, 362.8638, 362.9457, 363.0952, 363.4827, 
    363.8084, 363.142, 363.89, 361.0832, 362.5544, 360.2518, 360.9445, 
    361.4268, 361.2157, 362.3139, 362.5726, 363.6238, 363.0806, 366.3161, 
    364.8846, 368.8583, 367.7477, 360.2595, 360.6111, 361.8341, 361.2522, 
    362.9173, 363.3271, 363.6605, 364.0861, 364.1323, 364.3846, 363.9712, 
    364.3684, 362.8655, 363.5372, 361.6947, 362.1429, 361.9369, 361.7106, 
    362.409, 363.1524, 363.1689, 363.4072, 364.0777, 362.9241, 366.4997, 
    364.2904, 360.9944, 361.6707, 361.7681, 361.5059, 363.2859, 362.6409, 
    364.3785, 363.909, 364.6784, 364.296, 364.2397, 363.7487, 363.4429, 
    362.6703, 362.042, 361.544, 361.6599, 362.2068, 363.1981, 364.1362, 
    363.9306, 364.62, 362.7966, 363.5608, 363.2652, 364.0361, 362.3477, 
    363.7836, 361.9805, 362.1387, 362.6281, 363.6122, 363.8309, 364.0632, 
    363.92, 363.2233, 363.1095, 362.6163, 362.4799, 362.1043, 361.7932, 
    362.0773, 362.3756, 363.2239, 363.988, 364.8214, 365.0256, 365.9977, 
    365.2055, 366.5119, 365.3999, 367.3254, 363.8677, 365.3684, 362.6506, 
    362.9435, 363.4727, 364.6878, 364.0325, 364.7992, 363.1051, 362.2254, 
    361.9986, 361.5742, 362.0083, 361.973, 362.3884, 362.255, 363.252, 
    362.7165, 364.2382, 364.7933, 366.3618, 367.3229, 368.3023, 368.7343, 
    368.8658, 368.9208 ;

 FSH_NODYNLNDUSE =
  351.6926, 352.5784, 352.4064, 353.1205, 352.7246, 353.192, 351.8725, 
    352.6134, 352.1405, 351.7727, 354.5061, 353.1524, 355.9149, 355.051, 
    357.222, 355.7801, 357.5129, 357.181, 358.1813, 357.8948, 359.173, 
    358.3136, 359.8365, 358.9681, 359.1037, 358.2852, 353.4254, 354.3373, 
    353.3712, 353.5013, 353.443, 352.7326, 352.3741, 351.6253, 351.7614, 
    352.3116, 353.5598, 353.1364, 354.2047, 354.1805, 355.3696, 354.8335, 
    356.8327, 356.2646, 357.9068, 357.4937, 357.8873, 357.768, 357.8888, 
    357.283, 357.5425, 357.0096, 354.9337, 355.5436, 353.7245, 352.6302, 
    351.9048, 351.3898, 351.4626, 351.6013, 352.3148, 352.9862, 353.4977, 
    353.8398, 354.1771, 355.1964, 355.7372, 356.9473, 356.7294, 357.0989, 
    357.4526, 358.0458, 357.9482, 358.2095, 357.0895, 357.8336, 356.6052, 
    356.9411, 354.2668, 353.2507, 352.8173, 352.4394, 351.5185, 352.1543, 
    351.9036, 352.5005, 352.8794, 352.6921, 353.8492, 353.3992, 355.7692, 
    354.7483, 357.4113, 356.7741, 357.5641, 357.1611, 357.8515, 357.2302, 
    358.3069, 358.5411, 358.381, 358.9966, 357.1957, 357.8871, 352.6867, 
    352.7173, 352.8598, 352.2332, 352.195, 351.6215, 352.132, 352.3492, 
    352.9016, 353.2278, 353.5382, 354.2208, 354.9828, 356.049, 356.8154, 
    357.3291, 357.0143, 357.2922, 356.9814, 356.8358, 358.4532, 357.5448, 
    358.9081, 358.8327, 358.2156, 358.8412, 352.7388, 352.5629, 351.9518, 
    352.4301, 351.5591, 352.0464, 352.3264, 353.4082, 353.6464, 353.8666, 
    354.3022, 354.8609, 355.841, 356.6941, 357.4733, 357.4162, 357.4363, 
    357.6101, 357.1792, 357.6809, 357.7649, 357.545, 358.8226, 358.4576, 
    358.8311, 358.5935, 352.6201, 352.9161, 352.7561, 353.0568, 352.8448, 
    353.7869, 354.0695, 355.3921, 354.8498, 355.7135, 354.9377, 355.075, 
    355.7408, 354.9797, 356.6467, 355.5157, 357.6169, 356.4867, 357.6877, 
    357.4699, 357.8307, 358.1536, 358.5602, 359.3098, 359.1363, 359.7635, 
    353.3575, 353.7412, 353.7078, 354.1097, 354.4069, 355.0515, 356.085, 
    355.6964, 356.4102, 356.5533, 355.4692, 356.1345, 353.9984, 354.343, 
    354.1381, 353.3875, 355.7855, 354.5545, 356.828, 356.1612, 358.1075, 
    357.1392, 359.0407, 359.8526, 360.6185, 361.5114, 353.9511, 353.6903, 
    354.1576, 354.8036, 355.404, 356.2018, 356.2836, 356.433, 356.8203, 
    357.1457, 356.4798, 357.2274, 354.4223, 355.8925, 353.5913, 354.2837, 
    354.7657, 354.5546, 355.6521, 355.9107, 356.9613, 356.4184, 359.6519, 
    358.2213, 362.1925, 361.0826, 353.5991, 353.9504, 355.1726, 354.5911, 
    356.2552, 356.6647, 356.9979, 357.4233, 357.4695, 357.7216, 357.3084, 
    357.7054, 356.2035, 356.8747, 355.0334, 355.4813, 355.2754, 355.0492, 
    355.7472, 356.4902, 356.5067, 356.7448, 357.4149, 356.262, 359.8354, 
    357.6275, 354.3334, 355.0094, 355.1067, 354.8447, 356.6236, 355.9789, 
    357.7155, 357.2463, 358.0152, 357.6331, 357.5768, 357.0861, 356.7805, 
    356.0084, 355.3804, 354.8828, 354.9985, 355.5452, 356.5358, 357.4734, 
    357.2679, 357.9568, 356.1346, 356.8983, 356.6029, 357.3733, 355.686, 
    357.1209, 355.319, 355.4771, 355.9662, 356.9497, 357.1682, 357.4005, 
    357.2573, 356.5611, 356.4473, 355.9544, 355.8181, 355.4427, 355.1317, 
    355.4157, 355.7139, 356.5616, 357.3253, 358.1581, 358.3622, 359.3337, 
    358.542, 359.8476, 358.7363, 360.6606, 357.205, 358.7048, 355.9886, 
    356.2814, 356.8103, 358.0246, 357.3697, 358.136, 356.4428, 355.5638, 
    355.3371, 354.9129, 355.3468, 355.3115, 355.7267, 355.5933, 356.5898, 
    356.0545, 357.5753, 358.1301, 359.6976, 360.6581, 361.6368, 362.0685, 
    362.2, 362.2549 ;

 FSH_R =
  351.6926, 352.5784, 352.4064, 353.1205, 352.7246, 353.192, 351.8725, 
    352.6134, 352.1405, 351.7727, 354.5061, 353.1524, 355.9149, 355.051, 
    357.222, 355.7801, 357.5129, 357.181, 358.1813, 357.8948, 359.173, 
    358.3136, 359.8365, 358.9681, 359.1037, 358.2852, 353.4254, 354.3373, 
    353.3712, 353.5013, 353.443, 352.7326, 352.3741, 351.6253, 351.7614, 
    352.3116, 353.5598, 353.1364, 354.2047, 354.1805, 355.3696, 354.8335, 
    356.8327, 356.2646, 357.9068, 357.4937, 357.8873, 357.768, 357.8888, 
    357.283, 357.5425, 357.0096, 354.9337, 355.5436, 353.7245, 352.6302, 
    351.9048, 351.3898, 351.4626, 351.6013, 352.3148, 352.9862, 353.4977, 
    353.8398, 354.1771, 355.1964, 355.7372, 356.9473, 356.7294, 357.0989, 
    357.4526, 358.0458, 357.9482, 358.2095, 357.0895, 357.8336, 356.6052, 
    356.9411, 354.2668, 353.2507, 352.8173, 352.4394, 351.5185, 352.1543, 
    351.9036, 352.5005, 352.8794, 352.6921, 353.8492, 353.3992, 355.7692, 
    354.7483, 357.4113, 356.7741, 357.5641, 357.1611, 357.8515, 357.2302, 
    358.3069, 358.5411, 358.381, 358.9966, 357.1957, 357.8871, 352.6867, 
    352.7173, 352.8598, 352.2332, 352.195, 351.6215, 352.132, 352.3492, 
    352.9016, 353.2278, 353.5382, 354.2208, 354.9828, 356.049, 356.8154, 
    357.3291, 357.0143, 357.2922, 356.9814, 356.8358, 358.4532, 357.5448, 
    358.9081, 358.8327, 358.2156, 358.8412, 352.7388, 352.5629, 351.9518, 
    352.4301, 351.5591, 352.0464, 352.3264, 353.4082, 353.6464, 353.8666, 
    354.3022, 354.8609, 355.841, 356.6941, 357.4733, 357.4162, 357.4363, 
    357.6101, 357.1792, 357.6809, 357.7649, 357.545, 358.8226, 358.4576, 
    358.8311, 358.5935, 352.6201, 352.9161, 352.7561, 353.0568, 352.8448, 
    353.7869, 354.0695, 355.3921, 354.8498, 355.7135, 354.9377, 355.075, 
    355.7408, 354.9797, 356.6467, 355.5157, 357.6169, 356.4867, 357.6877, 
    357.4699, 357.8307, 358.1536, 358.5602, 359.3098, 359.1363, 359.7635, 
    353.3575, 353.7412, 353.7078, 354.1097, 354.4069, 355.0515, 356.085, 
    355.6964, 356.4102, 356.5533, 355.4692, 356.1345, 353.9984, 354.343, 
    354.1381, 353.3875, 355.7855, 354.5545, 356.828, 356.1612, 358.1075, 
    357.1392, 359.0407, 359.8526, 360.6185, 361.5114, 353.9511, 353.6903, 
    354.1576, 354.8036, 355.404, 356.2018, 356.2836, 356.433, 356.8203, 
    357.1457, 356.4798, 357.2274, 354.4223, 355.8925, 353.5913, 354.2837, 
    354.7657, 354.5546, 355.6521, 355.9107, 356.9613, 356.4184, 359.6519, 
    358.2213, 362.1925, 361.0826, 353.5991, 353.9504, 355.1726, 354.5911, 
    356.2552, 356.6647, 356.9979, 357.4233, 357.4695, 357.7216, 357.3084, 
    357.7054, 356.2035, 356.8747, 355.0334, 355.4813, 355.2754, 355.0492, 
    355.7472, 356.4902, 356.5067, 356.7448, 357.4149, 356.262, 359.8354, 
    357.6275, 354.3334, 355.0094, 355.1067, 354.8447, 356.6236, 355.9789, 
    357.7155, 357.2463, 358.0152, 357.6331, 357.5768, 357.0861, 356.7805, 
    356.0084, 355.3804, 354.8828, 354.9985, 355.5452, 356.5358, 357.4734, 
    357.2679, 357.9568, 356.1346, 356.8983, 356.6029, 357.3733, 355.686, 
    357.1209, 355.319, 355.4771, 355.9662, 356.9497, 357.1682, 357.4005, 
    357.2573, 356.5611, 356.4473, 355.9544, 355.8181, 355.4427, 355.1317, 
    355.4157, 355.7139, 356.5616, 357.3253, 358.1581, 358.3622, 359.3337, 
    358.542, 359.8476, 358.7363, 360.6606, 357.205, 358.7048, 355.9886, 
    356.2814, 356.8103, 358.0246, 357.3697, 358.136, 356.4428, 355.5638, 
    355.3371, 354.9129, 355.3468, 355.3115, 355.7267, 355.5933, 356.5898, 
    356.0545, 357.5753, 358.1301, 359.6976, 360.6581, 361.6368, 362.0685, 
    362.2, 362.2549 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.659273, -6.65982, -6.659716, -6.660152, -6.659914, -6.660197, -6.659389, 
    -6.659838, -6.659554, -6.659329, -6.660985, -6.660172, -6.661876, 
    -6.661349, -6.662688, -6.661788, -6.662872, -6.662673, -6.663299, 
    -6.66312, -6.663899, -6.663382, -6.664322, -6.663782, -6.663862, 
    -6.663363, -6.660347, -6.66088, -6.660312, -6.660389, -6.660357, 
    -6.659915, -6.659686, -6.659239, -6.659322, -6.659655, -6.660424, 
    -6.66017, -6.660831, -6.660817, -6.661548, -6.661218, -6.662457, 
    -6.662107, -6.663128, -6.662869, -6.663114, -6.663041, -6.663115, 
    -6.662736, -6.662898, -6.662568, -6.661277, -6.661653, -6.660529, 
    -6.659838, -6.659407, -6.659092, -6.659137, -6.659219, -6.659656, 
    -6.660077, -6.660394, -6.660605, -6.660815, -6.66142, -6.661766, 
    -6.662522, -6.662395, -6.662617, -6.662844, -6.663212, -6.663153, 
    -6.663312, -6.662618, -6.663076, -6.66232, -6.662525, -6.660834, 
    -6.66024, -6.659956, -6.659735, -6.65917, -6.659558, -6.659404, 
    -6.659778, -6.66001, -6.659897, -6.660611, -6.660332, -6.661786, 
    -6.66116, -6.662817, -6.662421, -6.662914, -6.662664, -6.663089, 
    -6.662707, -6.663375, -6.663517, -6.663419, -6.663806, -6.662685, 
    -6.663111, -6.659892, -6.65991, -6.66, -6.659606, -6.659584, -6.659235, 
    -6.659549, -6.65968, -6.660027, -6.660225, -6.660417, -6.660838, 
    -6.661303, -6.661964, -6.662446, -6.662769, -6.662574, -6.662745, 
    -6.662552, -6.662463, -6.663461, -6.662897, -6.663751, -6.663704, 
    -6.663315, -6.66371, -6.659924, -6.659818, -6.659437, -6.659735, 
    -6.659197, -6.659493, -6.659661, -6.66033, -6.660486, -6.660619, 
    -6.66089, -6.661234, -6.661837, -6.662368, -6.662858, -6.662823, 
    -6.662836, -6.662941, -6.662674, -6.662986, -6.663034, -6.662901, 
    -6.663698, -6.663471, -6.663703, -6.663557, -6.659853, -6.660034, 
    -6.659935, -6.660118, -6.659986, -6.660562, -6.660734, -6.661552, 
    -6.661225, -6.661756, -6.661282, -6.661364, -6.661758, -6.66131, 
    -6.662331, -6.661625, -6.662946, -6.662224, -6.66299, -6.662857, 
    -6.663081, -6.663279, -6.663534, -6.663995, -6.66389, -6.664282, 
    -6.660306, -6.660538, -6.660524, -6.660771, -6.660952, -6.661354, 
    -6.661991, -6.661754, -6.662198, -6.662284, -6.661614, -6.662019, 
    -6.660698, -6.660903, -6.660786, -6.660321, -6.661799, -6.661035, 
    -6.662453, -6.66204, -6.663249, -6.66264, -6.66383, -6.664322, -6.664819, 
    -6.665362, -6.660671, -6.660513, -6.660802, -6.66119, -6.66157, 
    -6.662064, -6.662118, -6.662209, -6.662453, -6.662654, -6.662231, 
    -6.662705, -6.660937, -6.661868, -6.660448, -6.660865, -6.66117, 
    -6.661044, -6.661728, -6.661887, -6.662532, -6.662203, -6.664195, 
    -6.663311, -6.6658, -6.665097, -6.660457, -6.660674, -6.661422, 
    -6.661067, -6.662101, -6.662353, -6.662563, -6.662822, -6.662855, 
    -6.663009, -6.662756, -6.663002, -6.662065, -6.662484, -6.661345, 
    -6.661618, -6.661494, -6.661354, -6.661786, -6.662236, -6.662257, 
    -6.662399, -6.662781, -6.662105, -6.664288, -6.662919, -6.660911, 
    -6.661315, -6.661386, -6.661227, -6.662327, -6.661927, -6.663007, 
    -6.662717, -6.663195, -6.662957, -6.662921, -6.662617, -6.662425, 
    -6.661943, -6.661554, -6.661252, -6.661323, -6.661655, -6.662266, 
    -6.662853, -6.662723, -6.663159, -6.662025, -6.662494, -6.662309, 
    -6.662794, -6.661745, -6.662604, -6.661521, -6.661619, -6.661919, 
    -6.662519, -6.662668, -6.662808, -6.662724, -6.662283, -6.662217, 
    -6.661914, -6.661825, -6.661598, -6.661406, -6.661579, -6.661759, 
    -6.662289, -6.66276, -6.66328, -6.663411, -6.663991, -6.663504, 
    -6.664294, -6.663599, -6.664814, -6.662671, -6.663601, -6.661936, 
    -6.662118, -6.662435, -6.663187, -6.662792, -6.663259, -6.662215, 
    -6.661661, -6.661532, -6.661268, -6.661538, -6.661517, -6.661774, 
    -6.661692, -6.662306, -6.661977, -6.662917, -6.663258, -6.664237, 
    -6.664832, -6.665456, -6.665727, -6.66581, -6.665844 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.484155e-43, 0, 1.912772e-42, 
    3.629363e-43, 4.945042e-41, 1.242251e-41, 5.060599e-39, 9.290469e-41, 
    9.736725e-38, 1.98011e-39, 3.686572e-39, 8.117582e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.165713e-44, 2.802597e-45, 1.31652e-41, 
    1.734807e-42, 1.19825e-41, 6.695404e-42, 1.207219e-41, 6.067622e-43, 
    2.209848e-42, 1.527415e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.107026e-43, 3.643376e-44, 2.39622e-43, 1.41391e-42, 2.581612e-41, 
    1.610512e-41, 5.664469e-41, 2.284116e-43, 9.242965e-42, 1.961818e-44, 
    1.079e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.151867e-42, 
    4.624285e-44, 2.457878e-42, 3.279038e-43, 1.007954e-41, 4.652311e-43, 
    9.005024e-41, 2.726717e-40, 1.280843e-40, 2.25279e-39, 3.909623e-43, 
    1.19839e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    5.605194e-44, 7.637077e-43, 1.555441e-43, 6.347882e-43, 1.317221e-43, 
    6.305843e-44, 1.803401e-40, 2.237874e-42, 1.5001e-39, 1.059208e-39, 
    5.835567e-41, 1.101639e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.082857e-44, 1.566652e-42, 1.178492e-42, 1.303208e-42, 3.085659e-42, 
    3.601337e-43, 4.37065e-42, 6.605721e-42, 2.235071e-42, 1.01087e-39, 
    1.837845e-40, 1.051384e-39, 3.479578e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.382207e-44, 0, 3.190757e-42, 9.809089e-45, 4.519188e-42, 
    1.540027e-42, 9.090223e-42, 4.333936e-41, 2.977451e-40, 9.368527e-39, 
    4.266976e-39, 7.056501e-38, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 
    7.006492e-45, 1.401298e-44, 0, 1.401298e-45, 0, 0, 0, 0, 0, 0, 
    6.025583e-44, 1.401298e-45, 3.474379e-41, 2.942727e-43, 2.759103e-39, 
    1.047586e-37, 2.781373e-36, 1.085173e-34, 0, 0, 0, 0, 0, 2.802597e-45, 
    4.203895e-45, 8.407791e-45, 5.745324e-44, 3.040818e-43, 9.809089e-45, 
    4.582246e-43, 0, 0, 0, 0, 0, 0, 0, 0, 1.191104e-43, 7.006492e-45, 
    4.333622e-38, 6.009609e-41, 1.567935e-33, 1.911503e-35, 0, 0, 0, 0, 
    2.802597e-45, 2.662467e-44, 1.429324e-43, 1.223334e-42, 1.537224e-42, 
    5.338947e-42, 6.880375e-43, 4.926965e-42, 2.802597e-45, 7.707142e-44, 0, 
    0, 0, 0, 0, 9.809089e-45, 1.121039e-44, 3.923636e-44, 1.1869e-42, 
    2.802597e-45, 9.780159e-38, 3.396747e-42, 0, 0, 0, 0, 2.101948e-44, 0, 
    5.179199e-42, 5.044674e-43, 2.225822e-41, 3.454201e-42, 2.617626e-42, 
    2.242078e-43, 4.764415e-44, 1.401298e-45, 0, 0, 0, 0, 1.261169e-44, 
    1.569454e-42, 5.63322e-43, 1.677915e-41, 1.401298e-45, 8.68805e-44, 
    1.821688e-44, 9.52883e-43, 0, 2.704506e-43, 0, 0, 0, 1.121039e-43, 
    3.405155e-43, 1.091612e-42, 5.324934e-43, 1.541428e-44, 8.407791e-45, 0, 
    0, 0, 0, 0, 0, 1.541428e-44, 7.496947e-43, 4.430766e-41, 1.170028e-40, 
    1.048755e-38, 2.749264e-40, 1.032221e-37, 6.868086e-40, 3.346619e-36, 
    4.119817e-43, 5.894758e-40, 1.401298e-45, 2.802597e-45, 5.465064e-44, 
    2.339888e-41, 9.360674e-43, 3.99356e-41, 8.407791e-45, 0, 0, 0, 0, 0, 0, 
    0, 1.821688e-44, 1.401298e-45, 2.599409e-42, 3.878654e-41, 5.282891e-38, 
    3.295288e-36, 1.781647e-34, 9.699692e-34, 1.611632e-33, 1.990581e-33 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.203895e-45, 0, 3.623758e-42, 
    1.401298e-45, 1.547874e-41, 2.938523e-42, 4.000861e-40, 1.005025e-40, 
    4.094323e-38, 7.516579e-40, 7.877586e-37, 1.602027e-38, 2.982655e-38, 
    6.567662e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.988623e-43, 2.522337e-44, 1.065127e-40, 1.40312e-41, 9.694043e-41, 
    5.41728e-41, 9.767611e-41, 4.907347e-42, 1.788477e-41, 1.233143e-42, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 8.996336e-43, 
    2.928714e-43, 1.9422e-42, 1.14402e-41, 2.088705e-40, 1.302941e-40, 
    4.582919e-40, 1.848313e-42, 7.478029e-41, 1.541428e-43, 8.68805e-43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 9.318635e-42, 
    3.685415e-43, 1.988583e-41, 2.654059e-42, 8.154436e-41, 3.759684e-42, 
    7.285603e-40, 2.20608e-39, 1.036277e-39, 1.822641e-38, 3.161329e-42, 
    9.695304e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.407791e-45, 
    4.568233e-43, 6.174121e-42, 1.261169e-42, 5.132956e-42, 1.066388e-42, 
    5.058687e-43, 1.459064e-39, 1.810197e-41, 1.213669e-38, 8.569614e-39, 
    4.721325e-40, 8.912917e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.802597e-45, 2.438259e-43, 1.267054e-41, 9.538639e-42, 1.054337e-41, 
    2.496413e-41, 2.909096e-42, 3.536317e-41, 5.344132e-41, 1.808936e-41, 
    8.178537e-39, 1.48693e-39, 8.506322e-39, 2.815182e-39, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.401298e-45, 0, 0, 1.401298e-45, 0, 1.919779e-43, 0, 
    2.580912e-41, 8.407791e-44, 3.655848e-41, 1.246035e-41, 7.354435e-41, 
    3.506371e-40, 2.408934e-39, 7.579692e-38, 3.452236e-38, 5.709127e-37, 0, 
    0, 0, 0, 0, 0, 9.809089e-45, 1.401298e-45, 5.605194e-44, 1.177091e-43, 0, 
    1.261169e-44, 0, 0, 0, 0, 1.401298e-45, 0, 4.876519e-43, 1.541428e-44, 
    2.811019e-40, 2.383609e-42, 2.232277e-38, 8.47559e-37, 2.250295e-35, 
    8.779691e-34, 0, 0, 0, 0, 0, 1.821688e-44, 2.802597e-44, 6.305843e-44, 
    4.680337e-43, 2.456476e-42, 7.987401e-44, 3.706434e-42, 0, 4.203895e-45, 
    0, 0, 0, 0, 1.401298e-45, 4.203895e-45, 9.654946e-43, 5.745324e-44, 
    3.506156e-37, 4.862099e-40, 1.268552e-32, 1.546519e-34, 0, 0, 0, 0, 
    2.522337e-44, 2.101948e-43, 1.160275e-42, 9.898772e-42, 1.243793e-41, 
    4.319222e-41, 5.56876e-42, 3.986414e-41, 1.821688e-44, 6.179726e-43, 0, 
    0, 0, 0, 1.401298e-45, 8.547921e-44, 9.24857e-44, 3.180948e-43, 
    9.603098e-42, 2.522337e-44, 7.912726e-37, 2.748367e-41, 0, 0, 0, 0, 
    1.695571e-43, 5.605194e-45, 4.190723e-41, 4.076377e-42, 1.800823e-40, 
    2.794189e-41, 2.117502e-41, 1.816083e-42, 3.811532e-43, 7.006492e-45, 0, 
    0, 0, 0, 1.079e-43, 1.269997e-41, 4.555621e-42, 1.35755e-40, 
    1.261169e-44, 6.992479e-43, 1.527415e-43, 7.70574e-42, 1.401298e-45, 
    2.191631e-42, 0, 0, 5.605194e-45, 9.122453e-43, 2.75215e-42, 
    8.833786e-42, 4.307591e-42, 1.21913e-43, 6.726233e-44, 5.605194e-45, 
    2.802597e-45, 0, 0, 0, 1.401298e-45, 1.233143e-43, 6.069024e-42, 
    3.584746e-40, 9.46622e-40, 8.485051e-38, 2.224322e-39, 8.351273e-37, 
    5.556685e-39, 2.707612e-35, 3.33509e-42, 4.769207e-39, 5.605194e-45, 
    2.802597e-44, 4.456129e-43, 1.893126e-40, 7.568413e-42, 3.230974e-40, 
    6.586103e-44, 0, 0, 0, 0, 0, 1.401298e-45, 0, 1.415311e-43, 8.407791e-45, 
    2.103069e-41, 3.13811e-40, 4.274171e-37, 2.666083e-35, 1.441458e-33, 
    7.847624e-33, 1.303905e-32, 1.610498e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.809089e-45, 0, 4.063766e-44, 
    8.407791e-45, 1.067789e-42, 2.690493e-43, 1.093321e-40, 2.006659e-42, 
    2.103568e-39, 4.277884e-41, 7.9647e-41, 1.754426e-42, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 2.844636e-43, 
    3.783506e-44, 2.592402e-43, 1.443337e-43, 2.606415e-43, 1.261169e-44, 
    4.764415e-44, 2.802597e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.802597e-45, 1.401298e-45, 5.605194e-45, 3.082857e-44, 5.577168e-43, 
    3.47522e-43, 1.223334e-42, 5.605194e-45, 2.003857e-43, 0, 2.802597e-45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.522337e-44, 1.401298e-45, 
    5.324934e-44, 7.006492e-45, 2.172013e-43, 9.809089e-45, 1.945002e-42, 
    5.891059e-42, 2.767564e-42, 4.86699e-41, 8.407791e-45, 2.592402e-43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 1.681558e-44, 
    2.802597e-45, 1.401298e-44, 2.802597e-45, 1.401298e-45, 3.89561e-42, 
    4.764415e-44, 3.240923e-41, 2.28832e-41, 1.261169e-42, 2.379965e-41, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.363116e-44, 2.522337e-44, 
    2.802597e-44, 6.726233e-44, 8.407791e-45, 9.3887e-44, 1.429324e-43, 
    4.764415e-44, 2.183924e-41, 3.969879e-42, 2.271505e-41, 7.517966e-42, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.866362e-44, 0, 
    9.809089e-44, 3.363116e-44, 1.961818e-43, 9.360674e-43, 6.43196e-42, 
    2.024021e-40, 9.218582e-41, 1.524519e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 7.51096e-43, 7.006492e-45, 
    5.960843e-41, 2.263253e-39, 6.009009e-38, 2.344459e-36, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.401298e-45, 7.006492e-45, 0, 9.809089e-45, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.802597e-45, 0, 9.362551e-40, 1.299004e-42, 3.387443e-35, 
    4.129701e-37, 0, 0, 0, 0, 0, 0, 2.802597e-45, 2.662467e-44, 3.363116e-44, 
    1.149065e-43, 1.541428e-44, 1.064987e-43, 0, 1.401298e-45, 0, 0, 0, 0, 0, 
    0, 0, 1.401298e-45, 2.522337e-44, 0, 2.112951e-39, 7.286752e-44, 0, 0, 0, 
    0, 0, 0, 1.121039e-43, 1.121039e-44, 4.806454e-43, 7.426882e-44, 
    5.605194e-44, 4.203895e-45, 1.401298e-45, 0, 0, 0, 0, 0, 0, 3.363116e-44, 
    1.261169e-44, 3.629363e-43, 0, 1.401298e-45, 0, 2.101948e-44, 0, 
    5.605194e-45, 0, 0, 0, 2.802597e-45, 7.006492e-45, 2.382207e-44, 
    1.121039e-44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.681558e-44, 9.570869e-43, 
    2.527942e-42, 2.265773e-40, 5.940104e-42, 2.230057e-39, 1.483835e-41, 
    7.230192e-38, 8.407791e-45, 1.2735e-41, 0, 0, 1.401298e-45, 5.058687e-43, 
    1.961818e-44, 8.631999e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.605194e-44, 
    8.379765e-43, 1.141339e-39, 7.119295e-38, 3.849155e-36, 2.095568e-35, 
    3.481846e-35, 4.300548e-35 ;

 F_N2O_NIT =
  2.298666e-14, 2.318478e-14, 2.314619e-14, 2.330649e-14, 2.32175e-14, 
    2.332256e-14, 2.302674e-14, 2.319264e-14, 2.308666e-14, 2.300444e-14, 
    2.36192e-14, 2.331364e-14, 2.393886e-14, 2.374234e-14, 2.423762e-14, 
    2.390821e-14, 2.430433e-14, 2.422809e-14, 2.445794e-14, 2.439197e-14, 
    2.468719e-14, 2.448841e-14, 2.484097e-14, 2.463964e-14, 2.467107e-14, 
    2.448185e-14, 2.337499e-14, 2.358106e-14, 2.336281e-14, 2.339213e-14, 
    2.337896e-14, 2.321932e-14, 2.313908e-14, 2.297154e-14, 2.30019e-14, 
    2.312498e-14, 2.34053e-14, 2.330995e-14, 2.355065e-14, 2.35452e-14, 
    2.381466e-14, 2.369297e-14, 2.414829e-14, 2.401841e-14, 2.439472e-14, 
    2.429979e-14, 2.439025e-14, 2.43628e-14, 2.43906e-14, 2.425146e-14, 
    2.431101e-14, 2.418877e-14, 2.371576e-14, 2.385428e-14, 2.344239e-14, 
    2.319652e-14, 2.303399e-14, 2.291902e-14, 2.293525e-14, 2.296622e-14, 
    2.31257e-14, 2.327618e-14, 2.339121e-14, 2.346831e-14, 2.354441e-14, 
    2.377554e-14, 2.389837e-14, 2.417458e-14, 2.412462e-14, 2.42093e-14, 
    2.429035e-14, 2.442674e-14, 2.440427e-14, 2.446445e-14, 2.420705e-14, 
    2.437795e-14, 2.409616e-14, 2.417306e-14, 2.356511e-14, 2.333566e-14, 
    2.323846e-14, 2.315358e-14, 2.294773e-14, 2.308978e-14, 2.303372e-14, 
    2.316719e-14, 2.325221e-14, 2.321014e-14, 2.347041e-14, 2.336904e-14, 
    2.390565e-14, 2.367373e-14, 2.428089e-14, 2.413487e-14, 2.431596e-14, 
    2.422346e-14, 2.438205e-14, 2.423929e-14, 2.448687e-14, 2.454095e-14, 
    2.450398e-14, 2.464614e-14, 2.423137e-14, 2.439022e-14, 2.320898e-14, 
    2.321583e-14, 2.32478e-14, 2.310745e-14, 2.309887e-14, 2.297068e-14, 
    2.308473e-14, 2.313338e-14, 2.325714e-14, 2.33305e-14, 2.340035e-14, 
    2.355432e-14, 2.372689e-14, 2.396933e-14, 2.414431e-14, 2.426197e-14, 
    2.418979e-14, 2.425351e-14, 2.418228e-14, 2.414893e-14, 2.452067e-14, 
    2.431156e-14, 2.462566e-14, 2.460823e-14, 2.446586e-14, 2.461018e-14, 
    2.322064e-14, 2.318119e-14, 2.304446e-14, 2.315142e-14, 2.295674e-14, 
    2.30656e-14, 2.312831e-14, 2.337114e-14, 2.342468e-14, 2.347437e-14, 
    2.357268e-14, 2.369916e-14, 2.39219e-14, 2.41166e-14, 2.429506e-14, 
    2.428196e-14, 2.428657e-14, 2.432652e-14, 2.422761e-14, 2.434277e-14, 
    2.436212e-14, 2.431153e-14, 2.460588e-14, 2.45216e-14, 2.460785e-14, 
    2.455294e-14, 2.319401e-14, 2.326043e-14, 2.322452e-14, 2.329206e-14, 
    2.324446e-14, 2.345649e-14, 2.352026e-14, 2.381986e-14, 2.369667e-14, 
    2.38929e-14, 2.371656e-14, 2.374775e-14, 2.389929e-14, 2.372607e-14, 
    2.410582e-14, 2.3848e-14, 2.432807e-14, 2.406934e-14, 2.434432e-14, 
    2.429427e-14, 2.437716e-14, 2.445153e-14, 2.454526e-14, 2.47187e-14, 
    2.467848e-14, 2.48239e-14, 2.335964e-14, 2.344614e-14, 2.343852e-14, 
    2.352921e-14, 2.359639e-14, 2.374237e-14, 2.397747e-14, 2.388892e-14, 
    2.405162e-14, 2.408436e-14, 2.383721e-14, 2.398879e-14, 2.35041e-14, 
    2.358204e-14, 2.353562e-14, 2.336642e-14, 2.390928e-14, 2.362985e-14, 
    2.414718e-14, 2.39948e-14, 2.444091e-14, 2.42185e-14, 2.465635e-14, 
    2.484477e-14, 2.502282e-14, 2.523169e-14, 2.349342e-14, 2.343456e-14, 
    2.354e-14, 2.368628e-14, 2.382245e-14, 2.400411e-14, 2.402274e-14, 
    2.405686e-14, 2.414537e-14, 2.421992e-14, 2.406764e-14, 2.423863e-14, 
    2.360012e-14, 2.393361e-14, 2.341229e-14, 2.356863e-14, 2.367761e-14, 
    2.362977e-14, 2.387878e-14, 2.393766e-14, 2.417772e-14, 2.405347e-14, 
    2.479818e-14, 2.446723e-14, 2.539137e-14, 2.513129e-14, 2.341401e-14, 
    2.349321e-14, 2.376994e-14, 2.363806e-14, 2.401626e-14, 2.410983e-14, 
    2.418604e-14, 2.428364e-14, 2.429419e-14, 2.435213e-14, 2.425722e-14, 
    2.434837e-14, 2.400447e-14, 2.415783e-14, 2.37382e-14, 2.383997e-14, 
    2.379312e-14, 2.374178e-14, 2.390041e-14, 2.407e-14, 2.407364e-14, 
    2.412815e-14, 2.42821e-14, 2.401774e-14, 2.484103e-14, 2.433085e-14, 
    2.357973e-14, 2.373296e-14, 2.37549e-14, 2.369545e-14, 2.410043e-14, 
    2.395327e-14, 2.435072e-14, 2.424296e-14, 2.441964e-14, 2.433176e-14, 
    2.431884e-14, 2.420624e-14, 2.413627e-14, 2.395999e-14, 2.381705e-14, 
    2.370403e-14, 2.373028e-14, 2.385452e-14, 2.408039e-14, 2.429511e-14, 
    2.424798e-14, 2.440615e-14, 2.398867e-14, 2.416326e-14, 2.40957e-14, 
    2.427207e-14, 2.388656e-14, 2.421466e-14, 2.380306e-14, 2.3839e-14, 
    2.395035e-14, 2.417516e-14, 2.422506e-14, 2.427839e-14, 2.424547e-14, 
    2.408616e-14, 2.406011e-14, 2.394762e-14, 2.391661e-14, 2.383114e-14, 
    2.37605e-14, 2.382503e-14, 2.38929e-14, 2.408621e-14, 2.426111e-14, 
    2.445255e-14, 2.449953e-14, 2.472442e-14, 2.454125e-14, 2.484387e-14, 
    2.458644e-14, 2.503297e-14, 2.423375e-14, 2.457896e-14, 2.395543e-14, 
    2.40222e-14, 2.414321e-14, 2.442198e-14, 2.427128e-14, 2.444757e-14, 
    2.405909e-14, 2.385881e-14, 2.380714e-14, 2.371089e-14, 2.380934e-14, 
    2.380132e-14, 2.389572e-14, 2.386536e-14, 2.409263e-14, 2.397041e-14, 
    2.431847e-14, 2.444615e-14, 2.48086e-14, 2.503217e-14, 2.526086e-14, 
    2.536216e-14, 2.539303e-14, 2.540594e-14 ;

 F_NIT =
  3.83111e-11, 3.86413e-11, 3.857699e-11, 3.884415e-11, 3.869583e-11, 
    3.887093e-11, 3.837791e-11, 3.86544e-11, 3.847777e-11, 3.834074e-11, 
    3.936533e-11, 3.885606e-11, 3.98981e-11, 3.957057e-11, 4.039603e-11, 
    3.984702e-11, 4.050721e-11, 4.038015e-11, 4.076324e-11, 4.065329e-11, 
    4.114531e-11, 4.081402e-11, 4.140161e-11, 4.106607e-11, 4.111845e-11, 
    4.080309e-11, 3.895832e-11, 3.930177e-11, 3.893801e-11, 3.898688e-11, 
    3.896494e-11, 3.869887e-11, 3.856513e-11, 3.828589e-11, 3.83365e-11, 
    3.854164e-11, 3.900883e-11, 3.884991e-11, 3.925108e-11, 3.9242e-11, 
    3.96911e-11, 3.948828e-11, 4.024715e-11, 4.003069e-11, 4.065787e-11, 
    4.049965e-11, 4.065042e-11, 4.060466e-11, 4.0651e-11, 4.04191e-11, 
    4.051836e-11, 4.031462e-11, 3.952627e-11, 3.975713e-11, 3.907066e-11, 
    3.866087e-11, 3.838999e-11, 3.819836e-11, 3.822542e-11, 3.827702e-11, 
    3.854283e-11, 3.879364e-11, 3.898534e-11, 3.911384e-11, 3.924068e-11, 
    3.962589e-11, 3.983061e-11, 4.029098e-11, 4.02077e-11, 4.034883e-11, 
    4.048392e-11, 4.071124e-11, 4.067378e-11, 4.077408e-11, 4.034509e-11, 
    4.062992e-11, 4.016026e-11, 4.028843e-11, 3.927519e-11, 3.889277e-11, 
    3.873077e-11, 3.85893e-11, 3.824622e-11, 3.848297e-11, 3.838954e-11, 
    3.861199e-11, 3.875368e-11, 3.868356e-11, 3.911736e-11, 3.89484e-11, 
    3.984275e-11, 3.945622e-11, 4.046816e-11, 4.022477e-11, 4.052659e-11, 
    4.037244e-11, 4.063675e-11, 4.039882e-11, 4.081144e-11, 4.090158e-11, 
    4.083996e-11, 4.107691e-11, 4.038562e-11, 4.065036e-11, 3.868163e-11, 
    3.869306e-11, 3.874633e-11, 3.851241e-11, 3.849812e-11, 3.828447e-11, 
    3.847454e-11, 3.855563e-11, 3.87619e-11, 3.888416e-11, 3.900058e-11, 
    3.925719e-11, 3.954482e-11, 3.994888e-11, 4.024052e-11, 4.043663e-11, 
    4.031632e-11, 4.042251e-11, 4.03038e-11, 4.024821e-11, 4.086778e-11, 
    4.051927e-11, 4.104277e-11, 4.101371e-11, 4.077643e-11, 4.101697e-11, 
    3.870107e-11, 3.863531e-11, 3.840744e-11, 3.85857e-11, 3.826124e-11, 
    3.844267e-11, 3.854719e-11, 3.89519e-11, 3.904113e-11, 3.912395e-11, 
    3.928781e-11, 3.949861e-11, 3.986984e-11, 4.019433e-11, 4.049177e-11, 
    4.046993e-11, 4.047761e-11, 4.054419e-11, 4.037935e-11, 4.057128e-11, 
    4.060353e-11, 4.051922e-11, 4.100981e-11, 4.086933e-11, 4.101307e-11, 
    4.092158e-11, 3.865668e-11, 3.876738e-11, 3.870753e-11, 3.88201e-11, 
    3.874076e-11, 3.909415e-11, 3.920043e-11, 3.969977e-11, 3.949445e-11, 
    3.98215e-11, 3.95276e-11, 3.957959e-11, 3.983215e-11, 3.954344e-11, 
    4.017638e-11, 3.974666e-11, 4.054677e-11, 4.011556e-11, 4.057387e-11, 
    4.049044e-11, 4.06286e-11, 4.075255e-11, 4.090877e-11, 4.119784e-11, 
    4.11308e-11, 4.137317e-11, 3.893274e-11, 3.90769e-11, 3.90642e-11, 
    3.921535e-11, 3.932732e-11, 3.957062e-11, 3.996246e-11, 3.981487e-11, 
    4.008604e-11, 4.014059e-11, 3.972869e-11, 3.998131e-11, 3.91735e-11, 
    3.93034e-11, 3.922603e-11, 3.894403e-11, 3.984879e-11, 3.938309e-11, 
    4.024529e-11, 3.999133e-11, 4.073485e-11, 4.036417e-11, 4.109392e-11, 
    4.140795e-11, 4.170469e-11, 4.205282e-11, 3.91557e-11, 3.90576e-11, 
    3.923334e-11, 3.947714e-11, 3.970408e-11, 4.000685e-11, 4.003789e-11, 
    4.009476e-11, 4.024229e-11, 4.036654e-11, 4.011273e-11, 4.039771e-11, 
    3.933354e-11, 3.988936e-11, 3.902048e-11, 3.928104e-11, 3.946269e-11, 
    3.938296e-11, 3.979796e-11, 3.989609e-11, 4.02962e-11, 4.008911e-11, 
    4.13303e-11, 4.077871e-11, 4.231895e-11, 4.188549e-11, 3.902335e-11, 
    3.915535e-11, 3.961657e-11, 3.939677e-11, 4.00271e-11, 4.018305e-11, 
    4.031007e-11, 4.047274e-11, 4.049032e-11, 4.058688e-11, 4.04287e-11, 
    4.058062e-11, 4.000745e-11, 4.026305e-11, 3.956367e-11, 3.973329e-11, 
    3.965521e-11, 3.956964e-11, 3.983401e-11, 4.011666e-11, 4.012272e-11, 
    4.021358e-11, 4.047016e-11, 4.002958e-11, 4.140172e-11, 4.055142e-11, 
    3.929955e-11, 3.955493e-11, 3.95915e-11, 3.949241e-11, 4.016739e-11, 
    3.992212e-11, 4.058453e-11, 4.040494e-11, 4.06994e-11, 4.055293e-11, 
    4.053139e-11, 4.034374e-11, 4.022712e-11, 3.993331e-11, 3.969508e-11, 
    3.950672e-11, 3.955047e-11, 3.975753e-11, 4.013398e-11, 4.049184e-11, 
    4.04133e-11, 4.067692e-11, 3.998112e-11, 4.027211e-11, 4.015949e-11, 
    4.045345e-11, 3.981093e-11, 4.035776e-11, 3.967177e-11, 3.973166e-11, 
    3.991725e-11, 4.029194e-11, 4.03751e-11, 4.046398e-11, 4.040912e-11, 
    4.01436e-11, 4.010018e-11, 3.991271e-11, 3.986101e-11, 3.971858e-11, 
    3.960084e-11, 3.970839e-11, 3.982149e-11, 4.014368e-11, 4.043518e-11, 
    4.075426e-11, 4.083255e-11, 4.120736e-11, 4.090208e-11, 4.140646e-11, 
    4.09774e-11, 4.172163e-11, 4.038958e-11, 4.096494e-11, 3.992571e-11, 
    4.003699e-11, 4.023868e-11, 4.070329e-11, 4.045212e-11, 4.074595e-11, 
    4.009848e-11, 3.976468e-11, 3.967857e-11, 3.951815e-11, 3.968223e-11, 
    3.966888e-11, 3.982619e-11, 3.97756e-11, 4.015439e-11, 3.995068e-11, 
    4.053079e-11, 4.074358e-11, 4.134767e-11, 4.172029e-11, 4.210143e-11, 
    4.227026e-11, 4.232172e-11, 4.234324e-11 ;

 F_NIT_vr =
  2.423523e-10, 2.434402e-10, 2.432282e-10, 2.441063e-10, 2.436189e-10, 
    2.441935e-10, 2.425716e-10, 2.434815e-10, 2.429003e-10, 2.424482e-10, 
    2.458103e-10, 2.441434e-10, 2.475471e-10, 2.464806e-10, 2.491616e-10, 
    2.473802e-10, 2.49521e-10, 2.491099e-10, 2.503476e-10, 2.499924e-10, 
    2.515763e-10, 2.505107e-10, 2.523989e-10, 2.513215e-10, 2.514894e-10, 
    2.504742e-10, 2.444809e-10, 2.456044e-10, 2.444138e-10, 2.44574e-10, 
    2.445019e-10, 2.436277e-10, 2.431873e-10, 2.422671e-10, 2.424337e-10, 
    2.431096e-10, 2.446441e-10, 2.441226e-10, 2.454369e-10, 2.454073e-10, 
    2.468725e-10, 2.462113e-10, 2.486789e-10, 2.479764e-10, 2.50007e-10, 
    2.494953e-10, 2.499823e-10, 2.498342e-10, 2.499835e-10, 2.492339e-10, 
    2.495544e-10, 2.488953e-10, 2.463382e-10, 2.4709e-10, 2.448481e-10, 
    2.43502e-10, 2.426103e-10, 2.419781e-10, 2.420669e-10, 2.422372e-10, 
    2.43113e-10, 2.439376e-10, 2.445667e-10, 2.449874e-10, 2.454023e-10, 
    2.466591e-10, 2.473258e-10, 2.4882e-10, 2.485504e-10, 2.49007e-10, 
    2.494442e-10, 2.50178e-10, 2.500571e-10, 2.503802e-10, 2.489938e-10, 
    2.499146e-10, 2.483944e-10, 2.488098e-10, 2.455162e-10, 2.442644e-10, 
    2.437316e-10, 2.432664e-10, 2.421353e-10, 2.42916e-10, 2.426078e-10, 
    2.433403e-10, 2.438061e-10, 2.435753e-10, 2.449986e-10, 2.444444e-10, 
    2.473649e-10, 2.461056e-10, 2.493935e-10, 2.486051e-10, 2.495818e-10, 
    2.490833e-10, 2.49937e-10, 2.491681e-10, 2.505002e-10, 2.507906e-10, 
    2.505915e-10, 2.513545e-10, 2.491238e-10, 2.499795e-10, 2.435703e-10, 
    2.436079e-10, 2.437828e-10, 2.430126e-10, 2.429655e-10, 2.422608e-10, 
    2.428872e-10, 2.431542e-10, 2.438325e-10, 2.442335e-10, 2.44615e-10, 
    2.454553e-10, 2.463942e-10, 2.477093e-10, 2.486559e-10, 2.492905e-10, 
    2.48901e-10, 2.492444e-10, 2.488599e-10, 2.486795e-10, 2.506809e-10, 
    2.495562e-10, 2.51244e-10, 2.511506e-10, 2.503857e-10, 2.511604e-10, 
    2.436338e-10, 2.434172e-10, 2.426666e-10, 2.432535e-10, 2.421837e-10, 
    2.42782e-10, 2.431257e-10, 2.444553e-10, 2.447478e-10, 2.450191e-10, 
    2.45555e-10, 2.462431e-10, 2.474521e-10, 2.485054e-10, 2.494686e-10, 
    2.493976e-10, 2.494223e-10, 2.496371e-10, 2.491038e-10, 2.497241e-10, 
    2.498278e-10, 2.495556e-10, 2.511373e-10, 2.50685e-10, 2.511475e-10, 
    2.508526e-10, 2.434872e-10, 2.438507e-10, 2.436537e-10, 2.440235e-10, 
    2.437623e-10, 2.449215e-10, 2.45269e-10, 2.468988e-10, 2.462294e-10, 
    2.47295e-10, 2.463372e-10, 2.465067e-10, 2.473282e-10, 2.463883e-10, 
    2.484462e-10, 2.470493e-10, 2.496451e-10, 2.482476e-10, 2.497322e-10, 
    2.494622e-10, 2.499083e-10, 2.503083e-10, 2.508113e-10, 2.517409e-10, 
    2.515251e-10, 2.523033e-10, 2.443933e-10, 2.448652e-10, 2.448238e-10, 
    2.453182e-10, 2.45684e-10, 2.464784e-10, 2.477535e-10, 2.472733e-10, 
    2.481542e-10, 2.483312e-10, 2.46992e-10, 2.478134e-10, 2.45179e-10, 
    2.456033e-10, 2.453505e-10, 2.444263e-10, 2.473812e-10, 2.458627e-10, 
    2.486683e-10, 2.478439e-10, 2.502504e-10, 2.490524e-10, 2.514063e-10, 
    2.52414e-10, 2.533645e-10, 2.544747e-10, 2.451232e-10, 2.448017e-10, 
    2.453767e-10, 2.461729e-10, 2.469125e-10, 2.478973e-10, 2.479979e-10, 
    2.481821e-10, 2.486603e-10, 2.490627e-10, 2.482395e-10, 2.491629e-10, 
    2.457009e-10, 2.475131e-10, 2.446765e-10, 2.455292e-10, 2.461223e-10, 
    2.458622e-10, 2.472151e-10, 2.475338e-10, 2.488316e-10, 2.481605e-10, 
    2.521642e-10, 2.503903e-10, 2.553217e-10, 2.539407e-10, 2.446891e-10, 
    2.451211e-10, 2.466271e-10, 2.459101e-10, 2.479625e-10, 2.484685e-10, 
    2.488797e-10, 2.49406e-10, 2.494624e-10, 2.497745e-10, 2.492627e-10, 
    2.497539e-10, 2.478965e-10, 2.487258e-10, 2.464522e-10, 2.470043e-10, 
    2.467501e-10, 2.464707e-10, 2.473314e-10, 2.482493e-10, 2.482691e-10, 
    2.485631e-10, 2.493923e-10, 2.479658e-10, 2.523914e-10, 2.496543e-10, 
    2.455925e-10, 2.464255e-10, 2.465449e-10, 2.462218e-10, 2.48417e-10, 
    2.476207e-10, 2.497669e-10, 2.491859e-10, 2.501372e-10, 2.496642e-10, 
    2.49594e-10, 2.489871e-10, 2.486086e-10, 2.47655e-10, 2.468794e-10, 
    2.462656e-10, 2.464077e-10, 2.470822e-10, 2.483048e-10, 2.49464e-10, 
    2.492096e-10, 2.500614e-10, 2.478079e-10, 2.487518e-10, 2.483861e-10, 
    2.493385e-10, 2.472594e-10, 2.490329e-10, 2.468062e-10, 2.470008e-10, 
    2.476041e-10, 2.488196e-10, 2.490889e-10, 2.493763e-10, 2.491984e-10, 
    2.48338e-10, 2.48197e-10, 2.475878e-10, 2.474192e-10, 2.46956e-10, 
    2.465718e-10, 2.469222e-10, 2.472896e-10, 2.483364e-10, 2.492802e-10, 
    2.503106e-10, 2.505631e-10, 2.517676e-10, 2.507858e-10, 2.524052e-10, 
    2.510268e-10, 2.534142e-10, 2.491357e-10, 2.509928e-10, 2.476318e-10, 
    2.479929e-10, 2.486466e-10, 2.501486e-10, 2.493373e-10, 2.502861e-10, 
    2.481913e-10, 2.471057e-10, 2.468254e-10, 2.463024e-10, 2.468368e-10, 
    2.467934e-10, 2.473052e-10, 2.471402e-10, 2.483704e-10, 2.477093e-10, 
    2.495885e-10, 2.502755e-10, 2.522184e-10, 2.53411e-10, 2.546277e-10, 
    2.551647e-10, 2.553282e-10, 2.553963e-10,
  1.242928e-10, 1.252339e-10, 1.250507e-10, 1.258112e-10, 1.253892e-10, 
    1.258874e-10, 1.244835e-10, 1.252712e-10, 1.247681e-10, 1.243775e-10, 
    1.272916e-10, 1.258452e-10, 1.288015e-10, 1.278741e-10, 1.302087e-10, 
    1.286569e-10, 1.305225e-10, 1.301641e-10, 1.312445e-10, 1.309347e-10, 
    1.323197e-10, 1.313876e-10, 1.330401e-10, 1.32097e-10, 1.322443e-10, 
    1.313569e-10, 1.26136e-10, 1.271111e-10, 1.260782e-10, 1.262171e-10, 
    1.261548e-10, 1.253979e-10, 1.250169e-10, 1.242211e-10, 1.243655e-10, 
    1.249501e-10, 1.262796e-10, 1.258278e-10, 1.269679e-10, 1.269421e-10, 
    1.282156e-10, 1.276409e-10, 1.297886e-10, 1.291768e-10, 1.309476e-10, 
    1.305014e-10, 1.309266e-10, 1.307977e-10, 1.309283e-10, 1.302741e-10, 
    1.305542e-10, 1.299792e-10, 1.277484e-10, 1.284025e-10, 1.264553e-10, 
    1.252895e-10, 1.245179e-10, 1.239714e-10, 1.240486e-10, 1.241958e-10, 
    1.249535e-10, 1.256677e-10, 1.26213e-10, 1.265782e-10, 1.269384e-10, 
    1.280306e-10, 1.286106e-10, 1.299123e-10, 1.296772e-10, 1.300757e-10, 
    1.304571e-10, 1.31098e-10, 1.309925e-10, 1.312751e-10, 1.300653e-10, 
    1.308688e-10, 1.295433e-10, 1.299053e-10, 1.270357e-10, 1.259497e-10, 
    1.254885e-10, 1.250859e-10, 1.241079e-10, 1.247829e-10, 1.245167e-10, 
    1.251507e-10, 1.255541e-10, 1.253545e-10, 1.265882e-10, 1.26108e-10, 
    1.28645e-10, 1.275499e-10, 1.304126e-10, 1.297254e-10, 1.305775e-10, 
    1.301425e-10, 1.308881e-10, 1.30217e-10, 1.313804e-10, 1.316342e-10, 
    1.314607e-10, 1.321277e-10, 1.301798e-10, 1.309265e-10, 1.253489e-10, 
    1.253814e-10, 1.255331e-10, 1.248669e-10, 1.248262e-10, 1.242171e-10, 
    1.247591e-10, 1.249901e-10, 1.255775e-10, 1.259253e-10, 1.262563e-10, 
    1.269853e-10, 1.278011e-10, 1.289454e-10, 1.297699e-10, 1.303237e-10, 
    1.299841e-10, 1.302839e-10, 1.299487e-10, 1.297918e-10, 1.31539e-10, 
    1.305568e-10, 1.320317e-10, 1.3195e-10, 1.312818e-10, 1.319592e-10, 
    1.254043e-10, 1.252171e-10, 1.245678e-10, 1.250758e-10, 1.241509e-10, 
    1.246682e-10, 1.24966e-10, 1.261179e-10, 1.263716e-10, 1.266069e-10, 
    1.270722e-10, 1.276702e-10, 1.287218e-10, 1.296394e-10, 1.304793e-10, 
    1.304177e-10, 1.304394e-10, 1.306272e-10, 1.301621e-10, 1.307036e-10, 
    1.307945e-10, 1.305568e-10, 1.31939e-10, 1.315436e-10, 1.319482e-10, 
    1.316907e-10, 1.252779e-10, 1.255931e-10, 1.254227e-10, 1.257431e-10, 
    1.255173e-10, 1.265221e-10, 1.26824e-10, 1.282402e-10, 1.276584e-10, 
    1.285849e-10, 1.277525e-10, 1.278998e-10, 1.286149e-10, 1.277975e-10, 
    1.295886e-10, 1.28373e-10, 1.306345e-10, 1.294166e-10, 1.307109e-10, 
    1.304757e-10, 1.308653e-10, 1.312146e-10, 1.316546e-10, 1.324678e-10, 
    1.322793e-10, 1.329605e-10, 1.260635e-10, 1.264732e-10, 1.264372e-10, 
    1.268665e-10, 1.271843e-10, 1.278744e-10, 1.289839e-10, 1.285663e-10, 
    1.293334e-10, 1.294876e-10, 1.283223e-10, 1.290372e-10, 1.267477e-10, 
    1.271164e-10, 1.26897e-10, 1.260957e-10, 1.286623e-10, 1.273426e-10, 
    1.297835e-10, 1.290657e-10, 1.311648e-10, 1.301192e-10, 1.321756e-10, 
    1.33058e-10, 1.338909e-10, 1.34866e-10, 1.266971e-10, 1.264185e-10, 
    1.269176e-10, 1.276092e-10, 1.282525e-10, 1.291094e-10, 1.291973e-10, 
    1.293581e-10, 1.29775e-10, 1.301259e-10, 1.294088e-10, 1.302139e-10, 
    1.272017e-10, 1.287771e-10, 1.263131e-10, 1.27053e-10, 1.275685e-10, 
    1.273424e-10, 1.285186e-10, 1.287964e-10, 1.299273e-10, 1.293423e-10, 
    1.328399e-10, 1.312882e-10, 1.356106e-10, 1.343975e-10, 1.263211e-10, 
    1.266962e-10, 1.280046e-10, 1.273814e-10, 1.291668e-10, 1.296076e-10, 
    1.299665e-10, 1.304255e-10, 1.304753e-10, 1.307476e-10, 1.303014e-10, 
    1.3073e-10, 1.291113e-10, 1.298338e-10, 1.278549e-10, 1.283354e-10, 
    1.281143e-10, 1.278719e-10, 1.286207e-10, 1.2942e-10, 1.294374e-10, 
    1.29694e-10, 1.304179e-10, 1.291741e-10, 1.330402e-10, 1.306473e-10, 
    1.271056e-10, 1.278298e-10, 1.279336e-10, 1.276528e-10, 1.295634e-10, 
    1.288699e-10, 1.30741e-10, 1.302344e-10, 1.310649e-10, 1.306519e-10, 
    1.305912e-10, 1.300616e-10, 1.297323e-10, 1.289016e-10, 1.282272e-10, 
    1.276935e-10, 1.278176e-10, 1.284041e-10, 1.29469e-10, 1.304797e-10, 
    1.30258e-10, 1.310017e-10, 1.29037e-10, 1.298594e-10, 1.295413e-10, 
    1.303715e-10, 1.285552e-10, 1.301006e-10, 1.281611e-10, 1.283308e-10, 
    1.288561e-10, 1.299151e-10, 1.301502e-10, 1.304009e-10, 1.302462e-10, 
    1.294962e-10, 1.293735e-10, 1.288434e-10, 1.286971e-10, 1.282939e-10, 
    1.279603e-10, 1.28265e-10, 1.285852e-10, 1.294966e-10, 1.303198e-10, 
    1.312195e-10, 1.314402e-10, 1.324944e-10, 1.316357e-10, 1.330535e-10, 
    1.318473e-10, 1.339381e-10, 1.301907e-10, 1.318123e-10, 1.288801e-10, 
    1.291949e-10, 1.297647e-10, 1.310756e-10, 1.303676e-10, 1.311959e-10, 
    1.293688e-10, 1.284242e-10, 1.281805e-10, 1.277259e-10, 1.28191e-10, 
    1.281531e-10, 1.285986e-10, 1.284554e-10, 1.295269e-10, 1.289509e-10, 
    1.305896e-10, 1.311894e-10, 1.32889e-10, 1.339346e-10, 1.350024e-10, 
    1.354747e-10, 1.356185e-10, 1.356787e-10,
  1.174375e-10, 1.184788e-10, 1.182761e-10, 1.191182e-10, 1.186508e-10, 
    1.192026e-10, 1.176483e-10, 1.185202e-10, 1.179633e-10, 1.175311e-10, 
    1.207595e-10, 1.191558e-10, 1.224355e-10, 1.214055e-10, 1.239999e-10, 
    1.222749e-10, 1.24349e-10, 1.239502e-10, 1.251526e-10, 1.248076e-10, 
    1.263507e-10, 1.253119e-10, 1.271538e-10, 1.261023e-10, 1.262665e-10, 
    1.252777e-10, 1.194779e-10, 1.205593e-10, 1.19414e-10, 1.195679e-10, 
    1.194988e-10, 1.186604e-10, 1.182387e-10, 1.173581e-10, 1.175178e-10, 
    1.181647e-10, 1.196371e-10, 1.191365e-10, 1.204001e-10, 1.203715e-10, 
    1.217847e-10, 1.211467e-10, 1.235325e-10, 1.228524e-10, 1.24822e-10, 
    1.243254e-10, 1.247987e-10, 1.246551e-10, 1.248005e-10, 1.240726e-10, 
    1.243842e-10, 1.237445e-10, 1.21266e-10, 1.219922e-10, 1.198318e-10, 
    1.185405e-10, 1.176865e-10, 1.170819e-10, 1.171673e-10, 1.173301e-10, 
    1.181685e-10, 1.189592e-10, 1.195632e-10, 1.19968e-10, 1.203674e-10, 
    1.215795e-10, 1.222234e-10, 1.236701e-10, 1.234086e-10, 1.238518e-10, 
    1.242761e-10, 1.249895e-10, 1.24872e-10, 1.251867e-10, 1.238402e-10, 
    1.247344e-10, 1.232597e-10, 1.236623e-10, 1.204757e-10, 1.192715e-10, 
    1.187609e-10, 1.18315e-10, 1.17233e-10, 1.179797e-10, 1.176851e-10, 
    1.183866e-10, 1.188333e-10, 1.186123e-10, 1.199791e-10, 1.194469e-10, 
    1.222616e-10, 1.210458e-10, 1.242266e-10, 1.234623e-10, 1.244101e-10, 
    1.239261e-10, 1.247558e-10, 1.24009e-10, 1.25304e-10, 1.255867e-10, 
    1.253934e-10, 1.261365e-10, 1.239676e-10, 1.247986e-10, 1.186061e-10, 
    1.186421e-10, 1.188101e-10, 1.180726e-10, 1.180276e-10, 1.173537e-10, 
    1.179533e-10, 1.182089e-10, 1.188592e-10, 1.192445e-10, 1.196113e-10, 
    1.204194e-10, 1.213246e-10, 1.225953e-10, 1.235118e-10, 1.241276e-10, 
    1.237499e-10, 1.240834e-10, 1.237106e-10, 1.23536e-10, 1.254807e-10, 
    1.243871e-10, 1.260295e-10, 1.259384e-10, 1.251942e-10, 1.259487e-10, 
    1.186674e-10, 1.184602e-10, 1.177416e-10, 1.183038e-10, 1.172804e-10, 
    1.178527e-10, 1.181823e-10, 1.194579e-10, 1.197391e-10, 1.199999e-10, 
    1.205158e-10, 1.211793e-10, 1.223469e-10, 1.233667e-10, 1.243008e-10, 
    1.242322e-10, 1.242564e-10, 1.244654e-10, 1.239479e-10, 1.245504e-10, 
    1.246517e-10, 1.24387e-10, 1.259262e-10, 1.254857e-10, 1.259365e-10, 
    1.256496e-10, 1.185275e-10, 1.188765e-10, 1.186879e-10, 1.190427e-10, 
    1.187926e-10, 1.19906e-10, 1.202407e-10, 1.21812e-10, 1.211662e-10, 
    1.221949e-10, 1.212705e-10, 1.214341e-10, 1.222283e-10, 1.213204e-10, 
    1.233103e-10, 1.219596e-10, 1.244735e-10, 1.231192e-10, 1.245586e-10, 
    1.242967e-10, 1.247304e-10, 1.251193e-10, 1.256094e-10, 1.265156e-10, 
    1.263055e-10, 1.27065e-10, 1.193976e-10, 1.198516e-10, 1.198117e-10, 
    1.202877e-10, 1.206402e-10, 1.214058e-10, 1.22638e-10, 1.221741e-10, 
    1.230265e-10, 1.231979e-10, 1.219031e-10, 1.226973e-10, 1.20156e-10, 
    1.20565e-10, 1.203215e-10, 1.194333e-10, 1.222808e-10, 1.208159e-10, 
    1.235269e-10, 1.22729e-10, 1.250638e-10, 1.239003e-10, 1.261899e-10, 
    1.271739e-10, 1.281032e-10, 1.291924e-10, 1.200999e-10, 1.19791e-10, 
    1.203444e-10, 1.211117e-10, 1.218257e-10, 1.227776e-10, 1.228752e-10, 
    1.230539e-10, 1.235174e-10, 1.239076e-10, 1.231103e-10, 1.240055e-10, 
    1.206598e-10, 1.224083e-10, 1.196742e-10, 1.204946e-10, 1.210664e-10, 
    1.208155e-10, 1.221211e-10, 1.224297e-10, 1.236869e-10, 1.230363e-10, 
    1.269307e-10, 1.252014e-10, 1.300245e-10, 1.28669e-10, 1.196831e-10, 
    1.200988e-10, 1.215504e-10, 1.208588e-10, 1.228413e-10, 1.233313e-10, 
    1.237303e-10, 1.24241e-10, 1.242963e-10, 1.245994e-10, 1.241029e-10, 
    1.245798e-10, 1.227796e-10, 1.235827e-10, 1.213842e-10, 1.219177e-10, 
    1.216722e-10, 1.21403e-10, 1.222345e-10, 1.231228e-10, 1.23142e-10, 
    1.234274e-10, 1.24233e-10, 1.228493e-10, 1.271543e-10, 1.244881e-10, 
    1.205529e-10, 1.213565e-10, 1.214716e-10, 1.211599e-10, 1.232821e-10, 
    1.225113e-10, 1.24592e-10, 1.240283e-10, 1.249526e-10, 1.244929e-10, 
    1.244253e-10, 1.238361e-10, 1.234699e-10, 1.225466e-10, 1.217976e-10, 
    1.212051e-10, 1.213428e-10, 1.21994e-10, 1.231773e-10, 1.243012e-10, 
    1.240547e-10, 1.248822e-10, 1.22697e-10, 1.236113e-10, 1.232576e-10, 
    1.241808e-10, 1.221617e-10, 1.238798e-10, 1.217241e-10, 1.219125e-10, 
    1.224961e-10, 1.236733e-10, 1.239346e-10, 1.242136e-10, 1.240414e-10, 
    1.232074e-10, 1.230711e-10, 1.224819e-10, 1.223194e-10, 1.218715e-10, 
    1.215012e-10, 1.218395e-10, 1.221952e-10, 1.232078e-10, 1.241234e-10, 
    1.251249e-10, 1.253705e-10, 1.265455e-10, 1.255885e-10, 1.271692e-10, 
    1.258245e-10, 1.281562e-10, 1.239799e-10, 1.257853e-10, 1.225227e-10, 
    1.228725e-10, 1.235061e-10, 1.249647e-10, 1.241765e-10, 1.250986e-10, 
    1.230657e-10, 1.220164e-10, 1.217457e-10, 1.212411e-10, 1.217573e-10, 
    1.217152e-10, 1.2221e-10, 1.220509e-10, 1.232415e-10, 1.226014e-10, 
    1.244236e-10, 1.250913e-10, 1.269853e-10, 1.281521e-10, 1.293446e-10, 
    1.298725e-10, 1.300333e-10, 1.301006e-10,
  1.205486e-10, 1.216954e-10, 1.21472e-10, 1.223999e-10, 1.218848e-10, 
    1.22493e-10, 1.207807e-10, 1.21741e-10, 1.211275e-10, 1.206517e-10, 
    1.242104e-10, 1.224414e-10, 1.260611e-10, 1.249233e-10, 1.27791e-10, 
    1.258837e-10, 1.281773e-10, 1.277359e-10, 1.290669e-10, 1.286849e-10, 
    1.303945e-10, 1.292434e-10, 1.31285e-10, 1.301191e-10, 1.303012e-10, 
    1.292055e-10, 1.227965e-10, 1.239895e-10, 1.22726e-10, 1.228957e-10, 
    1.228195e-10, 1.218954e-10, 1.21431e-10, 1.204612e-10, 1.20637e-10, 
    1.213494e-10, 1.22972e-10, 1.224201e-10, 1.238136e-10, 1.23782e-10, 
    1.253421e-10, 1.246375e-10, 1.272738e-10, 1.265218e-10, 1.287008e-10, 
    1.281511e-10, 1.28675e-10, 1.28516e-10, 1.28677e-10, 1.278713e-10, 
    1.282162e-10, 1.275084e-10, 1.247693e-10, 1.255713e-10, 1.231867e-10, 
    1.217635e-10, 1.208227e-10, 1.201573e-10, 1.202512e-10, 1.204305e-10, 
    1.213536e-10, 1.222247e-10, 1.228905e-10, 1.233369e-10, 1.237775e-10, 
    1.251156e-10, 1.258268e-10, 1.274261e-10, 1.271368e-10, 1.276272e-10, 
    1.280965e-10, 1.288863e-10, 1.287562e-10, 1.291047e-10, 1.276143e-10, 
    1.286039e-10, 1.269722e-10, 1.274174e-10, 1.238972e-10, 1.225689e-10, 
    1.220063e-10, 1.215149e-10, 1.203235e-10, 1.211457e-10, 1.208212e-10, 
    1.215938e-10, 1.220859e-10, 1.218424e-10, 1.233491e-10, 1.227623e-10, 
    1.25869e-10, 1.245262e-10, 1.280417e-10, 1.271962e-10, 1.282448e-10, 
    1.277092e-10, 1.286276e-10, 1.278009e-10, 1.292345e-10, 1.295477e-10, 
    1.293337e-10, 1.301569e-10, 1.277552e-10, 1.286749e-10, 1.218356e-10, 
    1.218753e-10, 1.220603e-10, 1.21248e-10, 1.211983e-10, 1.204564e-10, 
    1.211165e-10, 1.213981e-10, 1.221145e-10, 1.225392e-10, 1.229435e-10, 
    1.238349e-10, 1.24834e-10, 1.262377e-10, 1.272509e-10, 1.279322e-10, 
    1.275143e-10, 1.278832e-10, 1.274708e-10, 1.272777e-10, 1.294303e-10, 
    1.282194e-10, 1.300384e-10, 1.299374e-10, 1.29113e-10, 1.299488e-10, 
    1.219032e-10, 1.216748e-10, 1.208834e-10, 1.215025e-10, 1.203757e-10, 
    1.210058e-10, 1.213688e-10, 1.227745e-10, 1.230844e-10, 1.233721e-10, 
    1.239412e-10, 1.246735e-10, 1.259632e-10, 1.270905e-10, 1.281238e-10, 
    1.28048e-10, 1.280747e-10, 1.28306e-10, 1.277334e-10, 1.284002e-10, 
    1.285122e-10, 1.282193e-10, 1.299239e-10, 1.294358e-10, 1.299352e-10, 
    1.296173e-10, 1.21749e-10, 1.221335e-10, 1.219257e-10, 1.223167e-10, 
    1.220411e-10, 1.232686e-10, 1.236378e-10, 1.253723e-10, 1.246591e-10, 
    1.257952e-10, 1.247743e-10, 1.249549e-10, 1.258323e-10, 1.248294e-10, 
    1.270282e-10, 1.255354e-10, 1.28315e-10, 1.268169e-10, 1.284092e-10, 
    1.281194e-10, 1.285994e-10, 1.290301e-10, 1.295729e-10, 1.305772e-10, 
    1.303443e-10, 1.311865e-10, 1.227079e-10, 1.232086e-10, 1.231645e-10, 
    1.236895e-10, 1.240785e-10, 1.249236e-10, 1.262849e-10, 1.257722e-10, 
    1.267143e-10, 1.269038e-10, 1.254729e-10, 1.263505e-10, 1.235443e-10, 
    1.239956e-10, 1.237268e-10, 1.227473e-10, 1.258902e-10, 1.242724e-10, 
    1.272677e-10, 1.263854e-10, 1.289686e-10, 1.276808e-10, 1.302162e-10, 
    1.313073e-10, 1.323384e-10, 1.335481e-10, 1.234823e-10, 1.231416e-10, 
    1.237521e-10, 1.24599e-10, 1.253873e-10, 1.264391e-10, 1.26547e-10, 
    1.267446e-10, 1.272571e-10, 1.276888e-10, 1.268071e-10, 1.277971e-10, 
    1.241003e-10, 1.260311e-10, 1.230129e-10, 1.23918e-10, 1.24549e-10, 
    1.24272e-10, 1.257136e-10, 1.260546e-10, 1.274446e-10, 1.267252e-10, 
    1.310376e-10, 1.291211e-10, 1.344728e-10, 1.329667e-10, 1.230227e-10, 
    1.234812e-10, 1.250833e-10, 1.243198e-10, 1.265095e-10, 1.270513e-10, 
    1.274926e-10, 1.280578e-10, 1.281189e-10, 1.284544e-10, 1.279048e-10, 
    1.284327e-10, 1.264414e-10, 1.273294e-10, 1.248997e-10, 1.25489e-10, 
    1.252178e-10, 1.249205e-10, 1.25839e-10, 1.268209e-10, 1.26842e-10, 
    1.271576e-10, 1.280491e-10, 1.265184e-10, 1.312859e-10, 1.283315e-10, 
    1.239821e-10, 1.248693e-10, 1.249963e-10, 1.246521e-10, 1.26997e-10, 
    1.261449e-10, 1.284462e-10, 1.278223e-10, 1.288454e-10, 1.283365e-10, 
    1.282617e-10, 1.276097e-10, 1.272046e-10, 1.261839e-10, 1.253563e-10, 
    1.24702e-10, 1.24854e-10, 1.255733e-10, 1.268811e-10, 1.281244e-10, 
    1.278515e-10, 1.287675e-10, 1.263501e-10, 1.273611e-10, 1.269699e-10, 
    1.279911e-10, 1.257586e-10, 1.276584e-10, 1.252752e-10, 1.254832e-10, 
    1.26128e-10, 1.274297e-10, 1.277187e-10, 1.280274e-10, 1.278369e-10, 
    1.269144e-10, 1.267636e-10, 1.261123e-10, 1.259328e-10, 1.254379e-10, 
    1.250289e-10, 1.254026e-10, 1.257955e-10, 1.269148e-10, 1.279276e-10, 
    1.290362e-10, 1.293082e-10, 1.306106e-10, 1.295499e-10, 1.313024e-10, 
    1.298116e-10, 1.323975e-10, 1.27769e-10, 1.29768e-10, 1.261574e-10, 
    1.26544e-10, 1.272447e-10, 1.28859e-10, 1.279863e-10, 1.290072e-10, 
    1.267577e-10, 1.255981e-10, 1.25299e-10, 1.247417e-10, 1.253117e-10, 
    1.252653e-10, 1.258118e-10, 1.256361e-10, 1.269521e-10, 1.262444e-10, 
    1.282598e-10, 1.289991e-10, 1.310981e-10, 1.323928e-10, 1.337172e-10, 
    1.343038e-10, 1.344826e-10, 1.345574e-10,
  1.31568e-10, 1.327968e-10, 1.325574e-10, 1.335523e-10, 1.329999e-10, 
    1.336521e-10, 1.318166e-10, 1.328457e-10, 1.321882e-10, 1.316784e-10, 
    1.354953e-10, 1.335968e-10, 1.374836e-10, 1.362607e-10, 1.393446e-10, 
    1.372929e-10, 1.397604e-10, 1.392851e-10, 1.407185e-10, 1.40307e-10, 
    1.421497e-10, 1.409086e-10, 1.431104e-10, 1.418527e-10, 1.420491e-10, 
    1.408678e-10, 1.339775e-10, 1.352581e-10, 1.339019e-10, 1.34084e-10, 
    1.340023e-10, 1.330113e-10, 1.325135e-10, 1.314744e-10, 1.316627e-10, 
    1.32426e-10, 1.341659e-10, 1.335738e-10, 1.350689e-10, 1.350351e-10, 
    1.367106e-10, 1.359537e-10, 1.387879e-10, 1.379789e-10, 1.403241e-10, 
    1.397322e-10, 1.402963e-10, 1.401251e-10, 1.402985e-10, 1.394309e-10, 
    1.398023e-10, 1.390402e-10, 1.360953e-10, 1.36957e-10, 1.343962e-10, 
    1.3287e-10, 1.318617e-10, 1.311489e-10, 1.312495e-10, 1.314415e-10, 
    1.324305e-10, 1.333643e-10, 1.340784e-10, 1.345573e-10, 1.350302e-10, 
    1.364674e-10, 1.372317e-10, 1.389518e-10, 1.386404e-10, 1.391682e-10, 
    1.396734e-10, 1.40524e-10, 1.403838e-10, 1.407593e-10, 1.391542e-10, 
    1.402198e-10, 1.384633e-10, 1.389424e-10, 1.35159e-10, 1.337334e-10, 
    1.331302e-10, 1.326034e-10, 1.313269e-10, 1.322077e-10, 1.318601e-10, 
    1.326879e-10, 1.332155e-10, 1.329544e-10, 1.345704e-10, 1.339408e-10, 
    1.37277e-10, 1.358342e-10, 1.396144e-10, 1.387043e-10, 1.39833e-10, 
    1.392564e-10, 1.402453e-10, 1.393551e-10, 1.408992e-10, 1.412367e-10, 
    1.41006e-10, 1.418934e-10, 1.393059e-10, 1.402963e-10, 1.329471e-10, 
    1.329896e-10, 1.33188e-10, 1.323173e-10, 1.322641e-10, 1.314692e-10, 
    1.321764e-10, 1.324782e-10, 1.332461e-10, 1.337015e-10, 1.341353e-10, 
    1.350919e-10, 1.361648e-10, 1.376734e-10, 1.387632e-10, 1.394965e-10, 
    1.390466e-10, 1.394437e-10, 1.389998e-10, 1.38792e-10, 1.411102e-10, 
    1.398058e-10, 1.417656e-10, 1.416567e-10, 1.407682e-10, 1.41669e-10, 
    1.330195e-10, 1.327747e-10, 1.319267e-10, 1.325901e-10, 1.313828e-10, 
    1.320578e-10, 1.324468e-10, 1.33954e-10, 1.342864e-10, 1.345951e-10, 
    1.35206e-10, 1.359924e-10, 1.373782e-10, 1.385906e-10, 1.397028e-10, 
    1.396211e-10, 1.396499e-10, 1.39899e-10, 1.392824e-10, 1.400003e-10, 
    1.401211e-10, 1.398056e-10, 1.416421e-10, 1.41116e-10, 1.416544e-10, 
    1.413117e-10, 1.328542e-10, 1.332665e-10, 1.330436e-10, 1.334629e-10, 
    1.331675e-10, 1.344841e-10, 1.348803e-10, 1.367432e-10, 1.359769e-10, 
    1.371977e-10, 1.361006e-10, 1.362946e-10, 1.372377e-10, 1.361597e-10, 
    1.385236e-10, 1.369184e-10, 1.399087e-10, 1.382965e-10, 1.400101e-10, 
    1.396979e-10, 1.402149e-10, 1.406788e-10, 1.412638e-10, 1.423468e-10, 
    1.420956e-10, 1.43004e-10, 1.338825e-10, 1.344197e-10, 1.343724e-10, 
    1.349358e-10, 1.353534e-10, 1.36261e-10, 1.377241e-10, 1.371729e-10, 
    1.381858e-10, 1.383897e-10, 1.368511e-10, 1.377946e-10, 1.3478e-10, 
    1.352645e-10, 1.349759e-10, 1.339248e-10, 1.372998e-10, 1.355617e-10, 
    1.387813e-10, 1.378322e-10, 1.406126e-10, 1.392259e-10, 1.419574e-10, 
    1.431346e-10, 1.442477e-10, 1.45555e-10, 1.347134e-10, 1.343478e-10, 
    1.350029e-10, 1.359123e-10, 1.367593e-10, 1.378899e-10, 1.380059e-10, 
    1.382185e-10, 1.387699e-10, 1.392344e-10, 1.382857e-10, 1.39351e-10, 
    1.35377e-10, 1.374513e-10, 1.342097e-10, 1.351812e-10, 1.358586e-10, 
    1.355612e-10, 1.371099e-10, 1.374764e-10, 1.389717e-10, 1.381976e-10, 
    1.428436e-10, 1.40777e-10, 1.46555e-10, 1.449265e-10, 1.342202e-10, 
    1.347122e-10, 1.364327e-10, 1.356125e-10, 1.379656e-10, 1.385485e-10, 
    1.390233e-10, 1.396317e-10, 1.396974e-10, 1.400587e-10, 1.39467e-10, 
    1.400353e-10, 1.378924e-10, 1.388476e-10, 1.362353e-10, 1.368685e-10, 
    1.36577e-10, 1.362577e-10, 1.372446e-10, 1.383006e-10, 1.383232e-10, 
    1.386629e-10, 1.396227e-10, 1.379752e-10, 1.431117e-10, 1.399267e-10, 
    1.352499e-10, 1.362027e-10, 1.363391e-10, 1.359693e-10, 1.3849e-10, 
    1.375735e-10, 1.400499e-10, 1.393781e-10, 1.404798e-10, 1.399317e-10, 
    1.398512e-10, 1.391493e-10, 1.387133e-10, 1.376155e-10, 1.367259e-10, 
    1.360229e-10, 1.361862e-10, 1.369591e-10, 1.383654e-10, 1.397034e-10, 
    1.394097e-10, 1.403959e-10, 1.377942e-10, 1.388817e-10, 1.384608e-10, 
    1.395599e-10, 1.371582e-10, 1.39202e-10, 1.366387e-10, 1.368623e-10, 
    1.375554e-10, 1.389557e-10, 1.392666e-10, 1.39599e-10, 1.393938e-10, 
    1.384012e-10, 1.382389e-10, 1.375385e-10, 1.373455e-10, 1.368136e-10, 
    1.363741e-10, 1.367756e-10, 1.37198e-10, 1.384016e-10, 1.394915e-10, 
    1.406855e-10, 1.409785e-10, 1.423829e-10, 1.412391e-10, 1.431295e-10, 
    1.415215e-10, 1.443118e-10, 1.393209e-10, 1.414743e-10, 1.37587e-10, 
    1.380027e-10, 1.387566e-10, 1.404946e-10, 1.395547e-10, 1.406543e-10, 
    1.382326e-10, 1.369858e-10, 1.366643e-10, 1.360656e-10, 1.36678e-10, 
    1.366281e-10, 1.372155e-10, 1.370266e-10, 1.384417e-10, 1.376805e-10, 
    1.398492e-10, 1.406456e-10, 1.429087e-10, 1.443065e-10, 1.457376e-10, 
    1.463721e-10, 1.465655e-10, 1.466464e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24574.8, 24595.09, 24591.11, 24607.71, 24598.47, 24609.38, 24578.88, 
    24595.9, 24585.01, 24576.62, 24640.64, 24608.46, 24675.11, 24653.79, 
    24707.78, 24671.76, 24715.18, 24706.72, 24732.41, 24724.98, 24758.58, 
    24735.85, 24776.47, 24753.1, 24756.72, 24735.11, 24614.86, 24636.59, 
    24613.59, 24616.66, 24615.28, 24598.66, 24590.39, 24573.27, 24576.36, 
    24588.94, 24618.04, 24608.07, 24633.37, 24632.79, 24661.59, 24648.5, 
    24697.94, 24683.78, 24725.29, 24714.68, 24724.79, 24721.71, 24724.83, 
    24709.31, 24715.93, 24702.39, 24650.94, 24665.88, 24621.94, 24596.31, 
    24579.62, 24567.93, 24569.58, 24572.72, 24589.01, 24604.56, 24616.56, 
    24624.68, 24632.71, 24657.38, 24670.69, 24700.83, 24695.35, 24704.65, 
    24713.63, 24728.89, 24726.36, 24733.15, 24704.4, 24723.41, 24692.24, 
    24700.66, 24634.9, 24610.75, 24600.65, 24591.88, 24570.85, 24585.33, 
    24579.6, 24593.28, 24602.07, 24597.71, 24624.9, 24614.24, 24671.48, 
    24646.45, 24712.58, 24696.47, 24716.48, 24706.21, 24723.87, 24707.96, 
    24735.68, 24741.82, 24737.62, 24753.85, 24707.09, 24724.79, 24597.59, 
    24598.3, 24601.61, 24587.14, 24586.26, 24573.18, 24584.81, 24589.8, 
    24602.58, 24610.21, 24617.53, 24633.76, 24652.14, 24678.45, 24697.5, 
    24710.48, 24702.5, 24709.54, 24701.67, 24698.01, 24739.52, 24715.99, 
    24751.49, 24749.5, 24733.31, 24749.72, 24598.8, 24594.72, 24580.7, 
    24591.65, 24571.76, 24582.85, 24589.28, 24614.47, 24620.08, 24625.32, 
    24635.7, 24649.17, 24673.25, 24694.47, 24714.15, 24712.7, 24713.21, 
    24717.66, 24706.67, 24719.47, 24721.64, 24715.99, 24749.23, 24739.62, 
    24749.45, 24743.19, 24596.04, 24602.92, 24599.2, 24606.21, 24601.27, 
    24623.44, 24630.16, 24662.16, 24648.9, 24670.09, 24651.03, 24654.38, 
    24670.79, 24652.05, 24693.3, 24665.21, 24717.83, 24689.32, 24719.65, 
    24714.06, 24723.32, 24731.69, 24742.31, 24762.22, 24757.57, 24774.47, 
    24613.26, 24622.34, 24621.54, 24631.1, 24638.21, 24653.8, 24679.34, 
    24669.65, 24687.39, 24690.95, 24664.04, 24680.58, 24628.46, 24636.7, 
    24631.79, 24613.97, 24671.88, 24641.78, 24697.82, 24681.23, 24730.5, 
    24705.67, 24755.02, 24776.93, 24798.02, 24823.09, 24627.33, 24621.12, 
    24632.24, 24647.79, 24662.44, 24682.23, 24684.25, 24687.96, 24697.62, 
    24705.82, 24689.13, 24707.89, 24638.62, 24674.54, 24618.79, 24635.28, 
    24646.87, 24641.76, 24668.55, 24674.98, 24701.18, 24687.59, 24771.47, 
    24733.47, 24842.38, 24811.07, 24618.96, 24627.31, 24656.77, 24642.64, 
    24683.55, 24693.73, 24702.09, 24712.88, 24714.06, 24720.52, 24709.95, 
    24720.1, 24682.28, 24698.99, 24653.36, 24664.34, 24659.27, 24653.74, 
    24670.91, 24689.39, 24689.79, 24695.74, 24712.73, 24683.72, 24776.5, 
    24718.16, 24636.45, 24652.79, 24655.15, 24648.77, 24692.71, 24676.69, 
    24720.36, 24708.37, 24728.1, 24718.24, 24716.8, 24704.32, 24696.63, 
    24677.43, 24661.86, 24649.69, 24652.51, 24665.92, 24690.53, 24714.16, 
    24708.94, 24726.58, 24680.57, 24699.59, 24692.2, 24711.61, 24669.4, 
    24705.26, 24660.34, 24664.23, 24676.37, 24700.9, 24706.39, 24712.3, 
    24708.65, 24691.15, 24688.31, 24676.07, 24672.68, 24663.38, 24655.76, 
    24662.72, 24670.1, 24691.16, 24710.39, 24731.81, 24737.12, 24762.9, 
    24741.87, 24776.84, 24747.03, 24799.26, 24707.36, 24746.16, 24676.92, 
    24684.2, 24697.39, 24728.37, 24711.51, 24731.25, 24688.2, 24666.39, 
    24660.79, 24650.43, 24661.03, 24660.16, 24670.4, 24667.1, 24691.86, 
    24678.57, 24716.77, 24731.09, 24772.69, 24799.15, 24826.6, 24838.84, 
    24842.59, 24844.16 ;

 GC_ICE1 =
  17684.48, 17716.97, 17710.6, 17737.19, 17722.39, 17739.87, 17691.01, 
    17718.28, 17700.82, 17687.38, 17789.9, 17738.38, 17845.04, 17810.95, 
    17897.21, 17839.69, 17909.02, 17895.52, 17936.51, 17924.66, 17978.25, 
    17942, 18006.78, 17969.51, 17975.28, 17940.82, 17748.64, 17783.43, 
    17746.6, 17751.52, 17749.31, 17722.7, 17709.44, 17682.01, 17686.96, 
    17707.12, 17753.74, 17737.76, 17778.26, 17777.34, 17823.43, 17802.48, 
    17881.5, 17858.9, 17925.15, 17908.21, 17924.35, 17919.44, 17924.41, 
    17899.65, 17910.21, 17888.61, 17806.38, 17830.29, 17759.98, 17718.93, 
    17692.2, 17673.46, 17676.1, 17681.14, 17707.24, 17732.14, 17751.37, 
    17764.36, 17777.21, 17816.68, 17837.97, 17886.12, 17877.37, 17892.22, 
    17906.54, 17930.9, 17926.86, 17937.69, 17891.82, 17922.15, 17872.4, 
    17885.85, 17780.73, 17742.06, 17725.88, 17711.83, 17678.13, 17701.33, 
    17692.16, 17714.07, 17728.15, 17721.17, 17764.71, 17747.65, 17839.24, 
    17799.19, 17904.86, 17879.16, 17911.09, 17894.71, 17922.89, 17897.5, 
    17941.73, 17951.52, 17944.83, 17970.7, 17896.11, 17924.35, 17720.98, 
    17722.12, 17727.42, 17704.24, 17702.83, 17681.87, 17700.51, 17708.5, 
    17728.97, 17741.2, 17752.91, 17778.89, 17808.3, 17850.39, 17880.81, 
    17901.51, 17888.78, 17900.02, 17887.46, 17881.62, 17947.85, 17910.31, 
    17966.95, 17963.77, 17937.95, 17964.12, 17722.91, 17716.38, 17693.91, 
    17711.47, 17679.6, 17697.37, 17707.67, 17748.01, 17757, 17765.39, 17782, 
    17803.54, 17842.08, 17875.97, 17907.38, 17905.05, 17905.87, 17912.97, 
    17895.45, 17915.87, 17919.32, 17910.31, 17963.34, 17948.02, 17963.7, 
    17953.7, 17718.5, 17729.52, 17723.56, 17734.79, 17726.87, 17762.37, 
    17773.14, 17824.34, 17803.12, 17837.02, 17806.53, 17811.89, 17838.14, 
    17808.16, 17874.1, 17829.22, 17913.25, 17867.75, 17916.15, 17907.24, 
    17922.01, 17935.37, 17952.31, 17984.06, 17976.65, 18003.6, 17746.07, 
    17760.62, 17759.33, 17774.65, 17786.02, 17810.96, 17851.81, 17836.32, 
    17864.66, 17870.35, 17827.34, 17853.8, 17770.42, 17783.59, 17775.73, 
    17747.22, 17839.88, 17791.72, 17881.32, 17854.84, 17933.46, 17893.85, 
    17972.58, 18007.51, 18041.15, 18081.06, 17768.61, 17758.66, 17776.47, 
    17801.34, 17824.78, 17856.44, 17859.66, 17865.57, 17881, 17894.09, 
    17867.45, 17897.39, 17786.67, 17844.13, 17754.92, 17781.32, 17799.87, 
    17791.7, 17834.56, 17844.84, 17886.68, 17864.99, 17998.81, 17938.2, 
    18111.72, 18061.94, 17755.2, 17768.58, 17815.71, 17793.11, 17858.54, 
    17874.79, 17888.13, 17905.36, 17907.22, 17917.54, 17900.68, 17916.87, 
    17856.5, 17883.18, 17810.25, 17827.82, 17819.71, 17810.87, 17838.33, 
    17867.87, 17868.49, 17878, 17905.11, 17858.8, 18006.83, 17913.77, 
    17783.19, 17809.35, 17813.12, 17802.91, 17873.15, 17847.57, 17917.29, 
    17898.16, 17929.63, 17913.91, 17911.61, 17891.68, 17879.41, 17848.75, 
    17823.85, 17804.38, 17808.89, 17830.35, 17869.67, 17907.4, 17899.05, 
    17927.21, 17853.78, 17884.14, 17872.34, 17903.31, 17835.91, 17893.18, 
    17821.42, 17827.65, 17847.06, 17886.23, 17895, 17904.43, 17898.6, 
    17870.67, 17866.14, 17846.58, 17841.16, 17826.29, 17814.09, 17825.23, 
    17837.03, 17870.68, 17901.37, 17935.56, 17944.03, 17985.13, 17951.6, 
    18007.37, 17959.83, 18043.11, 17896.54, 17958.44, 17847.95, 17859.57, 
    17880.63, 17930.06, 17903.17, 17934.66, 17865.96, 17831.1, 17822.13, 
    17805.56, 17822.52, 17821.13, 17837.52, 17832.23, 17871.8, 17850.58, 
    17911.55, 17934.41, 18000.75, 18042.95, 18086.64, 18106.09, 18112.05, 
    18114.55 ;

 GC_LIQ1 =
  5232.647, 5234.676, 5234.278, 5235.939, 5235.014, 5236.107, 5233.055, 
    5234.757, 5233.667, 5232.828, 5239.248, 5236.014, 5242.726, 5240.575, 
    5246.076, 5242.388, 5246.837, 5245.967, 5248.61, 5247.845, 5251.311, 
    5248.965, 5253.16, 5250.745, 5251.119, 5248.889, 5236.656, 5238.839, 
    5236.528, 5236.836, 5236.697, 5235.033, 5234.206, 5232.494, 5232.802, 
    5234.061, 5236.975, 5235.975, 5238.514, 5238.456, 5241.362, 5240.041, 
    5245.063, 5243.608, 5247.877, 5246.785, 5247.825, 5247.509, 5247.83, 
    5246.233, 5246.914, 5245.521, 5240.287, 5241.795, 5237.365, 5234.798, 
    5233.129, 5231.962, 5232.126, 5232.44, 5234.068, 5235.624, 5236.826, 
    5237.639, 5238.447, 5240.936, 5242.28, 5245.361, 5244.797, 5245.754, 
    5246.677, 5248.248, 5247.987, 5248.686, 5245.729, 5247.684, 5244.478, 
    5245.343, 5238.669, 5236.244, 5235.232, 5234.354, 5232.253, 5233.699, 
    5233.126, 5234.495, 5235.375, 5234.938, 5237.662, 5236.594, 5242.36, 
    5239.833, 5246.569, 5244.913, 5246.97, 5245.915, 5247.731, 5246.095, 
    5248.948, 5249.581, 5249.147, 5250.822, 5246.005, 5247.826, 5234.926, 
    5234.997, 5235.328, 5233.88, 5233.792, 5232.485, 5233.647, 5234.147, 
    5235.425, 5236.19, 5236.922, 5238.553, 5240.408, 5243.063, 5245.019, 
    5246.353, 5245.533, 5246.256, 5245.448, 5245.071, 5249.343, 5246.92, 
    5250.58, 5250.374, 5248.703, 5250.396, 5235.047, 5234.639, 5233.236, 
    5234.332, 5232.344, 5233.452, 5234.095, 5236.616, 5237.179, 5237.704, 
    5238.749, 5240.107, 5242.539, 5244.707, 5246.731, 5246.581, 5246.634, 
    5247.092, 5245.962, 5247.278, 5247.501, 5246.92, 5250.346, 5249.354, 
    5250.369, 5249.722, 5234.771, 5235.459, 5235.087, 5235.789, 5235.294, 
    5237.515, 5238.191, 5241.419, 5240.081, 5242.22, 5240.296, 5240.634, 
    5242.291, 5240.398, 5244.586, 5241.727, 5247.109, 5244.178, 5247.296, 
    5246.722, 5247.675, 5248.536, 5249.631, 5251.688, 5251.208, 5252.954, 
    5236.495, 5237.405, 5237.325, 5238.286, 5239.002, 5240.575, 5243.154, 
    5242.176, 5243.979, 5244.345, 5241.608, 5243.279, 5238.019, 5238.85, 
    5238.354, 5236.566, 5242.4, 5239.362, 5245.052, 5243.346, 5248.413, 
    5245.859, 5250.944, 5253.207, 5255.388, 5258.006, 5237.905, 5237.283, 
    5238.4, 5239.969, 5241.447, 5243.449, 5243.657, 5244.038, 5245.031, 
    5245.875, 5244.158, 5246.087, 5239.043, 5242.669, 5237.049, 5238.707, 
    5239.875, 5239.361, 5242.064, 5242.713, 5245.397, 5244, 5252.644, 
    5248.72, 5260.051, 5256.74, 5237.066, 5237.903, 5240.875, 5239.449, 
    5243.584, 5244.631, 5245.49, 5246.601, 5246.721, 5247.386, 5246.299, 
    5247.343, 5243.454, 5245.172, 5240.53, 5241.639, 5241.127, 5240.569, 
    5242.303, 5244.185, 5244.226, 5244.837, 5246.584, 5243.602, 5253.163, 
    5247.143, 5238.824, 5240.474, 5240.711, 5240.067, 5244.525, 5242.886, 
    5247.37, 5246.137, 5248.166, 5247.152, 5247.004, 5245.719, 5244.929, 
    5242.96, 5241.389, 5240.161, 5240.445, 5241.799, 5244.301, 5246.732, 
    5246.194, 5248.01, 5243.278, 5245.233, 5244.473, 5246.469, 5242.15, 
    5245.816, 5241.235, 5241.628, 5242.854, 5245.368, 5245.933, 5246.541, 
    5246.165, 5244.366, 5244.074, 5242.823, 5242.481, 5241.542, 5240.772, 
    5241.476, 5242.22, 5244.367, 5246.344, 5248.549, 5249.096, 5251.757, 
    5249.585, 5253.198, 5250.118, 5255.516, 5246.032, 5250.029, 5242.91, 
    5243.651, 5245.007, 5248.193, 5246.459, 5248.491, 5244.063, 5241.846, 
    5241.28, 5240.235, 5241.304, 5241.217, 5242.251, 5241.917, 5244.438, 
    5243.076, 5247, 5248.474, 5252.769, 5255.505, 5258.377, 5259.674, 
    5260.073, 5260.24 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.721779e-09, 8.760239e-09, 8.752763e-09, 8.783783e-09, 8.766576e-09, 
    8.786889e-09, 8.729577e-09, 8.761765e-09, 8.741218e-09, 8.725243e-09, 
    8.843984e-09, 8.785168e-09, 8.905094e-09, 8.867578e-09, 8.961829e-09, 
    8.899256e-09, 8.974446e-09, 8.960026e-09, 9.003435e-09, 8.990999e-09, 
    9.046522e-09, 9.009176e-09, 9.075309e-09, 9.037604e-09, 9.043501e-09, 
    9.007944e-09, 8.797006e-09, 8.836661e-09, 8.794656e-09, 8.800311e-09, 
    8.797774e-09, 8.766931e-09, 8.751387e-09, 8.718841e-09, 8.72475e-09, 
    8.748655e-09, 8.802854e-09, 8.784457e-09, 8.830827e-09, 8.82978e-09, 
    8.881405e-09, 8.858128e-09, 8.944906e-09, 8.920241e-09, 8.991519e-09, 
    8.973593e-09, 8.990676e-09, 8.985496e-09, 8.990743e-09, 8.964453e-09, 
    8.975717e-09, 8.952584e-09, 8.862487e-09, 8.888963e-09, 8.809998e-09, 
    8.762518e-09, 8.730988e-09, 8.708613e-09, 8.711777e-09, 8.717806e-09, 
    8.748795e-09, 8.777933e-09, 8.800138e-09, 8.814992e-09, 8.829629e-09, 
    8.873928e-09, 8.897381e-09, 8.949892e-09, 8.940417e-09, 8.95647e-09, 
    8.971809e-09, 8.997559e-09, 8.993322e-09, 9.004666e-09, 8.956048e-09, 
    8.988359e-09, 8.93502e-09, 8.949608e-09, 8.833601e-09, 8.78942e-09, 
    8.770636e-09, 8.754199e-09, 8.714209e-09, 8.741825e-09, 8.730938e-09, 
    8.756841e-09, 8.773299e-09, 8.765158e-09, 8.815399e-09, 8.795866e-09, 
    8.898771e-09, 8.854444e-09, 8.970019e-09, 8.942362e-09, 8.97665e-09, 
    8.959153e-09, 8.989131e-09, 8.962152e-09, 9.008889e-09, 9.019065e-09, 
    9.012111e-09, 9.038828e-09, 8.960656e-09, 8.990675e-09, 8.76493e-09, 
    8.766258e-09, 8.772443e-09, 8.745254e-09, 8.743592e-09, 8.718678e-09, 
    8.740846e-09, 8.750287e-09, 8.774253e-09, 8.788429e-09, 8.801904e-09, 
    8.831535e-09, 8.864626e-09, 8.910904e-09, 8.944155e-09, 8.966444e-09, 
    8.952777e-09, 8.964842e-09, 8.951354e-09, 8.945032e-09, 9.015252e-09, 
    8.975822e-09, 9.034986e-09, 9.031712e-09, 9.004935e-09, 9.032081e-09, 
    8.76719e-09, 8.75955e-09, 8.733026e-09, 8.753783e-09, 8.715966e-09, 
    8.737134e-09, 8.749304e-09, 8.796273e-09, 8.806595e-09, 8.816163e-09, 
    8.835063e-09, 8.859319e-09, 8.901871e-09, 8.938898e-09, 8.972702e-09, 
    8.970225e-09, 8.971097e-09, 8.978648e-09, 8.959943e-09, 8.981718e-09, 
    8.985372e-09, 8.975817e-09, 9.031274e-09, 9.01543e-09, 9.031643e-09, 
    9.021327e-09, 8.762034e-09, 8.774888e-09, 8.767943e-09, 8.781004e-09, 
    8.771802e-09, 8.81272e-09, 8.82499e-09, 8.882402e-09, 8.858842e-09, 
    8.896341e-09, 8.862651e-09, 8.868621e-09, 8.897562e-09, 8.864472e-09, 
    8.936855e-09, 8.887779e-09, 8.978941e-09, 8.929927e-09, 8.982012e-09, 
    8.972555e-09, 8.988215e-09, 9.002238e-09, 9.019883e-09, 9.052438e-09, 
    9.0449e-09, 9.072127e-09, 8.794053e-09, 8.810726e-09, 8.80926e-09, 
    8.826709e-09, 8.839614e-09, 8.867588e-09, 8.912455e-09, 8.895584e-09, 
    8.926559e-09, 8.932777e-09, 8.885719e-09, 8.91461e-09, 8.821886e-09, 
    8.836865e-09, 8.827947e-09, 8.795368e-09, 8.89947e-09, 8.846041e-09, 
    8.944704e-09, 8.915759e-09, 9.000238e-09, 8.958223e-09, 9.040749e-09, 
    9.076029e-09, 9.109239e-09, 9.148044e-09, 8.819828e-09, 8.808498e-09, 
    8.828785e-09, 8.856851e-09, 8.882898e-09, 8.917524e-09, 8.921067e-09, 
    8.927554e-09, 8.944358e-09, 8.958486e-09, 8.929604e-09, 8.962028e-09, 
    8.840336e-09, 8.904108e-09, 8.804214e-09, 8.834291e-09, 8.855197e-09, 
    8.846028e-09, 8.893656e-09, 8.90488e-09, 8.950497e-09, 8.926917e-09, 
    9.06732e-09, 9.005198e-09, 9.177597e-09, 9.129415e-09, 8.804539e-09, 
    8.819789e-09, 8.872864e-09, 8.847611e-09, 8.919836e-09, 8.937614e-09, 
    8.952069e-09, 8.970544e-09, 8.97254e-09, 8.983486e-09, 8.965548e-09, 
    8.982778e-09, 8.917597e-09, 8.946725e-09, 8.866799e-09, 8.886251e-09, 
    8.877302e-09, 8.867486e-09, 8.897782e-09, 8.930058e-09, 8.93075e-09, 
    8.941099e-09, 8.970259e-09, 8.920129e-09, 9.075334e-09, 8.979476e-09, 
    8.836419e-09, 8.86579e-09, 8.869988e-09, 8.85861e-09, 8.935833e-09, 
    8.90785e-09, 8.98322e-09, 8.96285e-09, 8.996227e-09, 8.979641e-09, 
    8.9772e-09, 8.955899e-09, 8.942638e-09, 8.909133e-09, 8.881874e-09, 
    8.86026e-09, 8.865286e-09, 8.889029e-09, 8.932033e-09, 8.972719e-09, 
    8.963807e-09, 8.99369e-09, 8.914599e-09, 8.947762e-09, 8.934943e-09, 
    8.968366e-09, 8.895134e-09, 8.957489e-09, 8.879196e-09, 8.886061e-09, 
    8.907295e-09, 8.950009e-09, 8.959463e-09, 8.969553e-09, 8.963327e-09, 
    8.933125e-09, 8.928178e-09, 8.906779e-09, 8.90087e-09, 8.884567e-09, 
    8.871067e-09, 8.883401e-09, 8.896352e-09, 8.933139e-09, 8.966291e-09, 
    9.002437e-09, 9.011284e-09, 9.053515e-09, 9.019135e-09, 9.075867e-09, 
    9.027629e-09, 9.111137e-09, 8.961106e-09, 9.026214e-09, 8.908263e-09, 
    8.920969e-09, 8.943951e-09, 8.996667e-09, 8.968209e-09, 9.001493e-09, 
    8.927985e-09, 8.889847e-09, 8.879982e-09, 8.861574e-09, 8.880403e-09, 
    8.878872e-09, 8.896889e-09, 8.8911e-09, 8.93436e-09, 8.911123e-09, 
    8.977139e-09, 9.00123e-09, 9.069273e-09, 9.110987e-09, 9.153455e-09, 
    9.172203e-09, 9.17791e-09, 9.180296e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.152127, 6.181118, 6.175474, 6.19891, 6.185902, 6.201259, 6.157997, 
    6.182271, 6.166767, 6.154732, 6.244562, 6.199957, 6.291116, 6.262504, 
    6.33454, 6.286658, 6.344223, 6.333154, 6.366505, 6.356939, 6.399723, 
    6.370924, 6.421972, 6.392837, 6.397389, 6.369975, 6.208915, 6.238997, 
    6.207136, 6.211419, 6.209496, 6.186171, 6.174439, 6.149914, 6.154361, 
    6.172376, 6.213346, 6.199417, 6.234558, 6.233763, 6.273037, 6.255309, 
    6.321565, 6.302687, 6.357338, 6.343565, 6.356691, 6.352709, 6.356743, 
    6.336551, 6.345197, 6.327448, 6.258627, 6.278802, 6.218759, 6.182842, 
    6.15906, 6.142222, 6.144601, 6.149137, 6.172482, 6.194484, 6.211287, 
    6.222544, 6.233648, 6.267345, 6.285226, 6.325387, 6.318126, 6.330429, 
    6.342196, 6.361985, 6.358725, 6.367453, 6.330103, 6.354911, 6.313993, 
    6.325167, 6.236673, 6.203172, 6.188972, 6.176558, 6.14643, 6.167226, 
    6.159022, 6.17855, 6.190981, 6.184831, 6.222852, 6.208052, 6.286287, 
    6.252509, 6.340823, 6.319615, 6.345912, 6.332485, 6.355504, 6.334785, 
    6.370704, 6.378543, 6.373185, 6.39378, 6.333637, 6.356691, 6.184659, 
    6.185661, 6.190334, 6.169812, 6.168558, 6.149792, 6.166487, 6.173606, 
    6.191701, 6.202422, 6.212625, 6.235096, 6.260257, 6.295552, 6.320989, 
    6.338078, 6.327595, 6.336849, 6.326505, 6.321661, 6.375605, 6.345278, 
    6.390815, 6.38829, 6.367661, 6.388575, 6.186365, 6.180596, 6.160594, 
    6.176244, 6.147751, 6.16369, 6.172867, 6.208362, 6.216177, 6.223432, 
    6.237775, 6.256216, 6.288652, 6.316964, 6.342881, 6.34098, 6.341649, 
    6.347448, 6.33309, 6.349807, 6.352615, 6.345274, 6.387952, 6.37574, 
    6.388237, 6.380283, 6.182471, 6.192183, 6.186934, 6.196806, 6.18985, 
    6.220824, 6.230131, 6.2738, 6.255853, 6.284431, 6.258751, 6.263297, 
    6.285367, 6.260137, 6.315401, 6.2779, 6.347673, 6.310101, 6.350032, 
    6.342769, 6.354798, 6.365584, 6.37917, 6.404289, 6.398467, 6.419509, 
    6.206679, 6.219311, 6.218197, 6.231433, 6.241233, 6.26251, 6.296736, 
    6.283851, 6.307518, 6.312277, 6.276325, 6.298384, 6.227774, 6.239147, 
    6.232373, 6.207675, 6.286819, 6.246119, 6.32141, 6.29926, 6.364046, 
    6.331773, 6.395263, 6.422532, 6.448259, 6.478412, 6.226212, 6.21762, 
    6.233008, 6.254341, 6.274175, 6.30061, 6.303318, 6.30828, 6.321144, 
    6.331974, 6.30985, 6.33469, 6.241788, 6.29036, 6.214375, 6.237192, 
    6.253081, 6.246107, 6.282379, 6.290948, 6.32585, 6.307792, 6.415795, 
    6.367866, 6.501428, 6.463926, 6.214621, 6.226182, 6.26653, 6.24731, 
    6.302377, 6.31598, 6.327053, 6.341226, 6.342757, 6.351165, 6.33739, 
    6.350621, 6.300666, 6.322958, 6.261909, 6.276732, 6.269909, 6.262432, 
    6.285529, 6.310198, 6.310725, 6.318649, 6.341017, 6.3026, 6.422, 
    6.348093, 6.238804, 6.261144, 6.264338, 6.255675, 6.314616, 6.293218, 
    6.35096, 6.33532, 6.360959, 6.34821, 6.346336, 6.329989, 6.319827, 
    6.294198, 6.273396, 6.256931, 6.260757, 6.278851, 6.311709, 6.342896, 
    6.336056, 6.359008, 6.298373, 6.323753, 6.313936, 6.339554, 6.283509, 
    6.331217, 6.271353, 6.276586, 6.292793, 6.325478, 6.332722, 6.340465, 
    6.335686, 6.312545, 6.308758, 6.292399, 6.287888, 6.275446, 6.26516, 
    6.274558, 6.284439, 6.312554, 6.337962, 6.365738, 6.372547, 6.405127, 
    6.378599, 6.422414, 6.385153, 6.44974, 6.333988, 6.384058, 6.293531, 
    6.303243, 6.320835, 6.361302, 6.339433, 6.365013, 6.308609, 6.279477, 
    6.271952, 6.257931, 6.272273, 6.271106, 6.284847, 6.280429, 6.313488, 
    6.295716, 6.346289, 6.36481, 6.417302, 6.449619, 6.482619, 6.497222, 
    6.501671, 6.503531,
  3.942679, 3.961972, 3.958216, 3.9738, 3.965154, 3.975316, 3.946585, 
    3.96274, 3.952421, 3.944412, 4.003285, 3.974475, 4.03333, 4.01486, 
    4.061353, 4.030455, 4.0676, 4.060456, 4.081971, 4.0758, 4.103403, 
    4.084821, 4.11775, 4.098959, 4.101897, 4.08421, 3.980259, 3.999692, 
    3.97911, 3.981877, 3.980635, 3.965334, 3.95753, 3.941205, 3.944165, 
    3.956155, 3.983122, 3.974125, 3.996816, 3.996303, 4.021659, 4.010214, 
    4.052978, 4.040794, 4.076057, 4.067173, 4.075641, 4.073071, 4.075674, 
    4.062647, 4.068226, 4.056773, 4.012357, 4.025381, 3.986617, 3.963123, 
    3.947293, 3.936086, 3.937669, 3.940689, 3.956226, 3.970864, 3.98179, 
    3.989059, 3.996229, 4.017991, 4.029529, 4.055446, 4.050758, 4.058699, 
    4.066289, 4.079056, 4.076952, 4.082584, 4.058486, 4.074493, 4.04809, 
    4.055302, 3.998193, 3.97655, 3.967201, 3.958938, 3.938887, 3.952728, 
    3.947268, 3.960262, 3.968533, 3.964441, 3.989258, 3.979701, 4.030214, 
    4.008408, 4.065403, 4.051719, 4.068686, 4.060022, 4.074876, 4.061506, 
    4.084681, 4.089738, 4.086282, 4.099566, 4.060767, 4.075642, 3.964326, 
    3.964994, 3.968102, 3.954449, 3.953614, 3.941124, 3.952235, 3.956973, 
    3.969012, 3.976066, 3.982655, 3.997165, 4.013411, 4.036192, 4.052606, 
    4.063631, 4.056868, 4.062839, 4.056164, 4.053038, 4.087844, 4.068279, 
    4.097653, 4.096024, 4.082719, 4.096208, 3.965462, 3.961623, 3.948314, 
    3.958727, 3.939766, 3.950374, 3.956482, 3.979904, 3.984948, 3.989634, 
    3.998894, 4.0108, 4.031739, 4.050009, 4.06673, 4.065504, 4.065935, 
    4.069677, 4.060414, 4.071199, 4.073012, 4.068275, 4.095806, 4.087929, 
    4.095989, 4.090859, 3.96287, 3.969333, 3.96584, 3.97241, 3.967782, 
    3.987952, 3.993962, 4.022154, 4.010566, 4.029015, 4.012437, 4.015372, 
    4.029623, 4.01333, 4.049003, 4.024802, 4.069823, 4.045585, 4.071345, 
    4.066658, 4.074419, 4.081378, 4.090142, 4.106346, 4.102589, 4.11616, 
    3.978815, 3.986974, 3.986252, 3.994799, 4.001128, 4.014863, 4.036955, 
    4.028638, 4.043912, 4.046984, 4.02378, 4.038019, 3.992438, 3.999783, 
    3.995407, 3.979459, 4.030557, 4.004285, 4.052878, 4.038584, 4.080386, 
    4.059566, 4.100523, 4.118114, 4.134699, 4.154144, 3.991428, 3.98588, 
    3.995816, 4.009592, 4.022393, 4.039455, 4.041202, 4.044405, 4.052705, 
    4.059693, 4.04542, 4.061446, 4.001493, 4.032841, 3.983785, 3.998522, 
    4.008778, 4.004274, 4.027687, 4.033218, 4.055744, 4.044088, 4.11377, 
    4.082853, 4.168978, 4.144804, 3.983943, 3.991408, 4.017459, 4.005051, 
    4.040594, 4.049374, 4.056517, 4.065664, 4.06665, 4.072076, 4.063188, 
    4.071724, 4.039491, 4.053876, 4.014473, 4.024044, 4.019639, 4.014812, 
    4.02972, 4.045645, 4.045982, 4.051097, 4.06554, 4.040739, 4.117778, 
    4.070104, 3.999558, 4.013985, 4.016043, 4.01045, 4.048493, 4.034684, 
    4.071943, 4.061852, 4.078393, 4.070169, 4.06896, 4.058413, 4.051856, 
    4.035317, 4.02189, 4.011261, 4.01373, 4.025412, 4.046619, 4.066742, 
    4.062329, 4.077135, 4.038011, 4.05439, 4.048056, 4.064584, 4.028418, 
    4.059216, 4.02057, 4.023949, 4.03441, 4.055506, 4.060176, 4.065173, 
    4.062088, 4.047158, 4.044713, 4.034154, 4.031244, 4.023212, 4.016572, 
    4.02264, 4.029019, 4.047163, 4.063558, 4.081478, 4.085869, 4.106891, 
    4.089779, 4.118046, 4.094015, 4.135663, 4.060998, 4.093301, 4.034885, 
    4.041153, 4.052509, 4.078619, 4.064507, 4.081013, 4.044617, 4.025817, 
    4.020957, 4.011907, 4.021164, 4.020411, 4.029281, 4.026429, 4.047766, 
    4.036296, 4.068931, 4.080881, 4.114738, 4.135579, 4.156851, 4.166265, 
    4.169133, 4.170332,
  3.294122, 3.311954, 3.308482, 3.322676, 3.314897, 3.324076, 3.297731, 
    3.312665, 3.303126, 3.295723, 3.349906, 3.3233, 3.377674, 3.360601, 
    3.403591, 3.375016, 3.409371, 3.402761, 3.422672, 3.41696, 3.442516, 
    3.42531, 3.455805, 3.4384, 3.44112, 3.424744, 3.32864, 3.346587, 3.32758, 
    3.330134, 3.328987, 3.315063, 3.307848, 3.29276, 3.295495, 3.306578, 
    3.331284, 3.322977, 3.343931, 3.343457, 3.366886, 3.356309, 3.395843, 
    3.384576, 3.417198, 3.408976, 3.416812, 3.414434, 3.416843, 3.404789, 
    3.40995, 3.399354, 3.358289, 3.370326, 3.334511, 3.313019, 3.298386, 
    3.288029, 3.289492, 3.292283, 3.306643, 3.320035, 3.330054, 3.336766, 
    3.343389, 3.363494, 3.37416, 3.398126, 3.39379, 3.401135, 3.408158, 
    3.419974, 3.418027, 3.423239, 3.400939, 3.415751, 3.391322, 3.397993, 
    3.345202, 3.325216, 3.316754, 3.30915, 3.290618, 3.303409, 3.298363, 
    3.310374, 3.317947, 3.314237, 3.33695, 3.328125, 3.374793, 3.35464, 
    3.407339, 3.394679, 3.410377, 3.40236, 3.416105, 3.403733, 3.42518, 
    3.429862, 3.426662, 3.438962, 3.403049, 3.416813, 3.314132, 3.314749, 
    3.317561, 3.305, 3.304228, 3.292685, 3.302954, 3.307334, 3.318376, 
    3.324769, 3.330852, 3.344253, 3.359262, 3.38032, 3.395499, 3.405699, 
    3.399441, 3.404966, 3.398791, 3.395899, 3.428108, 3.409999, 3.437191, 
    3.435682, 3.423364, 3.435852, 3.315182, 3.311632, 3.29933, 3.308955, 
    3.29143, 3.301234, 3.30688, 3.328312, 3.33297, 3.337297, 3.34585, 
    3.35685, 3.376203, 3.393098, 3.408566, 3.407431, 3.407831, 3.411294, 
    3.402722, 3.412702, 3.41438, 3.409996, 3.43548, 3.428187, 3.43565, 
    3.4309, 3.312786, 3.318663, 3.315531, 3.321421, 3.317273, 3.335744, 
    3.341294, 3.367343, 3.356634, 3.373685, 3.358362, 3.361075, 3.374247, 
    3.359189, 3.392167, 3.36979, 3.411428, 3.389006, 3.412837, 3.408499, 
    3.415681, 3.422123, 3.430236, 3.445241, 3.441762, 3.454332, 3.327307, 
    3.33484, 3.334174, 3.342068, 3.347914, 3.360604, 3.381026, 3.373336, 
    3.387459, 3.390299, 3.368846, 3.38201, 3.339887, 3.346672, 3.342629, 
    3.327902, 3.37511, 3.35083, 3.395751, 3.382531, 3.421205, 3.401938, 
    3.439848, 3.456142, 3.471511, 3.489539, 3.338954, 3.33383, 3.343007, 
    3.355734, 3.367564, 3.383337, 3.384953, 3.387914, 3.395591, 3.402056, 
    3.388853, 3.403677, 3.348251, 3.377222, 3.331896, 3.345506, 3.354982, 
    3.350821, 3.372458, 3.377571, 3.398402, 3.387622, 3.452118, 3.423488, 
    3.503297, 3.480878, 3.332042, 3.338936, 3.363004, 3.351538, 3.384391, 
    3.39251, 3.399118, 3.40758, 3.408493, 3.413514, 3.405289, 3.413188, 
    3.383371, 3.396674, 3.360245, 3.36909, 3.365018, 3.360557, 3.374337, 
    3.389061, 3.389373, 3.394104, 3.407465, 3.384524, 3.455831, 3.411688, 
    3.346464, 3.359793, 3.361695, 3.356527, 3.391695, 3.378926, 3.413391, 
    3.404053, 3.41936, 3.411749, 3.41063, 3.400871, 3.394805, 3.379511, 
    3.367099, 3.357276, 3.359558, 3.370354, 3.389962, 3.408577, 3.404494, 
    3.418195, 3.382002, 3.39715, 3.391291, 3.406581, 3.373133, 3.401613, 
    3.365879, 3.369002, 3.378673, 3.398181, 3.402502, 3.407126, 3.404272, 
    3.39046, 3.3882, 3.378437, 3.375746, 3.368321, 3.362184, 3.367792, 
    3.373688, 3.390465, 3.405632, 3.422215, 3.42628, 3.445746, 3.429899, 
    3.456079, 3.433821, 3.472404, 3.403263, 3.433161, 3.379112, 3.384907, 
    3.39541, 3.419569, 3.406509, 3.421784, 3.388111, 3.370729, 3.366237, 
    3.357873, 3.366428, 3.365732, 3.37393, 3.371294, 3.391023, 3.380416, 
    3.410603, 3.421663, 3.453015, 3.472327, 3.492049, 3.500781, 3.503441, 
    3.504553,
  3.016762, 3.03369, 3.030393, 3.044087, 3.036484, 3.04546, 3.020187, 
    3.034364, 3.025308, 3.018281, 3.070795, 3.044699, 3.098064, 3.081296, 
    3.123541, 3.095452, 3.129226, 3.122725, 3.142315, 3.136694, 3.161406, 
    3.144912, 3.174079, 3.157482, 3.160076, 3.144355, 3.049935, 3.067538, 
    3.048895, 3.0514, 3.050275, 3.036642, 3.02979, 3.015469, 3.018065, 
    3.028584, 3.052527, 3.044382, 3.064934, 3.064469, 3.087467, 3.077082, 
    3.115922, 3.104846, 3.136928, 3.128838, 3.136548, 3.134209, 3.136579, 
    3.124719, 3.129797, 3.119375, 3.079025, 3.090845, 3.055692, 3.0347, 
    3.020808, 3.010981, 3.012369, 3.015017, 3.028646, 3.041499, 3.051321, 
    3.057905, 3.064402, 3.084135, 3.094611, 3.118167, 3.113904, 3.121126, 
    3.128034, 3.139659, 3.137743, 3.142874, 3.120934, 3.135503, 3.111478, 
    3.118036, 3.066179, 3.046577, 3.038282, 3.031027, 3.013437, 3.025577, 
    3.020787, 3.032189, 3.039452, 3.035858, 3.058085, 3.04943, 3.095233, 
    3.075443, 3.127228, 3.114778, 3.130217, 3.122331, 3.135852, 3.123682, 
    3.144784, 3.149346, 3.146243, 3.158018, 3.123008, 3.136549, 3.035758, 
    3.036344, 3.039074, 3.027086, 3.026354, 3.015399, 3.025144, 3.029302, 
    3.039872, 3.046139, 3.052104, 3.065249, 3.079981, 3.100664, 3.115584, 
    3.125615, 3.119461, 3.124894, 3.118821, 3.115978, 3.147666, 3.129845, 
    3.15633, 3.154892, 3.142996, 3.155055, 3.036755, 3.033384, 3.021704, 
    3.030842, 3.014207, 3.023511, 3.028871, 3.049613, 3.054182, 3.058425, 
    3.066817, 3.077613, 3.096618, 3.113223, 3.128436, 3.127319, 3.127712, 
    3.131118, 3.122687, 3.132504, 3.134155, 3.129842, 3.1547, 3.147744, 
    3.154862, 3.150335, 3.034479, 3.040154, 3.037087, 3.042857, 3.038792, 
    3.056901, 3.062346, 3.087915, 3.0774, 3.094145, 3.079098, 3.081761, 
    3.094696, 3.079909, 3.112308, 3.090319, 3.131251, 3.109199, 3.132637, 
    3.12837, 3.135436, 3.141775, 3.149702, 3.164004, 3.160688, 3.172674, 
    3.048627, 3.056015, 3.055363, 3.063106, 3.068842, 3.081299, 3.101357, 
    3.093803, 3.10768, 3.110472, 3.089392, 3.102324, 3.060966, 3.067622, 
    3.063656, 3.049211, 3.095545, 3.071703, 3.115832, 3.102837, 3.140871, 
    3.121916, 3.158863, 3.1744, 3.189066, 3.20628, 3.060051, 3.055025, 
    3.064027, 3.076516, 3.088133, 3.103629, 3.105217, 3.108128, 3.115675, 
    3.122031, 3.10905, 3.123626, 3.069171, 3.09762, 3.053128, 3.066478, 
    3.075778, 3.071695, 3.09294, 3.097963, 3.118438, 3.107841, 3.170562, 
    3.143118, 3.219428, 3.198009, 3.053271, 3.060033, 3.083655, 3.072399, 
    3.104665, 3.112645, 3.119142, 3.127465, 3.128363, 3.133302, 3.125211, 
    3.132982, 3.103662, 3.11674, 3.080946, 3.089631, 3.085633, 3.081253, 
    3.094786, 3.109255, 3.109561, 3.114212, 3.127349, 3.104796, 3.174103, 
    3.131504, 3.067419, 3.080501, 3.08237, 3.077296, 3.111845, 3.099294, 
    3.133182, 3.123996, 3.139056, 3.131566, 3.130465, 3.120867, 3.114902, 
    3.099869, 3.087676, 3.078031, 3.080271, 3.090873, 3.110141, 3.128446, 
    3.12443, 3.137909, 3.102317, 3.117207, 3.111447, 3.126482, 3.093603, 
    3.121594, 3.086478, 3.089545, 3.099045, 3.118221, 3.122471, 3.127018, 
    3.124211, 3.11063, 3.108408, 3.098814, 3.09617, 3.088877, 3.08285, 
    3.088357, 3.094148, 3.110635, 3.125548, 3.141866, 3.145867, 3.164485, 
    3.149381, 3.174339, 3.153117, 3.189918, 3.123218, 3.152488, 3.099477, 
    3.105172, 3.115496, 3.139261, 3.126411, 3.141441, 3.108321, 3.091241, 
    3.08683, 3.078617, 3.087018, 3.086334, 3.094387, 3.091797, 3.111183, 
    3.100759, 3.130439, 3.141321, 3.171418, 3.189845, 3.208679, 3.217023, 
    3.219565, 3.220629,
  2.987434, 3.004069, 3.000827, 3.014296, 3.006817, 3.015646, 2.990798, 
    3.004732, 2.995829, 2.988926, 3.0406, 3.014898, 3.06751, 3.050957, 
    3.092699, 3.064929, 3.098327, 3.091892, 3.111237, 3.105723, 3.12999, 
    3.113728, 3.142576, 3.126098, 3.12867, 3.113193, 3.020051, 3.037389, 
    3.019028, 3.021493, 3.020386, 3.006972, 3.000234, 2.986164, 2.988714, 
    2.999049, 3.022603, 3.014586, 3.034824, 3.034365, 3.057046, 3.0468, 
    3.085162, 3.074212, 3.105955, 3.097943, 3.105578, 3.103261, 3.105609, 
    3.093866, 3.098892, 3.088578, 3.048717, 3.060381, 3.025719, 3.005061, 
    2.991408, 2.981757, 2.98312, 2.98572, 2.99911, 3.011749, 3.021416, 
    3.027899, 3.0343, 3.053758, 3.0641, 3.087382, 3.083166, 3.09031, 
    3.097147, 3.10866, 3.106762, 3.111772, 3.09012, 3.104543, 3.080767, 
    3.087253, 3.036049, 3.016747, 3.008584, 3.00145, 2.984168, 2.996093, 
    2.991387, 3.002593, 3.009736, 3.006201, 3.028077, 3.019554, 3.064714, 
    3.045184, 3.096349, 3.084031, 3.099308, 3.091503, 3.104888, 3.092839, 
    3.113604, 3.118027, 3.115004, 3.12663, 3.092172, 3.105579, 3.006102, 
    3.006678, 3.009364, 2.997577, 2.996857, 2.986095, 2.995669, 2.999755, 
    3.010149, 3.016315, 3.022187, 3.035135, 3.049659, 3.070079, 3.084828, 
    3.094753, 3.088663, 3.094039, 3.08803, 3.085217, 3.116369, 3.098939, 
    3.124955, 3.123528, 3.111889, 3.123689, 3.007083, 3.003768, 2.992288, 
    3.001269, 2.984925, 2.994064, 2.999331, 3.019734, 3.024232, 3.028411, 
    3.03668, 3.047324, 3.066082, 3.082492, 3.097545, 3.096439, 3.096828, 
    3.100201, 3.091855, 3.101573, 3.103207, 3.098936, 3.123338, 3.116445, 
    3.123498, 3.119008, 3.004845, 3.010426, 3.007409, 3.013085, 3.009086, 
    3.02691, 3.032273, 3.057489, 3.047114, 3.063639, 3.048789, 3.051415, 
    3.064183, 3.049589, 3.081587, 3.059861, 3.100332, 3.078513, 3.101704, 
    3.097479, 3.104476, 3.110718, 3.118381, 3.13257, 3.129278, 3.141181, 
    3.018764, 3.026038, 3.025395, 3.033022, 3.038675, 3.05096, 3.070764, 
    3.063302, 3.077013, 3.079772, 3.058947, 3.071719, 3.030914, 3.037473, 
    3.033565, 3.019338, 3.065022, 3.041496, 3.085072, 3.072226, 3.109851, 
    3.091091, 3.127468, 3.142894, 3.157475, 3.174608, 3.030013, 3.025063, 
    3.03393, 3.046242, 3.057704, 3.073009, 3.074578, 3.077455, 3.084917, 
    3.091206, 3.078366, 3.092784, 3.038999, 3.067071, 3.023195, 3.036345, 
    3.045514, 3.041488, 3.06245, 3.067411, 3.087651, 3.077171, 3.139081, 
    3.112005, 3.18771, 3.166372, 3.023335, 3.029995, 3.053284, 3.042182, 
    3.074032, 3.081921, 3.088347, 3.096583, 3.097473, 3.102363, 3.094353, 
    3.102046, 3.073041, 3.08597, 3.050612, 3.059183, 3.055237, 3.050915, 
    3.064273, 3.078568, 3.078872, 3.08347, 3.096467, 3.074162, 3.142597, 
    3.100581, 3.037273, 3.050173, 3.052017, 3.047011, 3.081129, 3.068726, 
    3.102244, 3.09315, 3.108063, 3.100644, 3.099554, 3.090053, 3.084153, 
    3.069294, 3.057253, 3.047736, 3.049947, 3.060409, 3.079444, 3.097554, 
    3.093579, 3.106927, 3.071712, 3.086433, 3.080736, 3.095611, 3.063104, 
    3.090772, 3.056071, 3.059098, 3.06848, 3.087435, 3.09164, 3.096141, 
    3.093363, 3.079929, 3.077732, 3.068251, 3.065639, 3.058439, 3.052491, 
    3.057925, 3.063643, 3.079933, 3.094686, 3.110805, 3.114644, 3.133046, 
    3.118061, 3.142831, 3.121764, 3.158319, 3.092379, 3.121142, 3.068907, 
    3.074534, 3.08474, 3.108265, 3.095541, 3.110397, 3.077646, 3.060772, 
    3.056418, 3.048315, 3.056603, 3.055928, 3.063879, 3.061321, 3.080476, 
    3.070173, 3.099527, 3.110283, 3.139932, 3.158248, 3.176998, 3.185313, 
    3.187848, 3.188908,
  2.977508, 2.99592, 2.992333, 3.00725, 2.998963, 3.008748, 2.981243, 
    2.996654, 2.986804, 2.979175, 3.036464, 3.007918, 3.066465, 3.047998, 
    3.094651, 3.063583, 3.100963, 3.093748, 3.115525, 3.109266, 3.137337, 
    3.118419, 3.152011, 3.132804, 3.1358, 3.117797, 3.013634, 3.032892, 
    3.012498, 3.015234, 3.014005, 2.999135, 2.991677, 2.976059, 2.97894, 
    2.990366, 3.016465, 3.007573, 3.030041, 3.029531, 3.054786, 3.043367, 
    3.086207, 3.073955, 3.109527, 3.100533, 3.109104, 3.106502, 3.109138, 
    3.09596, 3.101598, 3.090033, 3.045502, 3.058506, 3.019925, 2.997019, 
    2.981917, 2.971032, 2.972586, 2.975552, 2.990433, 3.004428, 3.015148, 
    3.022346, 3.029458, 3.051119, 3.062657, 3.088693, 3.083972, 3.091974, 
    3.09964, 3.112566, 3.110434, 3.116146, 3.091761, 3.107941, 3.081287, 
    3.088549, 3.031402, 3.009968, 3.00092, 2.993022, 2.973782, 2.987096, 
    2.981894, 2.994287, 3.002197, 2.998281, 3.022543, 3.013082, 3.063342, 
    3.041567, 3.098744, 3.08494, 3.102064, 3.093311, 3.108329, 3.094809, 
    3.118275, 3.123415, 3.119901, 3.133424, 3.094062, 3.109105, 2.998172, 
    2.99881, 3.001785, 2.988737, 2.987941, 2.97598, 2.986627, 2.991147, 
    3.002655, 3.00949, 3.016003, 3.030387, 3.046552, 3.069335, 3.085833, 
    3.096954, 3.090128, 3.096154, 3.089419, 3.086269, 3.121488, 3.101651, 
    3.131474, 3.129814, 3.116282, 3.130002, 2.999258, 2.995588, 2.98289, 
    2.992822, 2.974645, 2.984853, 2.990678, 3.013281, 3.018274, 3.022915, 
    3.032105, 3.043951, 3.064871, 3.083218, 3.100086, 3.098846, 3.099283, 
    3.103066, 3.093706, 3.104606, 3.106441, 3.101648, 3.129592, 3.121576, 
    3.129779, 3.124556, 2.99678, 3.002962, 2.99962, 3.005909, 3.001477, 
    3.021247, 3.027205, 3.05528, 3.043717, 3.062143, 3.045582, 3.048509, 
    3.062749, 3.046474, 3.082204, 3.057926, 3.103213, 3.078765, 3.104754, 
    3.100013, 3.107867, 3.114922, 3.123827, 3.140343, 3.136508, 3.150383, 
    3.012206, 3.020278, 3.019565, 3.028038, 3.034324, 3.048002, 3.070101, 
    3.061767, 3.077087, 3.080174, 3.056907, 3.071168, 3.025695, 3.032986, 
    3.028641, 3.012843, 3.063686, 3.037462, 3.086107, 3.071735, 3.113915, 
    3.092849, 3.1344, 3.152382, 3.16942, 3.188975, 3.024694, 3.019196, 
    3.029047, 3.042746, 3.05552, 3.072609, 3.074364, 3.077581, 3.085933, 
    3.092978, 3.078601, 3.094747, 3.034683, 3.065975, 3.017122, 3.031732, 
    3.041935, 3.037453, 3.060816, 3.066355, 3.088994, 3.077264, 3.147933, 
    3.116417, 3.20387, 3.179629, 3.017279, 3.024674, 3.050592, 3.038226, 
    3.073754, 3.082579, 3.089775, 3.099008, 3.100005, 3.105494, 3.096507, 
    3.105138, 3.072646, 3.087113, 3.047614, 3.05717, 3.052769, 3.047951, 
    3.06285, 3.078827, 3.079167, 3.084313, 3.098876, 3.073899, 3.152035, 
    3.103492, 3.032765, 3.047124, 3.049179, 3.043602, 3.081693, 3.067823, 
    3.10536, 3.095158, 3.111895, 3.103564, 3.102341, 3.091687, 3.085077, 
    3.068458, 3.055017, 3.04441, 3.046872, 3.058538, 3.079807, 3.100097, 
    3.095638, 3.110619, 3.07116, 3.08763, 3.081252, 3.097917, 3.061546, 
    3.09249, 3.053699, 3.057076, 3.067549, 3.088753, 3.093466, 3.098511, 
    3.095396, 3.080349, 3.077891, 3.067293, 3.064376, 3.05634, 3.049707, 
    3.055767, 3.062147, 3.080354, 3.09688, 3.115023, 3.119483, 3.140897, 
    3.123454, 3.152308, 3.12776, 3.170407, 3.094292, 3.127037, 3.068026, 
    3.074315, 3.085734, 3.112121, 3.097838, 3.11455, 3.077795, 3.058943, 
    3.054086, 3.045054, 3.054293, 3.05354, 3.06241, 3.059556, 3.080961, 
    3.06944, 3.10231, 3.114417, 3.148926, 3.170324, 3.191691, 3.201143, 
    3.204026, 3.205233,
  3.255258, 3.278733, 3.274146, 3.293253, 3.282629, 3.295176, 3.259992, 
    3.279673, 3.267084, 3.257358, 3.330445, 3.29411, 3.368219, 3.344928, 
    3.404013, 3.364576, 3.41207, 3.402861, 3.430716, 3.422692, 3.458801, 
    3.434431, 3.477803, 3.45295, 3.456816, 3.433633, 3.301454, 3.32597, 
    3.299994, 3.303512, 3.301932, 3.282848, 3.273307, 3.253474, 3.257058, 
    3.271632, 3.305096, 3.293667, 3.322401, 3.321763, 3.353476, 3.339108, 
    3.393258, 3.377701, 3.423026, 3.41152, 3.422484, 3.419152, 3.422528, 
    3.405682, 3.412881, 3.398128, 3.341791, 3.358167, 3.309551, 3.280139, 
    3.260851, 3.247287, 3.249199, 3.252849, 3.271717, 3.289632, 3.303402, 
    3.312671, 3.321671, 3.348856, 3.363406, 3.396422, 3.390416, 3.4006, 
    3.410379, 3.426921, 3.424187, 3.431513, 3.400329, 3.420995, 3.387005, 
    3.396239, 3.324104, 3.296743, 3.285135, 3.275027, 3.25067, 3.267457, 
    3.260821, 3.276645, 3.286771, 3.281755, 3.312925, 3.300745, 3.364272, 
    3.336847, 3.409236, 3.391647, 3.413477, 3.402304, 3.421491, 3.404214, 
    3.434247, 3.440854, 3.436336, 3.453749, 3.403261, 3.422485, 3.281615, 
    3.282433, 3.286243, 3.269552, 3.268535, 3.253376, 3.266858, 3.27263, 
    3.287359, 3.296128, 3.304502, 3.322833, 3.34311, 3.37185, 3.392782, 
    3.406951, 3.398249, 3.40593, 3.397346, 3.393337, 3.438376, 3.412948, 
    3.451234, 3.449094, 3.431688, 3.449335, 3.283006, 3.278308, 3.262091, 
    3.27477, 3.251733, 3.264594, 3.27203, 3.301001, 3.307425, 3.313404, 
    3.324984, 3.339841, 3.366204, 3.389457, 3.410949, 3.409366, 3.409923, 
    3.414758, 3.402807, 3.416727, 3.419075, 3.412944, 3.448807, 3.438489, 
    3.449049, 3.442322, 3.279834, 3.287752, 3.283469, 3.291531, 3.285849, 
    3.311254, 3.318854, 3.354097, 3.339548, 3.362757, 3.341891, 3.345571, 
    3.363523, 3.343012, 3.388169, 3.357434, 3.414946, 3.383802, 3.416916, 
    3.410856, 3.420899, 3.429943, 3.441383, 3.462687, 3.457731, 3.47569, 
    3.299618, 3.310006, 3.309088, 3.319896, 3.327763, 3.344933, 3.372819, 
    3.362282, 3.381673, 3.385591, 3.356149, 3.374171, 3.316966, 3.326087, 
    3.32065, 3.300437, 3.364707, 3.331697, 3.393131, 3.374889, 3.428651, 
    3.401716, 3.455009, 3.478284, 3.500459, 3.526731, 3.315698, 3.308612, 
    3.321158, 3.338327, 3.354401, 3.375997, 3.37822, 3.3823, 3.39291, 
    3.40188, 3.383594, 3.404135, 3.328213, 3.3676, 3.305942, 3.324517, 
    3.33731, 3.331685, 3.361081, 3.36808, 3.396805, 3.381898, 3.472513, 
    3.431861, 3.546629, 3.514072, 3.306143, 3.315673, 3.348192, 3.332654, 
    3.377447, 3.388646, 3.397799, 3.409572, 3.410846, 3.417862, 3.406379, 
    3.417407, 3.376043, 3.39441, 3.344445, 3.356481, 3.350933, 3.344869, 
    3.363651, 3.383881, 3.384313, 3.39085, 3.409404, 3.37763, 3.477833, 
    3.415301, 3.32581, 3.343829, 3.346415, 3.339404, 3.38752, 3.369937, 
    3.417691, 3.404659, 3.42606, 3.415394, 3.41383, 3.400234, 3.391822, 
    3.37074, 3.353767, 3.340418, 3.343513, 3.358207, 3.385125, 3.410963, 
    3.405272, 3.424425, 3.374161, 3.395069, 3.38696, 3.40818, 3.362003, 
    3.401258, 3.352106, 3.356361, 3.36959, 3.396498, 3.402501, 3.408939, 
    3.404963, 3.385813, 3.382694, 3.369267, 3.365578, 3.355434, 3.34708, 
    3.354712, 3.362762, 3.38582, 3.406856, 3.430072, 3.435798, 3.463403, 
    3.440904, 3.478188, 3.446446, 3.501747, 3.403555, 3.445516, 3.370193, 
    3.378158, 3.392656, 3.42635, 3.408079, 3.429464, 3.382571, 3.358717, 
    3.352593, 3.341228, 3.352854, 3.351905, 3.363095, 3.359491, 3.38659, 
    3.371983, 3.413792, 3.429294, 3.473801, 3.501639, 3.530418, 3.543027, 
    3.546836, 3.548431,
  3.812406, 3.852937, 3.844965, 3.878337, 3.859726, 3.88172, 3.820528, 
    3.854572, 3.832743, 3.816005, 3.945441, 3.879844, 4.01692, 3.972602, 
    4.084903, 4.009935, 4.100404, 4.082694, 4.136674, 4.120997, 4.192388, 
    4.14397, 4.230848, 4.18067, 4.188406, 4.142401, 3.892799, 3.937109, 
    3.890218, 3.896441, 3.893644, 3.860109, 3.843509, 3.809353, 3.815492, 
    3.840606, 3.899248, 3.879065, 3.930483, 3.929301, 3.988774, 3.961651, 
    4.064368, 4.034976, 4.121648, 4.099342, 4.120593, 4.114115, 4.120677, 
    4.088106, 4.101969, 4.073643, 3.966693, 3.997694, 3.90716, 3.855384, 
    3.822005, 3.798792, 3.802051, 3.808284, 3.840755, 3.871978, 3.896246, 
    3.912715, 3.929131, 3.980019, 4.007696, 4.07039, 4.058971, 4.078366, 
    4.097143, 4.129248, 4.123912, 4.138238, 4.077848, 4.117695, 4.05251, 
    4.070041, 3.933642, 3.884481, 3.864103, 3.846494, 3.804561, 3.833386, 
    3.821953, 3.849304, 3.866965, 3.858202, 3.913168, 3.891545, 4.009353, 
    3.95741, 4.09494, 4.061307, 4.103121, 4.081628, 4.11866, 4.085288, 
    4.143606, 4.156633, 4.147718, 4.182268, 4.083461, 4.120595, 3.857958, 
    3.859383, 3.866041, 3.837007, 3.835249, 3.809186, 3.832352, 3.842335, 
    3.867995, 3.883397, 3.898195, 3.931285, 3.969176, 4.023901, 4.063463, 
    4.090544, 4.073875, 4.088581, 4.072153, 4.064517, 4.151739, 4.1021, 
    4.177247, 4.172982, 4.138582, 4.173461, 3.860385, 3.852197, 3.824137, 
    3.846049, 3.806376, 3.828447, 3.841297, 3.891997, 3.90338, 3.914023, 
    3.935276, 3.963027, 4.013053, 4.057154, 4.098242, 4.09519, 4.096264, 
    4.105598, 4.082592, 4.109411, 4.113965, 4.102093, 4.172411, 4.151962, 
    4.172891, 4.159538, 3.854853, 3.868683, 3.861193, 3.875312, 3.865352, 
    3.910191, 3.923916, 3.989954, 3.962476, 4.006454, 3.966881, 3.973815, 
    4.007919, 3.968991, 4.054713, 3.996299, 4.105962, 4.046459, 4.109776, 
    4.098062, 4.117509, 4.135159, 4.15768, 4.200201, 4.19024, 4.226542, 
    3.889555, 3.90797, 3.906336, 3.925843, 3.940444, 3.972611, 4.025769, 
    4.005546, 4.042445, 4.049838, 3.993853, 4.028357, 3.920427, 3.937326, 
    3.927238, 3.891, 4.010185, 3.947776, 4.064125, 4.029702, 4.13263, 
    4.080501, 4.184787, 4.231832, 4.277551, 4.33226, 3.918119, 3.905491, 
    3.92818, 3.960185, 3.99053, 4.031778, 4.03595, 4.043627, 4.063706, 
    4.080816, 4.046066, 4.085137, 3.941281, 4.015732, 3.900748, 3.93441, 
    3.958277, 3.947755, 4.003252, 4.016653, 4.07112, 4.042869, 4.220078, 
    4.138921, 4.374619, 4.306071, 3.901106, 3.918074, 3.978765, 3.949565, 
    4.034498, 4.055615, 4.073017, 4.095587, 4.098043, 4.111612, 4.089446, 
    4.110729, 4.031865, 4.066559, 3.971692, 3.994484, 3.983953, 3.972491, 
    4.008164, 4.046607, 4.047422, 4.059793, 4.095263, 4.034843, 4.23091, 
    4.10665, 3.936811, 3.97053, 3.975406, 3.962206, 4.053484, 4.020221, 
    4.111279, 4.086142, 4.127565, 4.106829, 4.103805, 4.077667, 4.061638, 
    4.021766, 3.989326, 3.964112, 3.969935, 3.99777, 4.048956, 4.098268, 
    4.087317, 4.124374, 4.028339, 4.067813, 4.052425, 4.092906, 4.005013, 
    4.079626, 3.986174, 3.994257, 4.019554, 4.070534, 4.082006, 4.094367, 
    4.086725, 4.050256, 4.044369, 4.018932, 4.011855, 3.992493, 3.976662, 
    3.991121, 4.006465, 4.050269, 4.09036, 4.135413, 4.146659, 4.201644, 
    4.156732, 4.231634, 4.167717, 4.280235, 4.084025, 4.165868, 4.020714, 
    4.035834, 4.063224, 4.128133, 4.092713, 4.134223, 4.044138, 3.998743, 
    3.987098, 3.965633, 3.987593, 3.985794, 4.007101, 4.000218, 4.051726, 
    4.024158, 4.10373, 4.133889, 4.222696, 4.280009, 4.33991, 4.366787, 
    4.37507, 4.378548,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24857.37, 24878.21, 24874.12, 24891.17, 24881.68, 24892.89, 24861.56, 
    24879.04, 24867.85, 24859.23, 24925, 24891.94, 24960.41, 24938.52, 
    24993.99, 24956.98, 25001.59, 24992.9, 25019.29, 25011.66, 25046.19, 
    25022.83, 25064.57, 25040.55, 25044.27, 25022.07, 24898.52, 24920.84, 
    24897.21, 24900.37, 24898.95, 24881.88, 24873.38, 24855.79, 24858.96, 
    24871.89, 24901.79, 24891.54, 24917.53, 24916.94, 24946.53, 24933.08, 
    24983.88, 24969.33, 25011.98, 25001.07, 25011.46, 25008.3, 25011.51, 
    24995.56, 25002.36, 24988.45, 24935.58, 24950.94, 24905.79, 24879.46, 
    24862.32, 24850.31, 24852, 24855.23, 24871.96, 24887.93, 24900.27, 
    24908.6, 24916.85, 24942.2, 24955.87, 24986.84, 24981.21, 24990.77, 
    24999.99, 25015.68, 25013.08, 25020.05, 24990.52, 25010.05, 24978.02, 
    24986.67, 24919.11, 24894.3, 24883.92, 24874.91, 24853.3, 24868.18, 
    24862.29, 24876.35, 24885.38, 24880.9, 24908.83, 24897.88, 24956.69, 
    24930.97, 24998.91, 24982.36, 25002.92, 24992.38, 25010.52, 24994.18, 
    25022.66, 25028.97, 25024.65, 25041.32, 24993.28, 25011.46, 24880.78, 
    24881.51, 24884.91, 24870.04, 24869.14, 24855.7, 24867.65, 24872.78, 
    24885.9, 24893.75, 24901.26, 24917.93, 24936.82, 24963.85, 24983.43, 
    24996.76, 24988.56, 24995.79, 24987.71, 24983.95, 25026.6, 25002.42, 
    25038.91, 25036.85, 25020.22, 25037.09, 24882.02, 24877.83, 24863.42, 
    24874.68, 24854.24, 24865.64, 24872.24, 24898.11, 24903.88, 24909.26, 
    24919.93, 24933.76, 24958.51, 24980.31, 25000.53, 24999.04, 24999.56, 
    25004.14, 24992.85, 25006, 25008.23, 25002.42, 25036.58, 25026.71, 
    25036.81, 25030.37, 24879.19, 24886.25, 24882.43, 24889.63, 24884.55, 
    24907.33, 24914.24, 24947.12, 24933.49, 24955.26, 24935.68, 24939.12, 
    24955.98, 24936.73, 24979.11, 24950.25, 25004.31, 24975.02, 25006.18, 
    25000.45, 25009.96, 25018.56, 25029.47, 25049.93, 25045.15, 25062.52, 
    24896.87, 24906.21, 24905.38, 24915.21, 24922.51, 24938.52, 24964.76, 
    24954.81, 24973.03, 24976.69, 24949.04, 24966.04, 24912.49, 24920.95, 
    24915.91, 24897.61, 24957.1, 24926.17, 24983.75, 24966.71, 25017.33, 
    24991.82, 25042.54, 25065.04, 25086.72, 25112.48, 24911.33, 24904.95, 
    24916.38, 24932.35, 24947.4, 24967.74, 24969.81, 24973.62, 24983.55, 
    24991.98, 24974.83, 24994.1, 24922.93, 24959.83, 24902.55, 24919.49, 
    24931.4, 24926.16, 24953.68, 24960.28, 24987.21, 24973.24, 25059.44, 
    25020.38, 25132.31, 25100.13, 24902.73, 24911.31, 24941.57, 24927.06, 
    24969.09, 24979.55, 24988.14, 24999.23, 25000.44, 25007.08, 24996.22, 
    25006.65, 24967.78, 24984.96, 24938.07, 24949.35, 24944.14, 24938.46, 
    24956.1, 24975.09, 24975.5, 24981.62, 24999.07, 24969.26, 25064.6, 
    25004.65, 24920.7, 24937.49, 24939.91, 24933.36, 24978.5, 24962.04, 
    25006.92, 24994.6, 25014.86, 25004.74, 25003.26, 24990.43, 24982.53, 
    24962.8, 24946.8, 24934.3, 24937.2, 24950.98, 24976.26, 25000.55, 
    24995.17, 25013.31, 24966.03, 24985.57, 24977.97, 24997.92, 24954.55, 
    24991.39, 24945.24, 24949.24, 24961.71, 24986.92, 24992.56, 24998.63, 
    24994.88, 24976.9, 24973.98, 24961.4, 24957.92, 24948.37, 24940.53, 
    24947.69, 24955.27, 24976.91, 24996.67, 25018.68, 25024.14, 25050.62, 
    25029.01, 25064.95, 25034.32, 25087.99, 24993.56, 25033.43, 24962.28, 
    24969.75, 24983.31, 25015.14, 24997.82, 25018.1, 24973.87, 24951.46, 
    24945.7, 24935.06, 24945.95, 24945.06, 24955.58, 24952.19, 24977.63, 
    24963.97, 25003.22, 25017.94, 25060.69, 25087.88, 25116.09, 25128.67, 
    25132.52, 25134.14 ;

 HCSOI =
  24857.37, 24878.21, 24874.12, 24891.17, 24881.68, 24892.89, 24861.56, 
    24879.04, 24867.85, 24859.23, 24925, 24891.94, 24960.41, 24938.52, 
    24993.99, 24956.98, 25001.59, 24992.9, 25019.29, 25011.66, 25046.19, 
    25022.83, 25064.57, 25040.55, 25044.27, 25022.07, 24898.52, 24920.84, 
    24897.21, 24900.37, 24898.95, 24881.88, 24873.38, 24855.79, 24858.96, 
    24871.89, 24901.79, 24891.54, 24917.53, 24916.94, 24946.53, 24933.08, 
    24983.88, 24969.33, 25011.98, 25001.07, 25011.46, 25008.3, 25011.51, 
    24995.56, 25002.36, 24988.45, 24935.58, 24950.94, 24905.79, 24879.46, 
    24862.32, 24850.31, 24852, 24855.23, 24871.96, 24887.93, 24900.27, 
    24908.6, 24916.85, 24942.2, 24955.87, 24986.84, 24981.21, 24990.77, 
    24999.99, 25015.68, 25013.08, 25020.05, 24990.52, 25010.05, 24978.02, 
    24986.67, 24919.11, 24894.3, 24883.92, 24874.91, 24853.3, 24868.18, 
    24862.29, 24876.35, 24885.38, 24880.9, 24908.83, 24897.88, 24956.69, 
    24930.97, 24998.91, 24982.36, 25002.92, 24992.38, 25010.52, 24994.18, 
    25022.66, 25028.97, 25024.65, 25041.32, 24993.28, 25011.46, 24880.78, 
    24881.51, 24884.91, 24870.04, 24869.14, 24855.7, 24867.65, 24872.78, 
    24885.9, 24893.75, 24901.26, 24917.93, 24936.82, 24963.85, 24983.43, 
    24996.76, 24988.56, 24995.79, 24987.71, 24983.95, 25026.6, 25002.42, 
    25038.91, 25036.85, 25020.22, 25037.09, 24882.02, 24877.83, 24863.42, 
    24874.68, 24854.24, 24865.64, 24872.24, 24898.11, 24903.88, 24909.26, 
    24919.93, 24933.76, 24958.51, 24980.31, 25000.53, 24999.04, 24999.56, 
    25004.14, 24992.85, 25006, 25008.23, 25002.42, 25036.58, 25026.71, 
    25036.81, 25030.37, 24879.19, 24886.25, 24882.43, 24889.63, 24884.55, 
    24907.33, 24914.24, 24947.12, 24933.49, 24955.26, 24935.68, 24939.12, 
    24955.98, 24936.73, 24979.11, 24950.25, 25004.31, 24975.02, 25006.18, 
    25000.45, 25009.96, 25018.56, 25029.47, 25049.93, 25045.15, 25062.52, 
    24896.87, 24906.21, 24905.38, 24915.21, 24922.51, 24938.52, 24964.76, 
    24954.81, 24973.03, 24976.69, 24949.04, 24966.04, 24912.49, 24920.95, 
    24915.91, 24897.61, 24957.1, 24926.17, 24983.75, 24966.71, 25017.33, 
    24991.82, 25042.54, 25065.04, 25086.72, 25112.48, 24911.33, 24904.95, 
    24916.38, 24932.35, 24947.4, 24967.74, 24969.81, 24973.62, 24983.55, 
    24991.98, 24974.83, 24994.1, 24922.93, 24959.83, 24902.55, 24919.49, 
    24931.4, 24926.16, 24953.68, 24960.28, 24987.21, 24973.24, 25059.44, 
    25020.38, 25132.31, 25100.13, 24902.73, 24911.31, 24941.57, 24927.06, 
    24969.09, 24979.55, 24988.14, 24999.23, 25000.44, 25007.08, 24996.22, 
    25006.65, 24967.78, 24984.96, 24938.07, 24949.35, 24944.14, 24938.46, 
    24956.1, 24975.09, 24975.5, 24981.62, 24999.07, 24969.26, 25064.6, 
    25004.65, 24920.7, 24937.49, 24939.91, 24933.36, 24978.5, 24962.04, 
    25006.92, 24994.6, 25014.86, 25004.74, 25003.26, 24990.43, 24982.53, 
    24962.8, 24946.8, 24934.3, 24937.2, 24950.98, 24976.26, 25000.55, 
    24995.17, 25013.31, 24966.03, 24985.57, 24977.97, 24997.92, 24954.55, 
    24991.39, 24945.24, 24949.24, 24961.71, 24986.92, 24992.56, 24998.63, 
    24994.88, 24976.9, 24973.98, 24961.4, 24957.92, 24948.37, 24940.53, 
    24947.69, 24955.27, 24976.91, 24996.67, 25018.68, 25024.14, 25050.62, 
    25029.01, 25064.95, 25034.32, 25087.99, 24993.56, 25033.43, 24962.28, 
    24969.75, 24983.31, 25015.14, 24997.82, 25018.1, 24973.87, 24951.46, 
    24945.7, 24935.06, 24945.95, 24945.06, 24955.58, 24952.19, 24977.63, 
    24963.97, 25003.22, 25017.94, 25060.69, 25087.88, 25116.09, 25128.67, 
    25132.52, 25134.14 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.191079e-08, 6.218382e-08, 6.213074e-08, 6.235096e-08, 6.22288e-08, 
    6.2373e-08, 6.196615e-08, 6.219464e-08, 6.204878e-08, 6.193537e-08, 
    6.277832e-08, 6.236078e-08, 6.321213e-08, 6.294581e-08, 6.361488e-08, 
    6.317068e-08, 6.370446e-08, 6.360209e-08, 6.391026e-08, 6.382197e-08, 
    6.421612e-08, 6.395101e-08, 6.442048e-08, 6.415281e-08, 6.419468e-08, 
    6.394226e-08, 6.244482e-08, 6.272633e-08, 6.242814e-08, 6.246828e-08, 
    6.245027e-08, 6.223132e-08, 6.212098e-08, 6.188993e-08, 6.193188e-08, 
    6.210158e-08, 6.248633e-08, 6.235573e-08, 6.268491e-08, 6.267748e-08, 
    6.304396e-08, 6.287872e-08, 6.349475e-08, 6.331966e-08, 6.382565e-08, 
    6.369839e-08, 6.381968e-08, 6.378291e-08, 6.382015e-08, 6.363351e-08, 
    6.371348e-08, 6.354926e-08, 6.290966e-08, 6.309762e-08, 6.253705e-08, 
    6.219999e-08, 6.197617e-08, 6.181733e-08, 6.183978e-08, 6.188259e-08, 
    6.210257e-08, 6.230942e-08, 6.246706e-08, 6.25725e-08, 6.267641e-08, 
    6.299089e-08, 6.315737e-08, 6.353015e-08, 6.346289e-08, 6.357685e-08, 
    6.368574e-08, 6.386854e-08, 6.383846e-08, 6.391899e-08, 6.357385e-08, 
    6.380323e-08, 6.342457e-08, 6.352813e-08, 6.270461e-08, 6.239097e-08, 
    6.225762e-08, 6.214094e-08, 6.185705e-08, 6.20531e-08, 6.197581e-08, 
    6.215969e-08, 6.227652e-08, 6.221874e-08, 6.257539e-08, 6.243673e-08, 
    6.316724e-08, 6.285257e-08, 6.367303e-08, 6.34767e-08, 6.37201e-08, 
    6.35959e-08, 6.380871e-08, 6.361718e-08, 6.394897e-08, 6.402121e-08, 
    6.397185e-08, 6.416151e-08, 6.360656e-08, 6.381967e-08, 6.221712e-08, 
    6.222654e-08, 6.227045e-08, 6.207744e-08, 6.206563e-08, 6.188878e-08, 
    6.204615e-08, 6.211316e-08, 6.22833e-08, 6.238393e-08, 6.247959e-08, 
    6.268994e-08, 6.292485e-08, 6.325337e-08, 6.348942e-08, 6.364765e-08, 
    6.355063e-08, 6.363629e-08, 6.354053e-08, 6.349565e-08, 6.399414e-08, 
    6.371423e-08, 6.413423e-08, 6.411099e-08, 6.392091e-08, 6.411361e-08, 
    6.223316e-08, 6.217893e-08, 6.199063e-08, 6.213799e-08, 6.186952e-08, 
    6.201979e-08, 6.210619e-08, 6.243962e-08, 6.251289e-08, 6.258082e-08, 
    6.271499e-08, 6.288717e-08, 6.318925e-08, 6.34521e-08, 6.369208e-08, 
    6.367449e-08, 6.368068e-08, 6.373428e-08, 6.36015e-08, 6.375608e-08, 
    6.378202e-08, 6.37142e-08, 6.410788e-08, 6.39954e-08, 6.411049e-08, 
    6.403727e-08, 6.219656e-08, 6.228781e-08, 6.22385e-08, 6.233122e-08, 
    6.22659e-08, 6.255637e-08, 6.264347e-08, 6.305104e-08, 6.288379e-08, 
    6.315e-08, 6.291083e-08, 6.295321e-08, 6.315866e-08, 6.292376e-08, 
    6.34376e-08, 6.30892e-08, 6.373637e-08, 6.338842e-08, 6.375817e-08, 
    6.369104e-08, 6.38022e-08, 6.390175e-08, 6.402701e-08, 6.425812e-08, 
    6.420461e-08, 6.43979e-08, 6.242386e-08, 6.254222e-08, 6.253181e-08, 
    6.265568e-08, 6.27473e-08, 6.294588e-08, 6.326439e-08, 6.314462e-08, 
    6.336451e-08, 6.340865e-08, 6.307459e-08, 6.327969e-08, 6.262145e-08, 
    6.272778e-08, 6.266447e-08, 6.243319e-08, 6.31722e-08, 6.279292e-08, 
    6.349332e-08, 6.328784e-08, 6.388755e-08, 6.358929e-08, 6.417515e-08, 
    6.442559e-08, 6.466136e-08, 6.493683e-08, 6.260683e-08, 6.25264e-08, 
    6.267042e-08, 6.286966e-08, 6.305456e-08, 6.330037e-08, 6.332552e-08, 
    6.337157e-08, 6.349087e-08, 6.359117e-08, 6.338612e-08, 6.361631e-08, 
    6.275242e-08, 6.320513e-08, 6.249599e-08, 6.27095e-08, 6.285792e-08, 
    6.279282e-08, 6.313093e-08, 6.321061e-08, 6.353445e-08, 6.336705e-08, 
    6.436377e-08, 6.392277e-08, 6.514664e-08, 6.480458e-08, 6.24983e-08, 
    6.260656e-08, 6.298333e-08, 6.280406e-08, 6.331678e-08, 6.3443e-08, 
    6.354561e-08, 6.367676e-08, 6.369093e-08, 6.376864e-08, 6.364129e-08, 
    6.376361e-08, 6.33009e-08, 6.350767e-08, 6.294027e-08, 6.307836e-08, 
    6.301484e-08, 6.294515e-08, 6.316022e-08, 6.338935e-08, 6.339426e-08, 
    6.346773e-08, 6.367474e-08, 6.331886e-08, 6.442066e-08, 6.374017e-08, 
    6.272461e-08, 6.293312e-08, 6.296292e-08, 6.288214e-08, 6.343034e-08, 
    6.32317e-08, 6.376674e-08, 6.362214e-08, 6.385908e-08, 6.374134e-08, 
    6.372401e-08, 6.35728e-08, 6.347865e-08, 6.32408e-08, 6.30473e-08, 
    6.289386e-08, 6.292954e-08, 6.309808e-08, 6.340337e-08, 6.36922e-08, 
    6.362893e-08, 6.384107e-08, 6.327961e-08, 6.351502e-08, 6.342403e-08, 
    6.36613e-08, 6.314143e-08, 6.358408e-08, 6.302828e-08, 6.307702e-08, 
    6.322776e-08, 6.353098e-08, 6.359809e-08, 6.366972e-08, 6.362552e-08, 
    6.341112e-08, 6.337601e-08, 6.322409e-08, 6.318215e-08, 6.306641e-08, 
    6.297058e-08, 6.305813e-08, 6.315008e-08, 6.341122e-08, 6.364657e-08, 
    6.390317e-08, 6.396598e-08, 6.426577e-08, 6.402171e-08, 6.442445e-08, 
    6.408201e-08, 6.467483e-08, 6.360975e-08, 6.407196e-08, 6.323462e-08, 
    6.332483e-08, 6.348797e-08, 6.386221e-08, 6.366019e-08, 6.389647e-08, 
    6.337463e-08, 6.310389e-08, 6.303387e-08, 6.290318e-08, 6.303685e-08, 
    6.302598e-08, 6.315389e-08, 6.311279e-08, 6.341989e-08, 6.325493e-08, 
    6.372358e-08, 6.38946e-08, 6.437764e-08, 6.467376e-08, 6.497525e-08, 
    6.510835e-08, 6.514885e-08, 6.516579e-08 ;

 HR_vr =
  2.673277e-07, 2.680603e-07, 2.67918e-07, 2.685084e-07, 2.68181e-07, 
    2.685675e-07, 2.674764e-07, 2.680892e-07, 2.676981e-07, 2.673938e-07, 
    2.696528e-07, 2.685347e-07, 2.708139e-07, 2.701017e-07, 2.718901e-07, 
    2.70703e-07, 2.721294e-07, 2.718562e-07, 2.726789e-07, 2.724433e-07, 
    2.73494e-07, 2.727876e-07, 2.740387e-07, 2.733255e-07, 2.73437e-07, 
    2.727642e-07, 2.687601e-07, 2.695135e-07, 2.687154e-07, 2.688229e-07, 
    2.687747e-07, 2.681877e-07, 2.678915e-07, 2.672719e-07, 2.673845e-07, 
    2.678397e-07, 2.688712e-07, 2.685214e-07, 2.694034e-07, 2.693835e-07, 
    2.703644e-07, 2.699223e-07, 2.715695e-07, 2.711017e-07, 2.724531e-07, 
    2.721134e-07, 2.724371e-07, 2.72339e-07, 2.724384e-07, 2.719401e-07, 
    2.721536e-07, 2.717152e-07, 2.70005e-07, 2.705079e-07, 2.690072e-07, 
    2.681033e-07, 2.675032e-07, 2.670769e-07, 2.671372e-07, 2.67252e-07, 
    2.678423e-07, 2.683972e-07, 2.688198e-07, 2.691023e-07, 2.693806e-07, 
    2.702219e-07, 2.706675e-07, 2.716639e-07, 2.714845e-07, 2.717887e-07, 
    2.720796e-07, 2.725675e-07, 2.724873e-07, 2.727021e-07, 2.717809e-07, 
    2.723931e-07, 2.713821e-07, 2.716587e-07, 2.694553e-07, 2.686158e-07, 
    2.682579e-07, 2.679453e-07, 2.671835e-07, 2.677096e-07, 2.675022e-07, 
    2.679957e-07, 2.68309e-07, 2.681541e-07, 2.6911e-07, 2.687385e-07, 
    2.706939e-07, 2.698521e-07, 2.720457e-07, 2.715213e-07, 2.721714e-07, 
    2.718398e-07, 2.724078e-07, 2.718966e-07, 2.727821e-07, 2.729747e-07, 
    2.72843e-07, 2.733489e-07, 2.718682e-07, 2.72437e-07, 2.681497e-07, 
    2.68175e-07, 2.682928e-07, 2.677749e-07, 2.677432e-07, 2.672687e-07, 
    2.676911e-07, 2.678708e-07, 2.683272e-07, 2.685969e-07, 2.688533e-07, 
    2.694168e-07, 2.700455e-07, 2.709243e-07, 2.715553e-07, 2.71978e-07, 
    2.717189e-07, 2.719476e-07, 2.716919e-07, 2.71572e-07, 2.729024e-07, 
    2.721556e-07, 2.732761e-07, 2.732142e-07, 2.727071e-07, 2.732212e-07, 
    2.681927e-07, 2.680473e-07, 2.675421e-07, 2.679375e-07, 2.67217e-07, 
    2.676203e-07, 2.67852e-07, 2.68746e-07, 2.689426e-07, 2.691245e-07, 
    2.694839e-07, 2.699449e-07, 2.707529e-07, 2.714555e-07, 2.720966e-07, 
    2.720496e-07, 2.720662e-07, 2.722092e-07, 2.718547e-07, 2.722674e-07, 
    2.723366e-07, 2.721556e-07, 2.732059e-07, 2.72906e-07, 2.732129e-07, 
    2.730176e-07, 2.680946e-07, 2.683393e-07, 2.682071e-07, 2.684556e-07, 
    2.682804e-07, 2.690589e-07, 2.692921e-07, 2.703831e-07, 2.699358e-07, 
    2.706479e-07, 2.700082e-07, 2.701215e-07, 2.706707e-07, 2.700428e-07, 
    2.714166e-07, 2.704851e-07, 2.722148e-07, 2.71285e-07, 2.72273e-07, 
    2.720938e-07, 2.723905e-07, 2.726561e-07, 2.729903e-07, 2.736062e-07, 
    2.734637e-07, 2.739787e-07, 2.68704e-07, 2.69021e-07, 2.689933e-07, 
    2.693251e-07, 2.695704e-07, 2.70102e-07, 2.709538e-07, 2.706337e-07, 
    2.712216e-07, 2.713395e-07, 2.704464e-07, 2.709947e-07, 2.692333e-07, 
    2.695179e-07, 2.693486e-07, 2.687289e-07, 2.707072e-07, 2.696924e-07, 
    2.715657e-07, 2.710166e-07, 2.726182e-07, 2.718219e-07, 2.733851e-07, 
    2.74052e-07, 2.746801e-07, 2.754124e-07, 2.691942e-07, 2.689788e-07, 
    2.693646e-07, 2.698978e-07, 2.703927e-07, 2.710501e-07, 2.711174e-07, 
    2.712404e-07, 2.715592e-07, 2.718271e-07, 2.712791e-07, 2.718943e-07, 
    2.695835e-07, 2.707953e-07, 2.688972e-07, 2.694689e-07, 2.698665e-07, 
    2.696923e-07, 2.705971e-07, 2.708102e-07, 2.716755e-07, 2.712284e-07, 
    2.738873e-07, 2.727119e-07, 2.759702e-07, 2.750608e-07, 2.689035e-07, 
    2.691935e-07, 2.702021e-07, 2.697224e-07, 2.71094e-07, 2.714312e-07, 
    2.717055e-07, 2.720556e-07, 2.720935e-07, 2.723009e-07, 2.71961e-07, 
    2.722875e-07, 2.710514e-07, 2.716041e-07, 2.700871e-07, 2.704564e-07, 
    2.702866e-07, 2.701001e-07, 2.706755e-07, 2.712877e-07, 2.713011e-07, 
    2.714973e-07, 2.720493e-07, 2.710996e-07, 2.740383e-07, 2.722241e-07, 
    2.695097e-07, 2.700675e-07, 2.701476e-07, 2.699315e-07, 2.713974e-07, 
    2.708665e-07, 2.722959e-07, 2.719098e-07, 2.725423e-07, 2.72228e-07, 
    2.721818e-07, 2.717781e-07, 2.715265e-07, 2.708908e-07, 2.703733e-07, 
    2.699629e-07, 2.700583e-07, 2.705091e-07, 2.713252e-07, 2.720968e-07, 
    2.719278e-07, 2.724943e-07, 2.709946e-07, 2.716236e-07, 2.713805e-07, 
    2.720144e-07, 2.706251e-07, 2.718074e-07, 2.703226e-07, 2.704529e-07, 
    2.70856e-07, 2.71666e-07, 2.718456e-07, 2.720368e-07, 2.719189e-07, 
    2.71346e-07, 2.712522e-07, 2.708462e-07, 2.70734e-07, 2.704246e-07, 
    2.701682e-07, 2.704024e-07, 2.706481e-07, 2.713464e-07, 2.719749e-07, 
    2.726598e-07, 2.728275e-07, 2.736261e-07, 2.729756e-07, 2.740484e-07, 
    2.731358e-07, 2.747152e-07, 2.718763e-07, 2.731096e-07, 2.708744e-07, 
    2.711155e-07, 2.715512e-07, 2.725503e-07, 2.720114e-07, 2.726418e-07, 
    2.712486e-07, 2.705245e-07, 2.703375e-07, 2.699878e-07, 2.703455e-07, 
    2.703164e-07, 2.706585e-07, 2.705486e-07, 2.713695e-07, 2.709287e-07, 
    2.721806e-07, 2.726369e-07, 2.739246e-07, 2.747128e-07, 2.755149e-07, 
    2.758686e-07, 2.759762e-07, 2.760212e-07,
  2.332861e-07, 2.341672e-07, 2.33996e-07, 2.347061e-07, 2.343123e-07, 
    2.347771e-07, 2.334648e-07, 2.34202e-07, 2.337316e-07, 2.333655e-07, 
    2.360823e-07, 2.347378e-07, 2.374777e-07, 2.366216e-07, 2.387709e-07, 
    2.373444e-07, 2.390583e-07, 2.3873e-07, 2.397183e-07, 2.394353e-07, 
    2.406978e-07, 2.398489e-07, 2.413518e-07, 2.404952e-07, 2.406292e-07, 
    2.398208e-07, 2.350087e-07, 2.35915e-07, 2.349549e-07, 2.350842e-07, 
    2.350262e-07, 2.343204e-07, 2.339643e-07, 2.332188e-07, 2.333542e-07, 
    2.339019e-07, 2.351424e-07, 2.347216e-07, 2.357821e-07, 2.357581e-07, 
    2.369373e-07, 2.364058e-07, 2.383855e-07, 2.378233e-07, 2.394471e-07, 
    2.39039e-07, 2.394279e-07, 2.3931e-07, 2.394295e-07, 2.388308e-07, 
    2.390873e-07, 2.385605e-07, 2.365053e-07, 2.371097e-07, 2.353058e-07, 
    2.342192e-07, 2.334972e-07, 2.329844e-07, 2.330569e-07, 2.331951e-07, 
    2.339051e-07, 2.345723e-07, 2.350804e-07, 2.354201e-07, 2.357547e-07, 
    2.367663e-07, 2.373017e-07, 2.384991e-07, 2.382833e-07, 2.38649e-07, 
    2.389984e-07, 2.395846e-07, 2.394881e-07, 2.397462e-07, 2.386394e-07, 
    2.393751e-07, 2.381603e-07, 2.384927e-07, 2.35845e-07, 2.348351e-07, 
    2.34405e-07, 2.340289e-07, 2.331126e-07, 2.337454e-07, 2.33496e-07, 
    2.340894e-07, 2.344662e-07, 2.342799e-07, 2.354294e-07, 2.349826e-07, 
    2.373334e-07, 2.363216e-07, 2.389577e-07, 2.383276e-07, 2.391086e-07, 
    2.387102e-07, 2.393927e-07, 2.387785e-07, 2.398423e-07, 2.400737e-07, 
    2.399156e-07, 2.405231e-07, 2.387444e-07, 2.394278e-07, 2.342746e-07, 
    2.34305e-07, 2.344466e-07, 2.33824e-07, 2.337859e-07, 2.332151e-07, 
    2.337231e-07, 2.339392e-07, 2.344881e-07, 2.348124e-07, 2.351207e-07, 
    2.357982e-07, 2.365541e-07, 2.376103e-07, 2.383684e-07, 2.388762e-07, 
    2.385649e-07, 2.388398e-07, 2.385325e-07, 2.383885e-07, 2.39987e-07, 
    2.390897e-07, 2.404358e-07, 2.403614e-07, 2.397524e-07, 2.403698e-07, 
    2.343264e-07, 2.341515e-07, 2.335439e-07, 2.340194e-07, 2.331529e-07, 
    2.33638e-07, 2.339167e-07, 2.349918e-07, 2.35228e-07, 2.354468e-07, 
    2.358789e-07, 2.36433e-07, 2.374043e-07, 2.382486e-07, 2.390187e-07, 
    2.389623e-07, 2.389822e-07, 2.391541e-07, 2.387281e-07, 2.39224e-07, 
    2.393072e-07, 2.390897e-07, 2.403514e-07, 2.399911e-07, 2.403598e-07, 
    2.401252e-07, 2.342083e-07, 2.345026e-07, 2.343436e-07, 2.346425e-07, 
    2.344319e-07, 2.35368e-07, 2.356485e-07, 2.369599e-07, 2.364221e-07, 
    2.372781e-07, 2.365091e-07, 2.366454e-07, 2.373057e-07, 2.365507e-07, 
    2.382019e-07, 2.370825e-07, 2.391608e-07, 2.380439e-07, 2.392307e-07, 
    2.390154e-07, 2.393719e-07, 2.39691e-07, 2.400924e-07, 2.408323e-07, 
    2.406611e-07, 2.412797e-07, 2.349412e-07, 2.353224e-07, 2.35289e-07, 
    2.356879e-07, 2.359829e-07, 2.366219e-07, 2.376457e-07, 2.372609e-07, 
    2.379674e-07, 2.381091e-07, 2.370358e-07, 2.376948e-07, 2.355776e-07, 
    2.359199e-07, 2.357162e-07, 2.349712e-07, 2.373494e-07, 2.361296e-07, 
    2.383809e-07, 2.377211e-07, 2.396455e-07, 2.386888e-07, 2.405667e-07, 
    2.41368e-07, 2.42122e-07, 2.430017e-07, 2.355306e-07, 2.352716e-07, 
    2.357354e-07, 2.363765e-07, 2.369713e-07, 2.377613e-07, 2.378422e-07, 
    2.3799e-07, 2.383731e-07, 2.38695e-07, 2.380367e-07, 2.387757e-07, 
    2.35999e-07, 2.374553e-07, 2.351735e-07, 2.35861e-07, 2.363388e-07, 
    2.361294e-07, 2.372169e-07, 2.37473e-07, 2.385129e-07, 2.379755e-07, 
    2.411702e-07, 2.397582e-07, 2.436712e-07, 2.425794e-07, 2.35181e-07, 
    2.355298e-07, 2.367422e-07, 2.361655e-07, 2.378141e-07, 2.382194e-07, 
    2.385488e-07, 2.389695e-07, 2.39015e-07, 2.392642e-07, 2.388558e-07, 
    2.392482e-07, 2.37763e-07, 2.38427e-07, 2.366039e-07, 2.370479e-07, 
    2.368437e-07, 2.366196e-07, 2.373111e-07, 2.38047e-07, 2.380629e-07, 
    2.382987e-07, 2.389626e-07, 2.378208e-07, 2.41352e-07, 2.391725e-07, 
    2.359099e-07, 2.365806e-07, 2.366766e-07, 2.364168e-07, 2.381787e-07, 
    2.375407e-07, 2.392582e-07, 2.387944e-07, 2.395543e-07, 2.391767e-07, 
    2.391212e-07, 2.386361e-07, 2.383339e-07, 2.375699e-07, 2.36948e-07, 
    2.364546e-07, 2.365693e-07, 2.371113e-07, 2.380921e-07, 2.390191e-07, 
    2.388161e-07, 2.394965e-07, 2.376946e-07, 2.384506e-07, 2.381584e-07, 
    2.3892e-07, 2.372506e-07, 2.386718e-07, 2.368869e-07, 2.370436e-07, 
    2.37528e-07, 2.385017e-07, 2.387172e-07, 2.38947e-07, 2.388053e-07, 
    2.38117e-07, 2.380042e-07, 2.375163e-07, 2.373815e-07, 2.370095e-07, 
    2.367013e-07, 2.369828e-07, 2.372783e-07, 2.381174e-07, 2.388727e-07, 
    2.396955e-07, 2.398968e-07, 2.408566e-07, 2.400751e-07, 2.41364e-07, 
    2.40268e-07, 2.421646e-07, 2.387544e-07, 2.402361e-07, 2.375501e-07, 
    2.378399e-07, 2.383637e-07, 2.395641e-07, 2.389164e-07, 2.396739e-07, 
    2.379999e-07, 2.371299e-07, 2.369049e-07, 2.364845e-07, 2.369145e-07, 
    2.368795e-07, 2.372907e-07, 2.371586e-07, 2.381452e-07, 2.376154e-07, 
    2.391197e-07, 2.39668e-07, 2.412148e-07, 2.421615e-07, 2.431245e-07, 
    2.435492e-07, 2.436784e-07, 2.437324e-07,
  2.190335e-07, 2.20003e-07, 2.198146e-07, 2.205963e-07, 2.201628e-07, 
    2.206745e-07, 2.192301e-07, 2.200415e-07, 2.195236e-07, 2.191208e-07, 
    2.221119e-07, 2.206312e-07, 2.236489e-07, 2.227056e-07, 2.250742e-07, 
    2.235021e-07, 2.25391e-07, 2.25029e-07, 2.261186e-07, 2.258066e-07, 
    2.271991e-07, 2.262626e-07, 2.279206e-07, 2.269756e-07, 2.271234e-07, 
    2.262317e-07, 2.209294e-07, 2.219276e-07, 2.208702e-07, 2.210126e-07, 
    2.209487e-07, 2.201717e-07, 2.197799e-07, 2.189594e-07, 2.191084e-07, 
    2.197111e-07, 2.210766e-07, 2.206133e-07, 2.217809e-07, 2.217545e-07, 
    2.230533e-07, 2.224679e-07, 2.246493e-07, 2.240296e-07, 2.258196e-07, 
    2.253696e-07, 2.257984e-07, 2.256684e-07, 2.258001e-07, 2.251402e-07, 
    2.25423e-07, 2.248421e-07, 2.225775e-07, 2.232434e-07, 2.212565e-07, 
    2.200604e-07, 2.192657e-07, 2.187014e-07, 2.187812e-07, 2.189333e-07, 
    2.197146e-07, 2.204489e-07, 2.210083e-07, 2.213823e-07, 2.217508e-07, 
    2.228652e-07, 2.23455e-07, 2.247745e-07, 2.245365e-07, 2.249397e-07, 
    2.253249e-07, 2.259712e-07, 2.258648e-07, 2.261495e-07, 2.249291e-07, 
    2.257403e-07, 2.24401e-07, 2.247674e-07, 2.218505e-07, 2.207383e-07, 
    2.20265e-07, 2.198508e-07, 2.188426e-07, 2.195389e-07, 2.192644e-07, 
    2.199174e-07, 2.203322e-07, 2.201271e-07, 2.213925e-07, 2.209007e-07, 
    2.234899e-07, 2.223752e-07, 2.252799e-07, 2.245854e-07, 2.254464e-07, 
    2.250071e-07, 2.257596e-07, 2.250824e-07, 2.262554e-07, 2.265107e-07, 
    2.263362e-07, 2.270063e-07, 2.250448e-07, 2.257984e-07, 2.201213e-07, 
    2.201547e-07, 2.203106e-07, 2.196253e-07, 2.195834e-07, 2.189553e-07, 
    2.195143e-07, 2.197522e-07, 2.203562e-07, 2.207133e-07, 2.210527e-07, 
    2.217987e-07, 2.226313e-07, 2.237949e-07, 2.246304e-07, 2.251902e-07, 
    2.24847e-07, 2.2515e-07, 2.248113e-07, 2.246525e-07, 2.26415e-07, 
    2.254256e-07, 2.269099e-07, 2.268279e-07, 2.261562e-07, 2.268371e-07, 
    2.201782e-07, 2.199857e-07, 2.193171e-07, 2.198404e-07, 2.188869e-07, 
    2.194206e-07, 2.197274e-07, 2.209108e-07, 2.211708e-07, 2.214117e-07, 
    2.218875e-07, 2.224979e-07, 2.235679e-07, 2.244984e-07, 2.253473e-07, 
    2.252851e-07, 2.25307e-07, 2.254965e-07, 2.250269e-07, 2.255736e-07, 
    2.256653e-07, 2.254255e-07, 2.268169e-07, 2.264195e-07, 2.268261e-07, 
    2.265674e-07, 2.200483e-07, 2.203722e-07, 2.201972e-07, 2.205263e-07, 
    2.202944e-07, 2.21325e-07, 2.216339e-07, 2.230784e-07, 2.224858e-07, 
    2.234289e-07, 2.225817e-07, 2.227318e-07, 2.234595e-07, 2.226275e-07, 
    2.24447e-07, 2.232135e-07, 2.255039e-07, 2.242729e-07, 2.25581e-07, 
    2.253436e-07, 2.257367e-07, 2.260885e-07, 2.265312e-07, 2.273474e-07, 
    2.271585e-07, 2.278409e-07, 2.20855e-07, 2.212748e-07, 2.21238e-07, 
    2.216773e-07, 2.220021e-07, 2.227059e-07, 2.23834e-07, 2.234099e-07, 
    2.241884e-07, 2.243446e-07, 2.231618e-07, 2.238881e-07, 2.215558e-07, 
    2.219328e-07, 2.217084e-07, 2.208881e-07, 2.235075e-07, 2.221637e-07, 
    2.246442e-07, 2.23917e-07, 2.260384e-07, 2.249837e-07, 2.270544e-07, 
    2.279385e-07, 2.287704e-07, 2.297416e-07, 2.21504e-07, 2.212188e-07, 
    2.217295e-07, 2.224357e-07, 2.230909e-07, 2.239613e-07, 2.240504e-07, 
    2.242134e-07, 2.246356e-07, 2.249904e-07, 2.242649e-07, 2.250793e-07, 
    2.220201e-07, 2.236241e-07, 2.211109e-07, 2.21868e-07, 2.223941e-07, 
    2.221634e-07, 2.233614e-07, 2.236436e-07, 2.247897e-07, 2.241974e-07, 
    2.277203e-07, 2.261628e-07, 2.304808e-07, 2.292754e-07, 2.211191e-07, 
    2.215031e-07, 2.228385e-07, 2.222033e-07, 2.240195e-07, 2.244661e-07, 
    2.248292e-07, 2.252931e-07, 2.253432e-07, 2.25618e-07, 2.251677e-07, 
    2.256002e-07, 2.239632e-07, 2.24695e-07, 2.22686e-07, 2.231752e-07, 
    2.229502e-07, 2.227033e-07, 2.234652e-07, 2.242762e-07, 2.242937e-07, 
    2.245536e-07, 2.252857e-07, 2.240268e-07, 2.27921e-07, 2.255171e-07, 
    2.219216e-07, 2.226606e-07, 2.227662e-07, 2.2248e-07, 2.244214e-07, 
    2.237182e-07, 2.256113e-07, 2.250999e-07, 2.259377e-07, 2.255215e-07, 
    2.254602e-07, 2.249254e-07, 2.245923e-07, 2.237504e-07, 2.230651e-07, 
    2.225216e-07, 2.22648e-07, 2.232451e-07, 2.243259e-07, 2.253477e-07, 
    2.251239e-07, 2.258741e-07, 2.238879e-07, 2.24721e-07, 2.24399e-07, 
    2.252384e-07, 2.233986e-07, 2.249651e-07, 2.229978e-07, 2.231705e-07, 
    2.237043e-07, 2.247774e-07, 2.250149e-07, 2.252682e-07, 2.251119e-07, 
    2.243533e-07, 2.242291e-07, 2.236913e-07, 2.235428e-07, 2.231329e-07, 
    2.227934e-07, 2.231036e-07, 2.234292e-07, 2.243537e-07, 2.251863e-07, 
    2.260935e-07, 2.263155e-07, 2.273743e-07, 2.265123e-07, 2.279344e-07, 
    2.267252e-07, 2.288178e-07, 2.25056e-07, 2.266899e-07, 2.237286e-07, 
    2.240479e-07, 2.246253e-07, 2.259487e-07, 2.252345e-07, 2.260698e-07, 
    2.242242e-07, 2.232656e-07, 2.230176e-07, 2.225546e-07, 2.230282e-07, 
    2.229897e-07, 2.234427e-07, 2.232972e-07, 2.243844e-07, 2.238005e-07, 
    2.254586e-07, 2.260632e-07, 2.277694e-07, 2.288141e-07, 2.29877e-07, 
    2.303459e-07, 2.304886e-07, 2.305483e-07,
  2.100144e-07, 2.110119e-07, 2.10818e-07, 2.116224e-07, 2.111762e-07, 
    2.11703e-07, 2.102167e-07, 2.110515e-07, 2.105186e-07, 2.101042e-07, 
    2.131833e-07, 2.116583e-07, 2.147672e-07, 2.137949e-07, 2.162373e-07, 
    2.146159e-07, 2.165642e-07, 2.161906e-07, 2.173151e-07, 2.16993e-07, 
    2.18431e-07, 2.174638e-07, 2.191764e-07, 2.182001e-07, 2.183528e-07, 
    2.174319e-07, 2.119653e-07, 2.129935e-07, 2.119044e-07, 2.12051e-07, 
    2.119852e-07, 2.111854e-07, 2.107823e-07, 2.099382e-07, 2.100914e-07, 
    2.107115e-07, 2.121169e-07, 2.116399e-07, 2.128422e-07, 2.12815e-07, 
    2.141532e-07, 2.135499e-07, 2.157988e-07, 2.151597e-07, 2.170064e-07, 
    2.16542e-07, 2.169846e-07, 2.168504e-07, 2.169863e-07, 2.163053e-07, 
    2.165971e-07, 2.159977e-07, 2.136629e-07, 2.143491e-07, 2.123022e-07, 
    2.11071e-07, 2.102533e-07, 2.096729e-07, 2.097549e-07, 2.099113e-07, 
    2.107151e-07, 2.114707e-07, 2.120465e-07, 2.124317e-07, 2.128111e-07, 
    2.139595e-07, 2.145673e-07, 2.15928e-07, 2.156825e-07, 2.160984e-07, 
    2.164958e-07, 2.171629e-07, 2.170531e-07, 2.17347e-07, 2.160875e-07, 
    2.169246e-07, 2.155427e-07, 2.159207e-07, 2.129141e-07, 2.117686e-07, 
    2.112815e-07, 2.108553e-07, 2.09818e-07, 2.105343e-07, 2.10252e-07, 
    2.109237e-07, 2.113506e-07, 2.111395e-07, 2.124422e-07, 2.119357e-07, 
    2.146033e-07, 2.134544e-07, 2.164495e-07, 2.157329e-07, 2.166212e-07, 
    2.16168e-07, 2.169446e-07, 2.162456e-07, 2.174564e-07, 2.1772e-07, 
    2.175398e-07, 2.182318e-07, 2.162069e-07, 2.169846e-07, 2.111336e-07, 
    2.11168e-07, 2.113284e-07, 2.106233e-07, 2.105801e-07, 2.09934e-07, 
    2.10509e-07, 2.107538e-07, 2.113753e-07, 2.117429e-07, 2.120923e-07, 
    2.128605e-07, 2.137184e-07, 2.149178e-07, 2.157794e-07, 2.163568e-07, 
    2.160027e-07, 2.163154e-07, 2.159659e-07, 2.158021e-07, 2.176212e-07, 
    2.165998e-07, 2.181323e-07, 2.180475e-07, 2.17354e-07, 2.18057e-07, 
    2.111921e-07, 2.10994e-07, 2.103061e-07, 2.108445e-07, 2.098636e-07, 
    2.104127e-07, 2.107283e-07, 2.119463e-07, 2.122139e-07, 2.12462e-07, 
    2.12952e-07, 2.135808e-07, 2.146837e-07, 2.156432e-07, 2.16519e-07, 
    2.164548e-07, 2.164774e-07, 2.16673e-07, 2.161884e-07, 2.167526e-07, 
    2.168472e-07, 2.165997e-07, 2.180361e-07, 2.176258e-07, 2.180457e-07, 
    2.177785e-07, 2.110584e-07, 2.113918e-07, 2.112117e-07, 2.115504e-07, 
    2.113117e-07, 2.123728e-07, 2.126908e-07, 2.141791e-07, 2.135684e-07, 
    2.145404e-07, 2.136671e-07, 2.138219e-07, 2.14572e-07, 2.137143e-07, 
    2.155902e-07, 2.143184e-07, 2.166806e-07, 2.154107e-07, 2.167602e-07, 
    2.165152e-07, 2.169208e-07, 2.172841e-07, 2.177411e-07, 2.185842e-07, 
    2.18389e-07, 2.190941e-07, 2.118887e-07, 2.123211e-07, 2.12283e-07, 
    2.127354e-07, 2.1307e-07, 2.137951e-07, 2.14958e-07, 2.145207e-07, 
    2.153234e-07, 2.154845e-07, 2.14265e-07, 2.150138e-07, 2.126104e-07, 
    2.129987e-07, 2.127675e-07, 2.119228e-07, 2.146214e-07, 2.132366e-07, 
    2.157936e-07, 2.150436e-07, 2.172323e-07, 2.161439e-07, 2.182815e-07, 
    2.191951e-07, 2.200549e-07, 2.210594e-07, 2.12557e-07, 2.122633e-07, 
    2.127892e-07, 2.135168e-07, 2.141919e-07, 2.150893e-07, 2.151811e-07, 
    2.153492e-07, 2.157846e-07, 2.161507e-07, 2.154023e-07, 2.162424e-07, 
    2.130887e-07, 2.147416e-07, 2.121522e-07, 2.12932e-07, 2.13474e-07, 
    2.132362e-07, 2.144707e-07, 2.147617e-07, 2.159437e-07, 2.153327e-07, 
    2.189696e-07, 2.173608e-07, 2.218242e-07, 2.205772e-07, 2.121606e-07, 
    2.12556e-07, 2.139319e-07, 2.132773e-07, 2.151492e-07, 2.156099e-07, 
    2.159844e-07, 2.164631e-07, 2.165148e-07, 2.167984e-07, 2.163336e-07, 
    2.1678e-07, 2.150912e-07, 2.15846e-07, 2.137747e-07, 2.142788e-07, 
    2.140469e-07, 2.137925e-07, 2.145777e-07, 2.154141e-07, 2.15432e-07, 
    2.157002e-07, 2.164557e-07, 2.151568e-07, 2.191771e-07, 2.166945e-07, 
    2.129871e-07, 2.137485e-07, 2.138573e-07, 2.135624e-07, 2.155637e-07, 
    2.148386e-07, 2.167914e-07, 2.162637e-07, 2.171284e-07, 2.166987e-07, 
    2.166355e-07, 2.160837e-07, 2.1574e-07, 2.148719e-07, 2.141654e-07, 
    2.136052e-07, 2.137354e-07, 2.143508e-07, 2.154653e-07, 2.165194e-07, 
    2.162885e-07, 2.170627e-07, 2.150135e-07, 2.158728e-07, 2.155407e-07, 
    2.164067e-07, 2.145091e-07, 2.161249e-07, 2.14096e-07, 2.142739e-07, 
    2.148242e-07, 2.159311e-07, 2.16176e-07, 2.164374e-07, 2.162761e-07, 
    2.154936e-07, 2.153654e-07, 2.148109e-07, 2.146577e-07, 2.142352e-07, 
    2.138853e-07, 2.14205e-07, 2.145406e-07, 2.154939e-07, 2.163529e-07, 
    2.172893e-07, 2.175184e-07, 2.186122e-07, 2.177218e-07, 2.19191e-07, 
    2.179418e-07, 2.201041e-07, 2.162186e-07, 2.179051e-07, 2.148493e-07, 
    2.151786e-07, 2.157741e-07, 2.171398e-07, 2.164026e-07, 2.172648e-07, 
    2.153604e-07, 2.143721e-07, 2.141164e-07, 2.136392e-07, 2.141273e-07, 
    2.140876e-07, 2.145546e-07, 2.144045e-07, 2.155256e-07, 2.149234e-07, 
    2.166339e-07, 2.17258e-07, 2.190202e-07, 2.201002e-07, 2.211994e-07, 
    2.216846e-07, 2.218323e-07, 2.218941e-07,
  2.030062e-07, 2.039531e-07, 2.037689e-07, 2.04533e-07, 2.041091e-07, 
    2.046095e-07, 2.031981e-07, 2.039907e-07, 2.034847e-07, 2.030914e-07, 
    2.060172e-07, 2.045671e-07, 2.07525e-07, 2.06599e-07, 2.089265e-07, 
    2.073809e-07, 2.092383e-07, 2.088818e-07, 2.099551e-07, 2.096475e-07, 
    2.110214e-07, 2.100971e-07, 2.117341e-07, 2.108006e-07, 2.109466e-07, 
    2.100666e-07, 2.048588e-07, 2.058366e-07, 2.048009e-07, 2.049403e-07, 
    2.048777e-07, 2.041179e-07, 2.037351e-07, 2.029339e-07, 2.030793e-07, 
    2.036678e-07, 2.050029e-07, 2.045496e-07, 2.056924e-07, 2.056666e-07, 
    2.069401e-07, 2.063658e-07, 2.085082e-07, 2.078989e-07, 2.096604e-07, 
    2.092171e-07, 2.096395e-07, 2.095114e-07, 2.096412e-07, 2.089913e-07, 
    2.092697e-07, 2.086979e-07, 2.064733e-07, 2.071267e-07, 2.05179e-07, 
    2.040093e-07, 2.032329e-07, 2.026822e-07, 2.0276e-07, 2.029085e-07, 
    2.036713e-07, 2.043888e-07, 2.04936e-07, 2.053021e-07, 2.056629e-07, 
    2.067558e-07, 2.073346e-07, 2.086314e-07, 2.083973e-07, 2.08794e-07, 
    2.091731e-07, 2.098098e-07, 2.09705e-07, 2.099856e-07, 2.087835e-07, 
    2.095823e-07, 2.082639e-07, 2.086244e-07, 2.057611e-07, 2.046718e-07, 
    2.042092e-07, 2.038043e-07, 2.028199e-07, 2.034997e-07, 2.032317e-07, 
    2.038693e-07, 2.042747e-07, 2.040742e-07, 2.053121e-07, 2.048307e-07, 
    2.073689e-07, 2.06275e-07, 2.091288e-07, 2.084453e-07, 2.092927e-07, 
    2.088602e-07, 2.096014e-07, 2.089343e-07, 2.1009e-07, 2.103418e-07, 
    2.101697e-07, 2.108308e-07, 2.088974e-07, 2.096395e-07, 2.040686e-07, 
    2.041013e-07, 2.042536e-07, 2.035841e-07, 2.035431e-07, 2.029299e-07, 
    2.034755e-07, 2.03708e-07, 2.042982e-07, 2.046474e-07, 2.049795e-07, 
    2.057099e-07, 2.065262e-07, 2.076684e-07, 2.084896e-07, 2.090404e-07, 
    2.087026e-07, 2.090009e-07, 2.086675e-07, 2.085113e-07, 2.102474e-07, 
    2.092723e-07, 2.107357e-07, 2.106547e-07, 2.099922e-07, 2.106638e-07, 
    2.041242e-07, 2.039361e-07, 2.03283e-07, 2.037941e-07, 2.028631e-07, 
    2.033841e-07, 2.036838e-07, 2.048408e-07, 2.050951e-07, 2.053309e-07, 
    2.057969e-07, 2.063952e-07, 2.074454e-07, 2.083598e-07, 2.091951e-07, 
    2.091339e-07, 2.091554e-07, 2.093421e-07, 2.088798e-07, 2.09418e-07, 
    2.095084e-07, 2.092722e-07, 2.106438e-07, 2.102518e-07, 2.10653e-07, 
    2.103977e-07, 2.039972e-07, 2.043138e-07, 2.041428e-07, 2.044645e-07, 
    2.042378e-07, 2.052462e-07, 2.055486e-07, 2.069648e-07, 2.063834e-07, 
    2.073089e-07, 2.064774e-07, 2.066247e-07, 2.073391e-07, 2.065223e-07, 
    2.083094e-07, 2.070975e-07, 2.093494e-07, 2.081383e-07, 2.094253e-07, 
    2.091915e-07, 2.095786e-07, 2.099255e-07, 2.10362e-07, 2.111678e-07, 
    2.109811e-07, 2.116553e-07, 2.04786e-07, 2.05197e-07, 2.051608e-07, 
    2.055909e-07, 2.059092e-07, 2.065992e-07, 2.077066e-07, 2.072901e-07, 
    2.080549e-07, 2.082085e-07, 2.070466e-07, 2.077599e-07, 2.05472e-07, 
    2.058414e-07, 2.056215e-07, 2.048184e-07, 2.073861e-07, 2.060677e-07, 
    2.085032e-07, 2.077882e-07, 2.09876e-07, 2.088373e-07, 2.108784e-07, 
    2.11752e-07, 2.125747e-07, 2.13537e-07, 2.054213e-07, 2.05142e-07, 
    2.056421e-07, 2.063344e-07, 2.06977e-07, 2.078318e-07, 2.079193e-07, 
    2.080795e-07, 2.084946e-07, 2.088438e-07, 2.081302e-07, 2.089313e-07, 
    2.059272e-07, 2.075006e-07, 2.050364e-07, 2.05778e-07, 2.062935e-07, 
    2.060673e-07, 2.072425e-07, 2.075196e-07, 2.086464e-07, 2.080638e-07, 
    2.115363e-07, 2.099988e-07, 2.142701e-07, 2.130749e-07, 2.050444e-07, 
    2.054203e-07, 2.067294e-07, 2.061064e-07, 2.078889e-07, 2.083281e-07, 
    2.086852e-07, 2.091418e-07, 2.091911e-07, 2.094618e-07, 2.090183e-07, 
    2.094442e-07, 2.078337e-07, 2.085531e-07, 2.065797e-07, 2.070597e-07, 
    2.068389e-07, 2.065967e-07, 2.073444e-07, 2.081415e-07, 2.081585e-07, 
    2.084142e-07, 2.091351e-07, 2.078961e-07, 2.11735e-07, 2.093629e-07, 
    2.058303e-07, 2.065549e-07, 2.066584e-07, 2.063776e-07, 2.08284e-07, 
    2.075929e-07, 2.094552e-07, 2.089516e-07, 2.097768e-07, 2.093667e-07, 
    2.093064e-07, 2.087798e-07, 2.084521e-07, 2.076246e-07, 2.069517e-07, 
    2.064184e-07, 2.065424e-07, 2.071283e-07, 2.081902e-07, 2.091956e-07, 
    2.089753e-07, 2.09714e-07, 2.077596e-07, 2.085788e-07, 2.082621e-07, 
    2.09088e-07, 2.07279e-07, 2.088194e-07, 2.068856e-07, 2.07055e-07, 
    2.075792e-07, 2.086344e-07, 2.088679e-07, 2.091173e-07, 2.089634e-07, 
    2.082172e-07, 2.08095e-07, 2.075665e-07, 2.074206e-07, 2.070181e-07, 
    2.06685e-07, 2.069894e-07, 2.073091e-07, 2.082175e-07, 2.090367e-07, 
    2.099304e-07, 2.101492e-07, 2.111946e-07, 2.103436e-07, 2.117482e-07, 
    2.10554e-07, 2.12622e-07, 2.089087e-07, 2.105188e-07, 2.076031e-07, 
    2.079169e-07, 2.084847e-07, 2.097878e-07, 2.090841e-07, 2.099071e-07, 
    2.080902e-07, 2.071486e-07, 2.06905e-07, 2.064508e-07, 2.069154e-07, 
    2.068776e-07, 2.073223e-07, 2.071794e-07, 2.082477e-07, 2.076737e-07, 
    2.093048e-07, 2.099006e-07, 2.115846e-07, 2.126181e-07, 2.13671e-07, 
    2.141362e-07, 2.142778e-07, 2.14337e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.191079e-08, 6.218382e-08, 6.213074e-08, 6.235096e-08, 6.22288e-08, 
    6.2373e-08, 6.196615e-08, 6.219464e-08, 6.204878e-08, 6.193537e-08, 
    6.277832e-08, 6.236078e-08, 6.321213e-08, 6.294581e-08, 6.361488e-08, 
    6.317068e-08, 6.370446e-08, 6.360209e-08, 6.391026e-08, 6.382197e-08, 
    6.421612e-08, 6.395101e-08, 6.442048e-08, 6.415281e-08, 6.419468e-08, 
    6.394226e-08, 6.244482e-08, 6.272633e-08, 6.242814e-08, 6.246828e-08, 
    6.245027e-08, 6.223132e-08, 6.212098e-08, 6.188993e-08, 6.193188e-08, 
    6.210158e-08, 6.248633e-08, 6.235573e-08, 6.268491e-08, 6.267748e-08, 
    6.304396e-08, 6.287872e-08, 6.349475e-08, 6.331966e-08, 6.382565e-08, 
    6.369839e-08, 6.381968e-08, 6.378291e-08, 6.382015e-08, 6.363351e-08, 
    6.371348e-08, 6.354926e-08, 6.290966e-08, 6.309762e-08, 6.253705e-08, 
    6.219999e-08, 6.197617e-08, 6.181733e-08, 6.183978e-08, 6.188259e-08, 
    6.210257e-08, 6.230942e-08, 6.246706e-08, 6.25725e-08, 6.267641e-08, 
    6.299089e-08, 6.315737e-08, 6.353015e-08, 6.346289e-08, 6.357685e-08, 
    6.368574e-08, 6.386854e-08, 6.383846e-08, 6.391899e-08, 6.357385e-08, 
    6.380323e-08, 6.342457e-08, 6.352813e-08, 6.270461e-08, 6.239097e-08, 
    6.225762e-08, 6.214094e-08, 6.185705e-08, 6.20531e-08, 6.197581e-08, 
    6.215969e-08, 6.227652e-08, 6.221874e-08, 6.257539e-08, 6.243673e-08, 
    6.316724e-08, 6.285257e-08, 6.367303e-08, 6.34767e-08, 6.37201e-08, 
    6.35959e-08, 6.380871e-08, 6.361718e-08, 6.394897e-08, 6.402121e-08, 
    6.397185e-08, 6.416151e-08, 6.360656e-08, 6.381967e-08, 6.221712e-08, 
    6.222654e-08, 6.227045e-08, 6.207744e-08, 6.206563e-08, 6.188878e-08, 
    6.204615e-08, 6.211316e-08, 6.22833e-08, 6.238393e-08, 6.247959e-08, 
    6.268994e-08, 6.292485e-08, 6.325337e-08, 6.348942e-08, 6.364765e-08, 
    6.355063e-08, 6.363629e-08, 6.354053e-08, 6.349565e-08, 6.399414e-08, 
    6.371423e-08, 6.413423e-08, 6.411099e-08, 6.392091e-08, 6.411361e-08, 
    6.223316e-08, 6.217893e-08, 6.199063e-08, 6.213799e-08, 6.186952e-08, 
    6.201979e-08, 6.210619e-08, 6.243962e-08, 6.251289e-08, 6.258082e-08, 
    6.271499e-08, 6.288717e-08, 6.318925e-08, 6.34521e-08, 6.369208e-08, 
    6.367449e-08, 6.368068e-08, 6.373428e-08, 6.36015e-08, 6.375608e-08, 
    6.378202e-08, 6.37142e-08, 6.410788e-08, 6.39954e-08, 6.411049e-08, 
    6.403727e-08, 6.219656e-08, 6.228781e-08, 6.22385e-08, 6.233122e-08, 
    6.22659e-08, 6.255637e-08, 6.264347e-08, 6.305104e-08, 6.288379e-08, 
    6.315e-08, 6.291083e-08, 6.295321e-08, 6.315866e-08, 6.292376e-08, 
    6.34376e-08, 6.30892e-08, 6.373637e-08, 6.338842e-08, 6.375817e-08, 
    6.369104e-08, 6.38022e-08, 6.390175e-08, 6.402701e-08, 6.425812e-08, 
    6.420461e-08, 6.43979e-08, 6.242386e-08, 6.254222e-08, 6.253181e-08, 
    6.265568e-08, 6.27473e-08, 6.294588e-08, 6.326439e-08, 6.314462e-08, 
    6.336451e-08, 6.340865e-08, 6.307459e-08, 6.327969e-08, 6.262145e-08, 
    6.272778e-08, 6.266447e-08, 6.243319e-08, 6.31722e-08, 6.279292e-08, 
    6.349332e-08, 6.328784e-08, 6.388755e-08, 6.358929e-08, 6.417515e-08, 
    6.442559e-08, 6.466136e-08, 6.493683e-08, 6.260683e-08, 6.25264e-08, 
    6.267042e-08, 6.286966e-08, 6.305456e-08, 6.330037e-08, 6.332552e-08, 
    6.337157e-08, 6.349087e-08, 6.359117e-08, 6.338612e-08, 6.361631e-08, 
    6.275242e-08, 6.320513e-08, 6.249599e-08, 6.27095e-08, 6.285792e-08, 
    6.279282e-08, 6.313093e-08, 6.321061e-08, 6.353445e-08, 6.336705e-08, 
    6.436377e-08, 6.392277e-08, 6.514664e-08, 6.480458e-08, 6.24983e-08, 
    6.260656e-08, 6.298333e-08, 6.280406e-08, 6.331678e-08, 6.3443e-08, 
    6.354561e-08, 6.367676e-08, 6.369093e-08, 6.376864e-08, 6.364129e-08, 
    6.376361e-08, 6.33009e-08, 6.350767e-08, 6.294027e-08, 6.307836e-08, 
    6.301484e-08, 6.294515e-08, 6.316022e-08, 6.338935e-08, 6.339426e-08, 
    6.346773e-08, 6.367474e-08, 6.331886e-08, 6.442066e-08, 6.374017e-08, 
    6.272461e-08, 6.293312e-08, 6.296292e-08, 6.288214e-08, 6.343034e-08, 
    6.32317e-08, 6.376674e-08, 6.362214e-08, 6.385908e-08, 6.374134e-08, 
    6.372401e-08, 6.35728e-08, 6.347865e-08, 6.32408e-08, 6.30473e-08, 
    6.289386e-08, 6.292954e-08, 6.309808e-08, 6.340337e-08, 6.36922e-08, 
    6.362893e-08, 6.384107e-08, 6.327961e-08, 6.351502e-08, 6.342403e-08, 
    6.36613e-08, 6.314143e-08, 6.358408e-08, 6.302828e-08, 6.307702e-08, 
    6.322776e-08, 6.353098e-08, 6.359809e-08, 6.366972e-08, 6.362552e-08, 
    6.341112e-08, 6.337601e-08, 6.322409e-08, 6.318215e-08, 6.306641e-08, 
    6.297058e-08, 6.305813e-08, 6.315008e-08, 6.341122e-08, 6.364657e-08, 
    6.390317e-08, 6.396598e-08, 6.426577e-08, 6.402171e-08, 6.442445e-08, 
    6.408201e-08, 6.467483e-08, 6.360975e-08, 6.407196e-08, 6.323462e-08, 
    6.332483e-08, 6.348797e-08, 6.386221e-08, 6.366019e-08, 6.389647e-08, 
    6.337463e-08, 6.310389e-08, 6.303387e-08, 6.290318e-08, 6.303685e-08, 
    6.302598e-08, 6.315389e-08, 6.311279e-08, 6.341989e-08, 6.325493e-08, 
    6.372358e-08, 6.38946e-08, 6.437764e-08, 6.467376e-08, 6.497525e-08, 
    6.510835e-08, 6.514885e-08, 6.516579e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.578916e-13, 9.605178e-13, 9.600076e-13, 9.621242e-13, 9.609506e-13, 
    9.62336e-13, 9.584246e-13, 9.606217e-13, 9.592195e-13, 9.581287e-13, 
    9.662267e-13, 9.622187e-13, 9.703888e-13, 9.678357e-13, 9.742465e-13, 
    9.699911e-13, 9.75104e-13, 9.741248e-13, 9.770735e-13, 9.762291e-13, 
    9.799954e-13, 9.774631e-13, 9.819474e-13, 9.793914e-13, 9.797909e-13, 
    9.773793e-13, 9.630265e-13, 9.657276e-13, 9.628662e-13, 9.632516e-13, 
    9.630789e-13, 9.609745e-13, 9.599129e-13, 9.576915e-13, 9.58095e-13, 
    9.59727e-13, 9.634249e-13, 9.621707e-13, 9.653326e-13, 9.652612e-13, 
    9.687773e-13, 9.671925e-13, 9.730971e-13, 9.714202e-13, 9.762643e-13, 
    9.750466e-13, 9.76207e-13, 9.758552e-13, 9.762115e-13, 9.744256e-13, 
    9.751908e-13, 9.736191e-13, 9.674891e-13, 9.692916e-13, 9.639123e-13, 
    9.606722e-13, 9.585208e-13, 9.569927e-13, 9.572087e-13, 9.576205e-13, 
    9.597364e-13, 9.617256e-13, 9.632404e-13, 9.642532e-13, 9.65251e-13, 
    9.682667e-13, 9.698639e-13, 9.734356e-13, 9.727922e-13, 9.738828e-13, 
    9.749255e-13, 9.766743e-13, 9.763866e-13, 9.771566e-13, 9.738547e-13, 
    9.760492e-13, 9.724254e-13, 9.734169e-13, 9.655189e-13, 9.625093e-13, 
    9.612264e-13, 9.601056e-13, 9.573748e-13, 9.592607e-13, 9.585173e-13, 
    9.602862e-13, 9.614093e-13, 9.608541e-13, 9.64281e-13, 9.629489e-13, 
    9.699585e-13, 9.669412e-13, 9.748039e-13, 9.729243e-13, 9.752544e-13, 
    9.740658e-13, 9.761018e-13, 9.742695e-13, 9.774434e-13, 9.781337e-13, 
    9.77662e-13, 9.79475e-13, 9.741678e-13, 9.762066e-13, 9.608384e-13, 
    9.609289e-13, 9.613511e-13, 9.594947e-13, 9.593813e-13, 9.576802e-13, 
    9.591942e-13, 9.598384e-13, 9.614747e-13, 9.624416e-13, 9.633607e-13, 
    9.653806e-13, 9.676344e-13, 9.707844e-13, 9.730462e-13, 9.745611e-13, 
    9.736325e-13, 9.744523e-13, 9.735357e-13, 9.731061e-13, 9.778749e-13, 
    9.751978e-13, 9.792142e-13, 9.789923e-13, 9.771748e-13, 9.790172e-13, 
    9.609926e-13, 9.604713e-13, 9.586601e-13, 9.600776e-13, 9.574949e-13, 
    9.589405e-13, 9.597711e-13, 9.629761e-13, 9.636806e-13, 9.643328e-13, 
    9.656211e-13, 9.672736e-13, 9.7017e-13, 9.726885e-13, 9.749864e-13, 
    9.748181e-13, 9.748773e-13, 9.7539e-13, 9.741193e-13, 9.755986e-13, 
    9.758466e-13, 9.751979e-13, 9.789625e-13, 9.778875e-13, 9.789875e-13, 
    9.782877e-13, 9.606409e-13, 9.615179e-13, 9.61044e-13, 9.61935e-13, 
    9.61307e-13, 9.640975e-13, 9.649336e-13, 9.688445e-13, 9.672408e-13, 
    9.697936e-13, 9.675005e-13, 9.679067e-13, 9.698754e-13, 9.676246e-13, 
    9.725491e-13, 9.692101e-13, 9.7541e-13, 9.720773e-13, 9.756186e-13, 
    9.749764e-13, 9.7604e-13, 9.769918e-13, 9.781895e-13, 9.803973e-13, 
    9.798863e-13, 9.817323e-13, 9.628253e-13, 9.639619e-13, 9.638625e-13, 
    9.650518e-13, 9.659311e-13, 9.678368e-13, 9.708903e-13, 9.697426e-13, 
    9.7185e-13, 9.722726e-13, 9.690713e-13, 9.710366e-13, 9.647228e-13, 
    9.65743e-13, 9.651361e-13, 9.629146e-13, 9.700063e-13, 9.663684e-13, 
    9.730834e-13, 9.711151e-13, 9.768561e-13, 9.740017e-13, 9.79605e-13, 
    9.819954e-13, 9.842463e-13, 9.868711e-13, 9.645827e-13, 9.638105e-13, 
    9.651934e-13, 9.671048e-13, 9.688789e-13, 9.712351e-13, 9.714765e-13, 
    9.719174e-13, 9.730602e-13, 9.740205e-13, 9.720563e-13, 9.742611e-13, 
    9.659784e-13, 9.703221e-13, 9.63518e-13, 9.655675e-13, 9.669924e-13, 
    9.66368e-13, 9.696115e-13, 9.703754e-13, 9.734769e-13, 9.718743e-13, 
    9.814051e-13, 9.771921e-13, 9.8887e-13, 9.85611e-13, 9.635406e-13, 
    9.645803e-13, 9.681955e-13, 9.664759e-13, 9.713927e-13, 9.726014e-13, 
    9.735844e-13, 9.748393e-13, 9.749752e-13, 9.757185e-13, 9.745003e-13, 
    9.756707e-13, 9.712401e-13, 9.73221e-13, 9.677831e-13, 9.691072e-13, 
    9.684984e-13, 9.6783e-13, 9.698924e-13, 9.720871e-13, 9.721349e-13, 
    9.728381e-13, 9.748172e-13, 9.714126e-13, 9.819465e-13, 9.754437e-13, 
    9.657136e-13, 9.677134e-13, 9.680001e-13, 9.672254e-13, 9.724803e-13, 
    9.705771e-13, 9.757006e-13, 9.74317e-13, 9.765839e-13, 9.754576e-13, 
    9.752918e-13, 9.738446e-13, 9.729431e-13, 9.706642e-13, 9.688092e-13, 
    9.67338e-13, 9.676801e-13, 9.692961e-13, 9.722214e-13, 9.749871e-13, 
    9.743814e-13, 9.764118e-13, 9.710364e-13, 9.73291e-13, 9.724195e-13, 
    9.746917e-13, 9.697119e-13, 9.7395e-13, 9.686273e-13, 9.690946e-13, 
    9.705394e-13, 9.734432e-13, 9.740868e-13, 9.74772e-13, 9.743494e-13, 
    9.722959e-13, 9.719598e-13, 9.705045e-13, 9.70102e-13, 9.689929e-13, 
    9.680739e-13, 9.689133e-13, 9.697944e-13, 9.722971e-13, 9.745503e-13, 
    9.770053e-13, 9.776061e-13, 9.80469e-13, 9.781374e-13, 9.819825e-13, 
    9.787117e-13, 9.843724e-13, 9.741969e-13, 9.786174e-13, 9.706054e-13, 
    9.714698e-13, 9.730316e-13, 9.766128e-13, 9.746809e-13, 9.769405e-13, 
    9.719467e-13, 9.693514e-13, 9.686808e-13, 9.674272e-13, 9.687095e-13, 
    9.686052e-13, 9.698316e-13, 9.694376e-13, 9.723803e-13, 9.707999e-13, 
    9.752873e-13, 9.76923e-13, 9.815385e-13, 9.843636e-13, 9.872382e-13, 
    9.885058e-13, 9.888916e-13, 9.890528e-13 ;

 LITR1C =
  3.06688e-05, 3.066868e-05, 3.066871e-05, 3.066861e-05, 3.066866e-05, 
    3.06686e-05, 3.066878e-05, 3.066868e-05, 3.066874e-05, 3.066879e-05, 
    3.066842e-05, 3.066861e-05, 3.066824e-05, 3.066835e-05, 3.066806e-05, 
    3.066826e-05, 3.066802e-05, 3.066807e-05, 3.066794e-05, 3.066797e-05, 
    3.06678e-05, 3.066792e-05, 3.066771e-05, 3.066783e-05, 3.066781e-05, 
    3.066792e-05, 3.066857e-05, 3.066845e-05, 3.066858e-05, 3.066856e-05, 
    3.066857e-05, 3.066866e-05, 3.066871e-05, 3.066881e-05, 3.066879e-05, 
    3.066872e-05, 3.066855e-05, 3.066861e-05, 3.066847e-05, 3.066847e-05, 
    3.066831e-05, 3.066838e-05, 3.066811e-05, 3.066819e-05, 3.066797e-05, 
    3.066803e-05, 3.066798e-05, 3.066799e-05, 3.066798e-05, 3.066806e-05, 
    3.066802e-05, 3.066809e-05, 3.066837e-05, 3.066829e-05, 3.066853e-05, 
    3.066867e-05, 3.066877e-05, 3.066884e-05, 3.066883e-05, 3.066881e-05, 
    3.066872e-05, 3.066863e-05, 3.066856e-05, 3.066851e-05, 3.066847e-05, 
    3.066833e-05, 3.066826e-05, 3.06681e-05, 3.066813e-05, 3.066808e-05, 
    3.066803e-05, 3.066795e-05, 3.066796e-05, 3.066793e-05, 3.066808e-05, 
    3.066798e-05, 3.066815e-05, 3.06681e-05, 3.066846e-05, 3.066859e-05, 
    3.066865e-05, 3.06687e-05, 3.066882e-05, 3.066874e-05, 3.066877e-05, 
    3.066869e-05, 3.066864e-05, 3.066867e-05, 3.066851e-05, 3.066857e-05, 
    3.066826e-05, 3.066839e-05, 3.066804e-05, 3.066812e-05, 3.066802e-05, 
    3.066807e-05, 3.066798e-05, 3.066806e-05, 3.066792e-05, 3.066789e-05, 
    3.066791e-05, 3.066783e-05, 3.066807e-05, 3.066798e-05, 3.066867e-05, 
    3.066866e-05, 3.066865e-05, 3.066873e-05, 3.066873e-05, 3.066881e-05, 
    3.066874e-05, 3.066871e-05, 3.066864e-05, 3.066859e-05, 3.066855e-05, 
    3.066846e-05, 3.066836e-05, 3.066822e-05, 3.066812e-05, 3.066805e-05, 
    3.066809e-05, 3.066805e-05, 3.06681e-05, 3.066811e-05, 3.06679e-05, 
    3.066802e-05, 3.066784e-05, 3.066785e-05, 3.066793e-05, 3.066785e-05, 
    3.066866e-05, 3.066869e-05, 3.066877e-05, 3.06687e-05, 3.066882e-05, 
    3.066875e-05, 3.066872e-05, 3.066857e-05, 3.066854e-05, 3.066851e-05, 
    3.066845e-05, 3.066838e-05, 3.066825e-05, 3.066813e-05, 3.066803e-05, 
    3.066804e-05, 3.066803e-05, 3.066801e-05, 3.066807e-05, 3.0668e-05, 
    3.066799e-05, 3.066802e-05, 3.066785e-05, 3.06679e-05, 3.066785e-05, 
    3.066788e-05, 3.066868e-05, 3.066864e-05, 3.066866e-05, 3.066862e-05, 
    3.066865e-05, 3.066852e-05, 3.066848e-05, 3.066831e-05, 3.066838e-05, 
    3.066826e-05, 3.066837e-05, 3.066835e-05, 3.066826e-05, 3.066836e-05, 
    3.066814e-05, 3.066829e-05, 3.066801e-05, 3.066816e-05, 3.0668e-05, 
    3.066803e-05, 3.066798e-05, 3.066794e-05, 3.066788e-05, 3.066779e-05, 
    3.066781e-05, 3.066772e-05, 3.066858e-05, 3.066853e-05, 3.066853e-05, 
    3.066848e-05, 3.066844e-05, 3.066835e-05, 3.066822e-05, 3.066827e-05, 
    3.066817e-05, 3.066815e-05, 3.06683e-05, 3.066821e-05, 3.066849e-05, 
    3.066845e-05, 3.066847e-05, 3.066858e-05, 3.066826e-05, 3.066842e-05, 
    3.066811e-05, 3.06682e-05, 3.066795e-05, 3.066807e-05, 3.066782e-05, 
    3.066771e-05, 3.066761e-05, 3.066749e-05, 3.06685e-05, 3.066853e-05, 
    3.066847e-05, 3.066839e-05, 3.066831e-05, 3.06682e-05, 3.066819e-05, 
    3.066817e-05, 3.066812e-05, 3.066807e-05, 3.066816e-05, 3.066806e-05, 
    3.066844e-05, 3.066824e-05, 3.066855e-05, 3.066846e-05, 3.066839e-05, 
    3.066842e-05, 3.066827e-05, 3.066824e-05, 3.06681e-05, 3.066817e-05, 
    3.066774e-05, 3.066793e-05, 3.06674e-05, 3.066755e-05, 3.066855e-05, 
    3.06685e-05, 3.066834e-05, 3.066841e-05, 3.066819e-05, 3.066814e-05, 
    3.066809e-05, 3.066804e-05, 3.066803e-05, 3.0668e-05, 3.066805e-05, 
    3.0668e-05, 3.06682e-05, 3.066811e-05, 3.066835e-05, 3.06683e-05, 
    3.066832e-05, 3.066835e-05, 3.066826e-05, 3.066816e-05, 3.066816e-05, 
    3.066812e-05, 3.066804e-05, 3.066819e-05, 3.066771e-05, 3.066801e-05, 
    3.066845e-05, 3.066836e-05, 3.066834e-05, 3.066838e-05, 3.066814e-05, 
    3.066823e-05, 3.0668e-05, 3.066806e-05, 3.066796e-05, 3.066801e-05, 
    3.066802e-05, 3.066808e-05, 3.066812e-05, 3.066822e-05, 3.066831e-05, 
    3.066838e-05, 3.066836e-05, 3.066829e-05, 3.066815e-05, 3.066803e-05, 
    3.066806e-05, 3.066796e-05, 3.066821e-05, 3.066811e-05, 3.066815e-05, 
    3.066804e-05, 3.066827e-05, 3.066808e-05, 3.066832e-05, 3.06683e-05, 
    3.066823e-05, 3.06681e-05, 3.066807e-05, 3.066804e-05, 3.066806e-05, 
    3.066815e-05, 3.066816e-05, 3.066823e-05, 3.066825e-05, 3.06683e-05, 
    3.066834e-05, 3.06683e-05, 3.066826e-05, 3.066815e-05, 3.066805e-05, 
    3.066794e-05, 3.066791e-05, 3.066778e-05, 3.066789e-05, 3.066771e-05, 
    3.066786e-05, 3.06676e-05, 3.066807e-05, 3.066787e-05, 3.066823e-05, 
    3.066819e-05, 3.066812e-05, 3.066796e-05, 3.066804e-05, 3.066794e-05, 
    3.066816e-05, 3.066829e-05, 3.066831e-05, 3.066837e-05, 3.066831e-05, 
    3.066832e-05, 3.066826e-05, 3.066828e-05, 3.066815e-05, 3.066822e-05, 
    3.066802e-05, 3.066794e-05, 3.066773e-05, 3.06676e-05, 3.066748e-05, 
    3.066742e-05, 3.06674e-05, 3.066739e-05 ;

 LITR1C_TO_SOIL1C =
  6.37999e-13, 6.397478e-13, 6.394081e-13, 6.408175e-13, 6.40036e-13, 
    6.409586e-13, 6.38354e-13, 6.39817e-13, 6.388833e-13, 6.381569e-13, 
    6.435494e-13, 6.408805e-13, 6.463211e-13, 6.44621e-13, 6.4889e-13, 
    6.460563e-13, 6.49461e-13, 6.48809e-13, 6.507725e-13, 6.502102e-13, 
    6.527183e-13, 6.51032e-13, 6.540181e-13, 6.52316e-13, 6.525822e-13, 
    6.509762e-13, 6.414185e-13, 6.432171e-13, 6.413117e-13, 6.415683e-13, 
    6.414533e-13, 6.40052e-13, 6.39345e-13, 6.378657e-13, 6.381345e-13, 
    6.392212e-13, 6.416837e-13, 6.408485e-13, 6.429541e-13, 6.429066e-13, 
    6.45248e-13, 6.441926e-13, 6.481246e-13, 6.470079e-13, 6.502337e-13, 
    6.494228e-13, 6.501955e-13, 6.499613e-13, 6.501985e-13, 6.490093e-13, 
    6.495189e-13, 6.484722e-13, 6.443901e-13, 6.455905e-13, 6.420083e-13, 
    6.398506e-13, 6.38418e-13, 6.374004e-13, 6.375443e-13, 6.378184e-13, 
    6.392275e-13, 6.405521e-13, 6.415609e-13, 6.422353e-13, 6.428997e-13, 
    6.44908e-13, 6.459716e-13, 6.4835e-13, 6.479215e-13, 6.486478e-13, 
    6.493422e-13, 6.505067e-13, 6.503151e-13, 6.508279e-13, 6.48629e-13, 
    6.500905e-13, 6.476773e-13, 6.483376e-13, 6.430781e-13, 6.410739e-13, 
    6.402197e-13, 6.394733e-13, 6.376549e-13, 6.389107e-13, 6.384156e-13, 
    6.395936e-13, 6.403415e-13, 6.399717e-13, 6.422538e-13, 6.413668e-13, 
    6.460346e-13, 6.440253e-13, 6.492612e-13, 6.480095e-13, 6.495612e-13, 
    6.487697e-13, 6.501255e-13, 6.489053e-13, 6.510189e-13, 6.514786e-13, 
    6.511644e-13, 6.523717e-13, 6.488376e-13, 6.501953e-13, 6.399613e-13, 
    6.400216e-13, 6.403028e-13, 6.390665e-13, 6.38991e-13, 6.378583e-13, 
    6.388665e-13, 6.392955e-13, 6.40385e-13, 6.410289e-13, 6.416409e-13, 
    6.42986e-13, 6.444869e-13, 6.465846e-13, 6.480907e-13, 6.490995e-13, 
    6.484811e-13, 6.490271e-13, 6.484167e-13, 6.481306e-13, 6.513062e-13, 
    6.495235e-13, 6.521981e-13, 6.520502e-13, 6.5084e-13, 6.520669e-13, 
    6.40064e-13, 6.397169e-13, 6.385107e-13, 6.394547e-13, 6.377349e-13, 
    6.386974e-13, 6.392506e-13, 6.413848e-13, 6.41854e-13, 6.422883e-13, 
    6.431462e-13, 6.442466e-13, 6.461754e-13, 6.478525e-13, 6.493827e-13, 
    6.492706e-13, 6.4931e-13, 6.496515e-13, 6.488053e-13, 6.497904e-13, 
    6.499555e-13, 6.495235e-13, 6.520305e-13, 6.513146e-13, 6.520471e-13, 
    6.515811e-13, 6.398298e-13, 6.404138e-13, 6.400982e-13, 6.406915e-13, 
    6.402734e-13, 6.421316e-13, 6.426884e-13, 6.452927e-13, 6.442248e-13, 
    6.459247e-13, 6.443977e-13, 6.446682e-13, 6.459793e-13, 6.444804e-13, 
    6.477597e-13, 6.455362e-13, 6.496648e-13, 6.474456e-13, 6.498037e-13, 
    6.493761e-13, 6.500843e-13, 6.507182e-13, 6.515158e-13, 6.529859e-13, 
    6.526457e-13, 6.538749e-13, 6.412844e-13, 6.420413e-13, 6.419751e-13, 
    6.427671e-13, 6.433527e-13, 6.446217e-13, 6.466551e-13, 6.458908e-13, 
    6.472941e-13, 6.475756e-13, 6.454438e-13, 6.467525e-13, 6.42548e-13, 
    6.432274e-13, 6.428232e-13, 6.413439e-13, 6.460664e-13, 6.436438e-13, 
    6.481155e-13, 6.468048e-13, 6.506278e-13, 6.48727e-13, 6.524583e-13, 
    6.540501e-13, 6.55549e-13, 6.572969e-13, 6.424547e-13, 6.419405e-13, 
    6.428614e-13, 6.441342e-13, 6.453157e-13, 6.468847e-13, 6.470454e-13, 
    6.473391e-13, 6.481001e-13, 6.487395e-13, 6.474315e-13, 6.488998e-13, 
    6.433842e-13, 6.462767e-13, 6.417457e-13, 6.431105e-13, 6.440594e-13, 
    6.436436e-13, 6.458035e-13, 6.463122e-13, 6.483775e-13, 6.473103e-13, 
    6.53657e-13, 6.508515e-13, 6.58628e-13, 6.564578e-13, 6.417607e-13, 
    6.424531e-13, 6.448606e-13, 6.437155e-13, 6.469896e-13, 6.477946e-13, 
    6.484491e-13, 6.492848e-13, 6.493753e-13, 6.498703e-13, 6.49059e-13, 
    6.498384e-13, 6.46888e-13, 6.482071e-13, 6.44586e-13, 6.454677e-13, 
    6.450622e-13, 6.446172e-13, 6.459905e-13, 6.47452e-13, 6.474839e-13, 
    6.479522e-13, 6.492701e-13, 6.470029e-13, 6.540176e-13, 6.496872e-13, 
    6.432078e-13, 6.445395e-13, 6.447304e-13, 6.442146e-13, 6.477139e-13, 
    6.464465e-13, 6.498583e-13, 6.48937e-13, 6.504465e-13, 6.496965e-13, 
    6.495861e-13, 6.486224e-13, 6.48022e-13, 6.465046e-13, 6.452692e-13, 
    6.442895e-13, 6.445174e-13, 6.455935e-13, 6.475415e-13, 6.493832e-13, 
    6.489798e-13, 6.503319e-13, 6.467523e-13, 6.482537e-13, 6.476734e-13, 
    6.491864e-13, 6.458703e-13, 6.486925e-13, 6.451481e-13, 6.454593e-13, 
    6.464214e-13, 6.483551e-13, 6.487837e-13, 6.492399e-13, 6.489585e-13, 
    6.475911e-13, 6.473673e-13, 6.463981e-13, 6.461302e-13, 6.453916e-13, 
    6.447796e-13, 6.453386e-13, 6.459253e-13, 6.475919e-13, 6.490923e-13, 
    6.507271e-13, 6.511273e-13, 6.530336e-13, 6.51481e-13, 6.540415e-13, 
    6.518634e-13, 6.55633e-13, 6.488569e-13, 6.518007e-13, 6.464654e-13, 
    6.47041e-13, 6.48081e-13, 6.504657e-13, 6.491793e-13, 6.50684e-13, 
    6.473585e-13, 6.456303e-13, 6.451837e-13, 6.443489e-13, 6.452028e-13, 
    6.451334e-13, 6.459501e-13, 6.456877e-13, 6.476472e-13, 6.465949e-13, 
    6.495831e-13, 6.506723e-13, 6.537459e-13, 6.556272e-13, 6.575414e-13, 
    6.583855e-13, 6.586424e-13, 6.587497e-13 ;

 LITR1C_vr =
  0.00175122, 0.001751213, 0.001751215, 0.001751209, 0.001751212, 
    0.001751209, 0.001751219, 0.001751213, 0.001751217, 0.00175122, 
    0.001751199, 0.001751209, 0.001751188, 0.001751195, 0.001751178, 
    0.001751189, 0.001751176, 0.001751178, 0.001751171, 0.001751173, 
    0.001751163, 0.00175117, 0.001751158, 0.001751165, 0.001751164, 
    0.00175117, 0.001751207, 0.0017512, 0.001751207, 0.001751206, 
    0.001751207, 0.001751212, 0.001751215, 0.001751221, 0.00175122, 
    0.001751216, 0.001751206, 0.001751209, 0.001751201, 0.001751201, 
    0.001751192, 0.001751196, 0.001751181, 0.001751185, 0.001751173, 
    0.001751176, 0.001751173, 0.001751174, 0.001751173, 0.001751178, 
    0.001751176, 0.00175118, 0.001751196, 0.001751191, 0.001751205, 
    0.001751213, 0.001751219, 0.001751223, 0.001751222, 0.001751221, 
    0.001751215, 0.00175121, 0.001751206, 0.001751204, 0.001751201, 
    0.001751194, 0.001751189, 0.00175118, 0.001751182, 0.001751179, 
    0.001751176, 0.001751172, 0.001751173, 0.001751171, 0.001751179, 
    0.001751173, 0.001751183, 0.00175118, 0.001751201, 0.001751208, 
    0.001751212, 0.001751214, 0.001751222, 0.001751217, 0.001751219, 
    0.001751214, 0.001751211, 0.001751213, 0.001751204, 0.001751207, 
    0.001751189, 0.001751197, 0.001751177, 0.001751181, 0.001751175, 
    0.001751179, 0.001751173, 0.001751178, 0.00175117, 0.001751168, 
    0.001751169, 0.001751165, 0.001751178, 0.001751173, 0.001751213, 
    0.001751212, 0.001751211, 0.001751216, 0.001751216, 0.001751221, 
    0.001751217, 0.001751215, 0.001751211, 0.001751209, 0.001751206, 
    0.001751201, 0.001751195, 0.001751187, 0.001751181, 0.001751177, 
    0.00175118, 0.001751178, 0.00175118, 0.001751181, 0.001751169, 
    0.001751176, 0.001751165, 0.001751166, 0.00175117, 0.001751166, 
    0.001751212, 0.001751214, 0.001751218, 0.001751215, 0.001751221, 
    0.001751218, 0.001751215, 0.001751207, 0.001751205, 0.001751204, 
    0.0017512, 0.001751196, 0.001751189, 0.001751182, 0.001751176, 
    0.001751177, 0.001751176, 0.001751175, 0.001751178, 0.001751175, 
    0.001751174, 0.001751176, 0.001751166, 0.001751169, 0.001751166, 
    0.001751168, 0.001751213, 0.001751211, 0.001751212, 0.00175121, 
    0.001751211, 0.001751204, 0.001751202, 0.001751192, 0.001751196, 
    0.00175119, 0.001751196, 0.001751194, 0.001751189, 0.001751195, 
    0.001751182, 0.001751191, 0.001751175, 0.001751184, 0.001751175, 
    0.001751176, 0.001751173, 0.001751171, 0.001751168, 0.001751162, 
    0.001751164, 0.001751159, 0.001751208, 0.001751205, 0.001751205, 
    0.001751202, 0.001751199, 0.001751195, 0.001751187, 0.00175119, 
    0.001751184, 0.001751183, 0.001751191, 0.001751186, 0.001751203, 
    0.0017512, 0.001751202, 0.001751207, 0.001751189, 0.001751198, 
    0.001751181, 0.001751186, 0.001751171, 0.001751179, 0.001751164, 
    0.001751158, 0.001751152, 0.001751146, 0.001751203, 0.001751205, 
    0.001751201, 0.001751196, 0.001751192, 0.001751186, 0.001751185, 
    0.001751184, 0.001751181, 0.001751179, 0.001751184, 0.001751178, 
    0.001751199, 0.001751188, 0.001751206, 0.0017512, 0.001751197, 
    0.001751198, 0.00175119, 0.001751188, 0.00175118, 0.001751184, 
    0.00175116, 0.00175117, 0.00175114, 0.001751149, 0.001751206, 
    0.001751203, 0.001751194, 0.001751198, 0.001751185, 0.001751182, 
    0.00175118, 0.001751177, 0.001751176, 0.001751174, 0.001751177, 
    0.001751174, 0.001751186, 0.001751181, 0.001751195, 0.001751191, 
    0.001751193, 0.001751195, 0.001751189, 0.001751184, 0.001751184, 
    0.001751182, 0.001751177, 0.001751185, 0.001751158, 0.001751175, 
    0.0017512, 0.001751195, 0.001751194, 0.001751196, 0.001751183, 
    0.001751187, 0.001751174, 0.001751178, 0.001751172, 0.001751175, 
    0.001751175, 0.001751179, 0.001751181, 0.001751187, 0.001751192, 
    0.001751196, 0.001751195, 0.001751191, 0.001751183, 0.001751176, 
    0.001751178, 0.001751172, 0.001751186, 0.001751181, 0.001751183, 
    0.001751177, 0.00175119, 0.001751179, 0.001751193, 0.001751191, 
    0.001751188, 0.00175118, 0.001751179, 0.001751177, 0.001751178, 
    0.001751183, 0.001751184, 0.001751188, 0.001751189, 0.001751192, 
    0.001751194, 0.001751192, 0.00175119, 0.001751183, 0.001751177, 
    0.001751171, 0.001751169, 0.001751162, 0.001751168, 0.001751158, 
    0.001751167, 0.001751152, 0.001751178, 0.001751167, 0.001751187, 
    0.001751185, 0.001751181, 0.001751172, 0.001751177, 0.001751171, 
    0.001751184, 0.001751191, 0.001751192, 0.001751196, 0.001751192, 
    0.001751193, 0.001751189, 0.001751191, 0.001751183, 0.001751187, 
    0.001751175, 0.001751171, 0.001751159, 0.001751152, 0.001751145, 
    0.001751141, 0.00175114, 0.00175114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.733138e-07, 9.733101e-07, 9.733108e-07, 9.733078e-07, 9.733094e-07, 
    9.733075e-07, 9.73313e-07, 9.7331e-07, 9.733119e-07, 9.733135e-07, 
    9.733019e-07, 9.733076e-07, 9.732959e-07, 9.732996e-07, 9.732904e-07, 
    9.732964e-07, 9.732892e-07, 9.732905e-07, 9.732863e-07, 9.732876e-07, 
    9.732821e-07, 9.732858e-07, 9.732794e-07, 9.73283e-07, 9.732825e-07, 
    9.732859e-07, 9.733064e-07, 9.733026e-07, 9.733067e-07, 9.733061e-07, 
    9.733064e-07, 9.733094e-07, 9.733109e-07, 9.733141e-07, 9.733135e-07, 
    9.733112e-07, 9.733059e-07, 9.733077e-07, 9.733031e-07, 9.733033e-07, 
    9.732983e-07, 9.733005e-07, 9.73292e-07, 9.732944e-07, 9.732875e-07, 
    9.732893e-07, 9.732876e-07, 9.732881e-07, 9.732876e-07, 9.732902e-07, 
    9.73289e-07, 9.732913e-07, 9.733001e-07, 9.732975e-07, 9.733052e-07, 
    9.733099e-07, 9.733129e-07, 9.733151e-07, 9.733149e-07, 9.733142e-07, 
    9.733112e-07, 9.733084e-07, 9.733062e-07, 9.733047e-07, 9.733033e-07, 
    9.732989e-07, 9.732967e-07, 9.732915e-07, 9.732925e-07, 9.732909e-07, 
    9.732894e-07, 9.732869e-07, 9.732873e-07, 9.732862e-07, 9.73291e-07, 
    9.732878e-07, 9.73293e-07, 9.732915e-07, 9.733029e-07, 9.733072e-07, 
    9.733091e-07, 9.733106e-07, 9.733145e-07, 9.733119e-07, 9.733129e-07, 
    9.733104e-07, 9.733088e-07, 9.733096e-07, 9.733046e-07, 9.733066e-07, 
    9.732966e-07, 9.733009e-07, 9.732896e-07, 9.732922e-07, 9.732889e-07, 
    9.732906e-07, 9.732877e-07, 9.732904e-07, 9.732859e-07, 9.732848e-07, 
    9.732855e-07, 9.732829e-07, 9.732905e-07, 9.732876e-07, 9.733096e-07, 
    9.733095e-07, 9.733088e-07, 9.733116e-07, 9.733117e-07, 9.733142e-07, 
    9.73312e-07, 9.73311e-07, 9.733087e-07, 9.733074e-07, 9.73306e-07, 
    9.733031e-07, 9.732998e-07, 9.732953e-07, 9.732921e-07, 9.7329e-07, 
    9.732913e-07, 9.732901e-07, 9.732914e-07, 9.73292e-07, 9.732852e-07, 
    9.73289e-07, 9.732832e-07, 9.732836e-07, 9.732862e-07, 9.732836e-07, 
    9.733094e-07, 9.733101e-07, 9.733127e-07, 9.733106e-07, 9.733144e-07, 
    9.733124e-07, 9.733111e-07, 9.733066e-07, 9.733055e-07, 9.733046e-07, 
    9.733028e-07, 9.733004e-07, 9.732962e-07, 9.732926e-07, 9.732893e-07, 
    9.732896e-07, 9.732895e-07, 9.732887e-07, 9.732905e-07, 9.732885e-07, 
    9.732881e-07, 9.73289e-07, 9.732836e-07, 9.732852e-07, 9.732836e-07, 
    9.732846e-07, 9.733099e-07, 9.733086e-07, 9.733093e-07, 9.73308e-07, 
    9.733089e-07, 9.73305e-07, 9.733037e-07, 9.732981e-07, 9.733004e-07, 
    9.732968e-07, 9.733001e-07, 9.732995e-07, 9.732967e-07, 9.732998e-07, 
    9.732928e-07, 9.732976e-07, 9.732887e-07, 9.732935e-07, 9.732885e-07, 
    9.732894e-07, 9.732878e-07, 9.732864e-07, 9.732847e-07, 9.732815e-07, 
    9.732823e-07, 9.732796e-07, 9.733068e-07, 9.733051e-07, 9.733053e-07, 
    9.733036e-07, 9.733023e-07, 9.732996e-07, 9.732952e-07, 9.732969e-07, 
    9.732938e-07, 9.732933e-07, 9.732978e-07, 9.73295e-07, 9.733041e-07, 
    9.733026e-07, 9.733035e-07, 9.733067e-07, 9.732964e-07, 9.733017e-07, 
    9.73292e-07, 9.732948e-07, 9.732867e-07, 9.732908e-07, 9.732827e-07, 
    9.732793e-07, 9.732761e-07, 9.732723e-07, 9.733043e-07, 9.733053e-07, 
    9.733034e-07, 9.733006e-07, 9.73298e-07, 9.732947e-07, 9.732944e-07, 
    9.732937e-07, 9.732921e-07, 9.732908e-07, 9.732935e-07, 9.732904e-07, 
    9.733022e-07, 9.73296e-07, 9.733058e-07, 9.733028e-07, 9.733008e-07, 
    9.733017e-07, 9.73297e-07, 9.73296e-07, 9.732915e-07, 9.732938e-07, 
    9.732802e-07, 9.732862e-07, 9.732694e-07, 9.732742e-07, 9.733058e-07, 
    9.733043e-07, 9.732991e-07, 9.733016e-07, 9.732945e-07, 9.732928e-07, 
    9.732913e-07, 9.732895e-07, 9.732894e-07, 9.732883e-07, 9.732901e-07, 
    9.732884e-07, 9.732947e-07, 9.732919e-07, 9.732996e-07, 9.732978e-07, 
    9.732986e-07, 9.732996e-07, 9.732967e-07, 9.732935e-07, 9.732934e-07, 
    9.732925e-07, 9.732896e-07, 9.732945e-07, 9.732794e-07, 9.732887e-07, 
    9.733026e-07, 9.732997e-07, 9.732994e-07, 9.733004e-07, 9.732929e-07, 
    9.732956e-07, 9.732883e-07, 9.732903e-07, 9.73287e-07, 9.732887e-07, 
    9.732889e-07, 9.73291e-07, 9.732922e-07, 9.732955e-07, 9.732981e-07, 
    9.733003e-07, 9.732998e-07, 9.732975e-07, 9.732933e-07, 9.732893e-07, 
    9.732902e-07, 9.732873e-07, 9.73295e-07, 9.732918e-07, 9.73293e-07, 
    9.732897e-07, 9.732969e-07, 9.732909e-07, 9.732985e-07, 9.732978e-07, 
    9.732958e-07, 9.732915e-07, 9.732906e-07, 9.732896e-07, 9.732903e-07, 
    9.732931e-07, 9.732937e-07, 9.732958e-07, 9.732963e-07, 9.732979e-07, 
    9.732993e-07, 9.73298e-07, 9.732968e-07, 9.732931e-07, 9.7329e-07, 
    9.732864e-07, 9.732855e-07, 9.732814e-07, 9.732848e-07, 9.732793e-07, 
    9.73284e-07, 9.732759e-07, 9.732904e-07, 9.732842e-07, 9.732956e-07, 
    9.732944e-07, 9.732921e-07, 9.73287e-07, 9.732897e-07, 9.732865e-07, 
    9.732937e-07, 9.732975e-07, 9.732984e-07, 9.733002e-07, 9.732984e-07, 
    9.732985e-07, 9.732967e-07, 9.732972e-07, 9.73293e-07, 9.732953e-07, 
    9.732889e-07, 9.732865e-07, 9.7328e-07, 9.732759e-07, 9.732718e-07, 
    9.732699e-07, 9.732694e-07, 9.732692e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  -3.823413e-25, 2.107779e-25, 3.38225e-25, -7.548789e-25, 3.38225e-25, 
    -8.284061e-25, 1.56858e-25, -1.56858e-25, 1.617598e-25, 2.058761e-25, 
    -2.843051e-25, -6.078246e-25, 2.843051e-25, 1.230355e-24, -7.842898e-26, 
    -6.372354e-26, 9.019333e-25, -2.843051e-25, -2.254833e-25, -1.81367e-25, 
    5.490028e-25, -7.156644e-25, 5.686101e-25, -2.254833e-25, 3.235195e-25, 
    2.107779e-25, 1.323489e-25, -3.725376e-25, -3.529304e-25, -1.470543e-25, 
    1.078398e-25, -3.137159e-25, 3.578322e-25, 7.450753e-25, -4.852793e-25, 
    -3.431268e-26, 2.205815e-25, -5.882173e-26, -7.548789e-25, 3.921449e-26, 
    5.784137e-25, 3.088141e-25, -1.862688e-25, 8.529151e-25, 6.813517e-25, 
    -1.078398e-25, -2.745014e-25, 9.313441e-26, -6.372354e-25, 4.117521e-25, 
    -1.274471e-25, -4.705739e-25, 8.333079e-25, -9.803622e-26, -6.47039e-25, 
    -1.117613e-24, 8.235043e-25, 7.989952e-25, 1.56858e-25, -5.98021e-25, 
    6.862535e-26, 4.607703e-25, -3.62734e-25, -1.960724e-25, 5.391992e-25, 
    3.061136e-41, -1.225453e-25, 6.960572e-25, 5.833155e-25, -1.078398e-25, 
    -6.666463e-25, -2.156797e-25, -7.352717e-25, -1.063693e-24, 
    -1.019577e-24, -1.470543e-25, 1.132318e-24, -6.862535e-25, 6.862535e-26, 
    7.695843e-25, -1.176435e-25, 2.254833e-25, 4.019485e-25, -4.509666e-25, 
    2.401887e-25, -7.842898e-26, 2.205815e-25, -1.019577e-24, 2.843051e-25, 
    -2.941087e-26, -1.186238e-24, -6.274318e-25, 4.607703e-25, 5.391992e-25, 
    -7.25468e-25, -1.666616e-25, 2.843051e-25, -1.372507e-25, 1.960724e-26, 
    -6.078246e-25, -4.705739e-25, 2.254833e-25, -4.852793e-25, 1.019577e-24, 
    -5.293956e-25, -5.293956e-25, 6.715481e-25, -2.156797e-25, 1.421525e-25, 
    2.745014e-25, 8.333079e-26, -6.666463e-25, 5.539047e-25, 2.107779e-25, 
    8.82326e-25, 7.646825e-25, 2.892069e-25, -2.794032e-25, -5.490028e-25, 
    6.274318e-25, -4.068503e-25, 1.078398e-25, 5.19592e-25, -2.450906e-25, 
    -5.686101e-25, -3.872431e-25, -1.274471e-25, -7.450753e-25, 7.744861e-25, 
    6.029227e-25, 0, 3.333231e-25, -4.901811e-27, 1.960724e-26, 1.960724e-25, 
    4.852793e-25, 5.244938e-25, -1.764652e-25, 5.048866e-25, 1.56858e-25, 
    -4.264576e-25, -3.921449e-26, -2.548942e-25, 5.490028e-25, 4.607703e-25, 
    1.274471e-25, -1.470543e-25, 9.411477e-25, 3.62734e-25, 3.823413e-25, 
    -8.186024e-25, -1.960724e-25, 2.254833e-25, 1.470543e-25, -3.235195e-25, 
    3.62734e-25, -1.960724e-26, -1.519561e-25, -5.588064e-25, 1.274471e-25, 
    1.56858e-25, 7.352717e-25, 3.529304e-25, -1.372507e-25, -1.401918e-24, 
    7.450753e-25, -6.372354e-25, 8.431115e-25, 5.98021e-25, 2.745014e-25, 
    -2.548942e-25, 8.82326e-26, -5.048866e-25, -4.41163e-25, 5.588064e-25, 
    -3.431268e-25, 1.960724e-25, -4.215557e-25, -1.470543e-25, -2.843051e-25, 
    -2.499924e-25, 1.475445e-24, -9.803622e-27, -3.039123e-25, -1.470543e-26, 
    3.970467e-25, -4.41163e-25, 3.921449e-26, -1.274471e-25, 5.588064e-25, 
    2.59796e-25, -4.460648e-25, -6.862535e-26, 3.921449e-26, 1.960724e-25, 
    2.401887e-25, 6.666463e-25, -1.56858e-25, -6.862535e-26, -1.81367e-25, 
    3.235195e-25, 8.82326e-26, -4.901811e-25, -2.941087e-25, -1.960724e-25, 
    2.941087e-25, 1.960724e-26, -4.019485e-25, 8.03897e-25, -6.274318e-25, 
    6.666463e-25, -1.166631e-24, -6.122413e-41, -1.176435e-25, 9.705585e-25, 
    -3.431268e-25, 4.999847e-25, -4.901811e-26, 2.303851e-25, 1.56858e-25, 
    -1.078398e-25, 4.901811e-27, 4.313593e-25, -2.058761e-25, -9.803622e-27, 
    -1.048988e-24, 2.352869e-25, 5.588064e-25, 9.999695e-25, -1.960724e-25, 
    4.950829e-25, 1.470543e-25, -7.156644e-25, 1.127417e-25, -1.960724e-26, 
    4.509666e-25, 5.539047e-25, 1.862688e-25, 6.960572e-25, 4.41163e-25, 
    4.509666e-25, -1.470543e-25, 4.509666e-25, 3.480286e-25, -1.862688e-25, 
    4.460648e-25, 4.754757e-25, 1.02938e-25, -1.470543e-26, 7.744861e-25, 
    -8.82326e-26, 3.921449e-26, -3.039123e-25, -6.862535e-26, -9.803622e-26, 
    2.450906e-25, 2.450906e-25, 1.372507e-25, 1.078398e-25, 8.82326e-26, 
    6.862535e-25, 5.19592e-25, 2.843051e-25, 6.960572e-25, 2.745014e-25, 
    -2.058761e-25, 1.117613e-24, 2.401887e-25, 7.25468e-25, -3.235195e-25, 
    -1.274471e-25, 1.176435e-25, 6.715481e-25, 5.784137e-25, -3.774394e-25, 
    8.284061e-25, 8.431115e-25, -2.745014e-25, 3.431268e-25, 1.470543e-25, 
    2.843051e-25, -2.59796e-25, -3.088141e-25, -9.803622e-26, 1.470543e-25, 
    2.941087e-26, 2.548942e-25, -2.646978e-25, -7.940934e-25, -5.391992e-26, 
    -1.372507e-25, 9.901658e-25, 3.62734e-25, 3.039123e-25, 2.843051e-25, 
    -5.490028e-25, -7.842898e-26, -4.607703e-25, 5.882173e-26, -9.803622e-27, 
    -2.254833e-25, -4.41163e-26, 1.372507e-25, -6.372354e-25, 9.803622e-26, 
    9.705585e-25, 2.254833e-25, -9.803622e-26, 2.303851e-25, 8.333079e-25, 
    -6.862535e-25, -7.842898e-26, -2.352869e-25, -8.82326e-26, -2.303851e-25, 
    3.186177e-25, -4.509666e-25, 9.068351e-25, 9.019333e-25, 8.921296e-25, 
    1.294078e-24, 1.421525e-25, 2.843051e-25, 7.25468e-25, -5.686101e-25, 
    3.725376e-25, -6.372354e-26, 7.058608e-25, -4.558684e-25, -6.862535e-25, 
    3.235195e-25, -5.097883e-25, -2.303851e-25, 2.941087e-26, -3.578322e-25, 
    -3.62734e-25, -2.450906e-25, 3.333231e-25,
  9.436979e-32, 9.436942e-32, 9.436949e-32, 9.436918e-32, 9.436935e-32, 
    9.436915e-32, 9.436972e-32, 9.43694e-32, 9.43696e-32, 9.436976e-32, 
    9.436859e-32, 9.436917e-32, 9.436799e-32, 9.436836e-32, 9.436744e-32, 
    9.436805e-32, 9.436732e-32, 9.436746e-32, 9.436703e-32, 9.436715e-32, 
    9.436661e-32, 9.436698e-32, 9.436633e-32, 9.43667e-32, 9.436664e-32, 
    9.436699e-32, 9.436905e-32, 9.436866e-32, 9.436907e-32, 9.436902e-32, 
    9.436905e-32, 9.436935e-32, 9.43695e-32, 9.436982e-32, 9.436976e-32, 
    9.436953e-32, 9.4369e-32, 9.436917e-32, 9.436872e-32, 9.436873e-32, 
    9.436823e-32, 9.436845e-32, 9.436761e-32, 9.436785e-32, 9.436715e-32, 
    9.436732e-32, 9.436716e-32, 9.436721e-32, 9.436715e-32, 9.436741e-32, 
    9.43673e-32, 9.436753e-32, 9.436841e-32, 9.436815e-32, 9.436893e-32, 
    9.436939e-32, 9.43697e-32, 9.436992e-32, 9.436989e-32, 9.436983e-32, 
    9.436953e-32, 9.436924e-32, 9.436902e-32, 9.436887e-32, 9.436873e-32, 
    9.43683e-32, 9.436807e-32, 9.436755e-32, 9.436765e-32, 9.436749e-32, 
    9.436734e-32, 9.436709e-32, 9.436713e-32, 9.436702e-32, 9.436749e-32, 
    9.436718e-32, 9.43677e-32, 9.436756e-32, 9.436869e-32, 9.436913e-32, 
    9.436931e-32, 9.436947e-32, 9.436987e-32, 9.43696e-32, 9.43697e-32, 
    9.436944e-32, 9.436929e-32, 9.436937e-32, 9.436887e-32, 9.436906e-32, 
    9.436806e-32, 9.436849e-32, 9.436736e-32, 9.436763e-32, 9.436729e-32, 
    9.436746e-32, 9.436717e-32, 9.436743e-32, 9.436698e-32, 9.436688e-32, 
    9.436695e-32, 9.436669e-32, 9.436745e-32, 9.436716e-32, 9.436937e-32, 
    9.436936e-32, 9.436929e-32, 9.436956e-32, 9.436958e-32, 9.436982e-32, 
    9.43696e-32, 9.436951e-32, 9.436927e-32, 9.436914e-32, 9.4369e-32, 
    9.436872e-32, 9.436839e-32, 9.436793e-32, 9.436761e-32, 9.436739e-32, 
    9.436753e-32, 9.436741e-32, 9.436754e-32, 9.436761e-32, 9.436692e-32, 
    9.43673e-32, 9.436672e-32, 9.436675e-32, 9.436702e-32, 9.436675e-32, 
    9.436934e-32, 9.436942e-32, 9.436968e-32, 9.436948e-32, 9.436985e-32, 
    9.436964e-32, 9.436952e-32, 9.436906e-32, 9.436896e-32, 9.436886e-32, 
    9.436868e-32, 9.436844e-32, 9.436802e-32, 9.436766e-32, 9.436733e-32, 
    9.436736e-32, 9.436735e-32, 9.436728e-32, 9.436746e-32, 9.436724e-32, 
    9.436721e-32, 9.43673e-32, 9.436676e-32, 9.436691e-32, 9.436675e-32, 
    9.436686e-32, 9.43694e-32, 9.436927e-32, 9.436934e-32, 9.436921e-32, 
    9.43693e-32, 9.43689e-32, 9.436878e-32, 9.436822e-32, 9.436845e-32, 
    9.436808e-32, 9.436841e-32, 9.436835e-32, 9.436807e-32, 9.436839e-32, 
    9.436768e-32, 9.436816e-32, 9.436727e-32, 9.436775e-32, 9.436724e-32, 
    9.436733e-32, 9.436718e-32, 9.436704e-32, 9.436687e-32, 9.436655e-32, 
    9.436662e-32, 9.436636e-32, 9.436908e-32, 9.436892e-32, 9.436893e-32, 
    9.436876e-32, 9.436863e-32, 9.436836e-32, 9.436792e-32, 9.436809e-32, 
    9.436778e-32, 9.436772e-32, 9.436818e-32, 9.43679e-32, 9.436881e-32, 
    9.436866e-32, 9.436875e-32, 9.436907e-32, 9.436805e-32, 9.436857e-32, 
    9.436761e-32, 9.436789e-32, 9.436706e-32, 9.436748e-32, 9.436666e-32, 
    9.436632e-32, 9.4366e-32, 9.436562e-32, 9.436883e-32, 9.436894e-32, 
    9.436874e-32, 9.436846e-32, 9.436821e-32, 9.436787e-32, 9.436783e-32, 
    9.436778e-32, 9.436761e-32, 9.436747e-32, 9.436775e-32, 9.436743e-32, 
    9.436863e-32, 9.4368e-32, 9.436898e-32, 9.436869e-32, 9.436848e-32, 
    9.436857e-32, 9.43681e-32, 9.436799e-32, 9.436755e-32, 9.436778e-32, 
    9.436641e-32, 9.436701e-32, 9.436533e-32, 9.43658e-32, 9.436898e-32, 
    9.436883e-32, 9.436831e-32, 9.436856e-32, 9.436785e-32, 9.436768e-32, 
    9.436753e-32, 9.436735e-32, 9.436733e-32, 9.436723e-32, 9.43674e-32, 
    9.436723e-32, 9.436787e-32, 9.436759e-32, 9.436837e-32, 9.436818e-32, 
    9.436826e-32, 9.436836e-32, 9.436806e-32, 9.436775e-32, 9.436774e-32, 
    9.436764e-32, 9.436736e-32, 9.436785e-32, 9.436633e-32, 9.436726e-32, 
    9.436867e-32, 9.436838e-32, 9.436834e-32, 9.436845e-32, 9.436769e-32, 
    9.436796e-32, 9.436723e-32, 9.436743e-32, 9.43671e-32, 9.436726e-32, 
    9.436729e-32, 9.436749e-32, 9.436763e-32, 9.436795e-32, 9.436822e-32, 
    9.436843e-32, 9.436838e-32, 9.436815e-32, 9.436773e-32, 9.436733e-32, 
    9.436742e-32, 9.436713e-32, 9.43679e-32, 9.436758e-32, 9.43677e-32, 
    9.436738e-32, 9.436809e-32, 9.436748e-32, 9.436825e-32, 9.436818e-32, 
    9.436797e-32, 9.436755e-32, 9.436746e-32, 9.436736e-32, 9.436742e-32, 
    9.436772e-32, 9.436777e-32, 9.436798e-32, 9.436803e-32, 9.436819e-32, 
    9.436833e-32, 9.43682e-32, 9.436808e-32, 9.436772e-32, 9.436739e-32, 
    9.436704e-32, 9.436695e-32, 9.436654e-32, 9.436688e-32, 9.436632e-32, 
    9.436679e-32, 9.436598e-32, 9.436745e-32, 9.436681e-32, 9.436796e-32, 
    9.436784e-32, 9.436761e-32, 9.43671e-32, 9.436738e-32, 9.436705e-32, 
    9.436777e-32, 9.436814e-32, 9.436824e-32, 9.436842e-32, 9.436823e-32, 
    9.436825e-32, 9.436808e-32, 9.436813e-32, 9.43677e-32, 9.436793e-32, 
    9.436729e-32, 9.436705e-32, 9.436639e-32, 9.436598e-32, 9.436557e-32, 
    9.436538e-32, 9.436533e-32, 9.436531e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.499488e-14, 4.511822e-14, 4.509426e-14, 4.519366e-14, 4.513855e-14, 
    4.520361e-14, 4.501992e-14, 4.51231e-14, 4.505725e-14, 4.500602e-14, 
    4.538633e-14, 4.51981e-14, 4.55818e-14, 4.54619e-14, 4.576297e-14, 
    4.556313e-14, 4.580325e-14, 4.575726e-14, 4.589574e-14, 4.585608e-14, 
    4.603296e-14, 4.591404e-14, 4.612464e-14, 4.600459e-14, 4.602336e-14, 
    4.59101e-14, 4.523604e-14, 4.536289e-14, 4.522851e-14, 4.524661e-14, 
    4.52385e-14, 4.513967e-14, 4.508981e-14, 4.498549e-14, 4.500444e-14, 
    4.508108e-14, 4.525475e-14, 4.519585e-14, 4.534434e-14, 4.534099e-14, 
    4.550612e-14, 4.543169e-14, 4.570899e-14, 4.563024e-14, 4.585774e-14, 
    4.580055e-14, 4.585504e-14, 4.583853e-14, 4.585526e-14, 4.577138e-14, 
    4.580732e-14, 4.573351e-14, 4.544562e-14, 4.553027e-14, 4.527764e-14, 
    4.512547e-14, 4.502444e-14, 4.495267e-14, 4.496282e-14, 4.498215e-14, 
    4.508153e-14, 4.517494e-14, 4.524609e-14, 4.529365e-14, 4.534051e-14, 
    4.548214e-14, 4.555715e-14, 4.572489e-14, 4.569467e-14, 4.574589e-14, 
    4.579486e-14, 4.587699e-14, 4.586348e-14, 4.589964e-14, 4.574457e-14, 
    4.584764e-14, 4.567745e-14, 4.572401e-14, 4.53531e-14, 4.521175e-14, 
    4.51515e-14, 4.509886e-14, 4.497062e-14, 4.505918e-14, 4.502427e-14, 
    4.510735e-14, 4.516009e-14, 4.513402e-14, 4.529495e-14, 4.52324e-14, 
    4.556159e-14, 4.541989e-14, 4.578915e-14, 4.570088e-14, 4.581031e-14, 
    4.575449e-14, 4.585011e-14, 4.576406e-14, 4.591311e-14, 4.594553e-14, 
    4.592338e-14, 4.600852e-14, 4.575928e-14, 4.585503e-14, 4.513328e-14, 
    4.513753e-14, 4.515736e-14, 4.507018e-14, 4.506485e-14, 4.498496e-14, 
    4.505606e-14, 4.508632e-14, 4.516316e-14, 4.520857e-14, 4.525173e-14, 
    4.534659e-14, 4.545245e-14, 4.560038e-14, 4.57066e-14, 4.577775e-14, 
    4.573414e-14, 4.577264e-14, 4.572959e-14, 4.570941e-14, 4.593338e-14, 
    4.580765e-14, 4.599628e-14, 4.598585e-14, 4.59005e-14, 4.598702e-14, 
    4.514052e-14, 4.511604e-14, 4.503098e-14, 4.509755e-14, 4.497626e-14, 
    4.504414e-14, 4.508315e-14, 4.523367e-14, 4.526676e-14, 4.529739e-14, 
    4.53579e-14, 4.54355e-14, 4.557152e-14, 4.56898e-14, 4.579772e-14, 
    4.578982e-14, 4.57926e-14, 4.581668e-14, 4.5757e-14, 4.582647e-14, 
    4.583812e-14, 4.580765e-14, 4.598445e-14, 4.593397e-14, 4.598563e-14, 
    4.595276e-14, 4.5124e-14, 4.516519e-14, 4.514293e-14, 4.518478e-14, 
    4.515529e-14, 4.528634e-14, 4.532561e-14, 4.550927e-14, 4.543396e-14, 
    4.555385e-14, 4.544616e-14, 4.546524e-14, 4.555769e-14, 4.545199e-14, 
    4.568325e-14, 4.552645e-14, 4.581761e-14, 4.56611e-14, 4.582741e-14, 
    4.579725e-14, 4.58472e-14, 4.589191e-14, 4.594816e-14, 4.605184e-14, 
    4.602784e-14, 4.611453e-14, 4.522659e-14, 4.527997e-14, 4.52753e-14, 
    4.533116e-14, 4.537245e-14, 4.546195e-14, 4.560536e-14, 4.555145e-14, 
    4.565042e-14, 4.567028e-14, 4.551993e-14, 4.561223e-14, 4.53157e-14, 
    4.536362e-14, 4.533511e-14, 4.523079e-14, 4.556384e-14, 4.539299e-14, 
    4.570835e-14, 4.561592e-14, 4.588553e-14, 4.575148e-14, 4.601462e-14, 
    4.612689e-14, 4.62326e-14, 4.635587e-14, 4.530912e-14, 4.527286e-14, 
    4.533781e-14, 4.542757e-14, 4.551089e-14, 4.562155e-14, 4.563288e-14, 
    4.565359e-14, 4.570726e-14, 4.575236e-14, 4.566011e-14, 4.576366e-14, 
    4.537467e-14, 4.557867e-14, 4.525912e-14, 4.535538e-14, 4.542229e-14, 
    4.539297e-14, 4.55453e-14, 4.558117e-14, 4.572683e-14, 4.565157e-14, 
    4.609917e-14, 4.590131e-14, 4.644975e-14, 4.629669e-14, 4.526018e-14, 
    4.530901e-14, 4.547879e-14, 4.539804e-14, 4.562895e-14, 4.568572e-14, 
    4.573188e-14, 4.579081e-14, 4.57972e-14, 4.583211e-14, 4.577489e-14, 
    4.582986e-14, 4.562178e-14, 4.571481e-14, 4.545943e-14, 4.552161e-14, 
    4.549302e-14, 4.546163e-14, 4.555849e-14, 4.566156e-14, 4.566381e-14, 
    4.569683e-14, 4.578978e-14, 4.562989e-14, 4.61246e-14, 4.58192e-14, 
    4.536224e-14, 4.545616e-14, 4.546962e-14, 4.543324e-14, 4.568003e-14, 
    4.559065e-14, 4.583127e-14, 4.576628e-14, 4.587275e-14, 4.581985e-14, 
    4.581206e-14, 4.57441e-14, 4.570176e-14, 4.559474e-14, 4.550762e-14, 
    4.543852e-14, 4.545459e-14, 4.553049e-14, 4.566787e-14, 4.579775e-14, 
    4.576931e-14, 4.586466e-14, 4.561222e-14, 4.57181e-14, 4.567717e-14, 
    4.578388e-14, 4.555001e-14, 4.574905e-14, 4.549908e-14, 4.552102e-14, 
    4.558887e-14, 4.572525e-14, 4.575547e-14, 4.578765e-14, 4.576781e-14, 
    4.567137e-14, 4.565558e-14, 4.558724e-14, 4.556834e-14, 4.551625e-14, 
    4.547309e-14, 4.551251e-14, 4.555389e-14, 4.567143e-14, 4.577724e-14, 
    4.589254e-14, 4.592076e-14, 4.60552e-14, 4.59457e-14, 4.612628e-14, 
    4.597268e-14, 4.623852e-14, 4.576064e-14, 4.596825e-14, 4.559198e-14, 
    4.563257e-14, 4.570592e-14, 4.58741e-14, 4.578338e-14, 4.58895e-14, 
    4.565497e-14, 4.553308e-14, 4.550159e-14, 4.544271e-14, 4.550293e-14, 
    4.549804e-14, 4.555564e-14, 4.553713e-14, 4.567533e-14, 4.560111e-14, 
    4.581185e-14, 4.588867e-14, 4.610543e-14, 4.623811e-14, 4.637311e-14, 
    4.643264e-14, 4.645076e-14, 4.645833e-14 ;

 LITR1N_vr =
  5.557722e-05, 5.557701e-05, 5.557705e-05, 5.557688e-05, 5.557698e-05, 
    5.557686e-05, 5.557718e-05, 5.5577e-05, 5.557711e-05, 5.557721e-05, 
    5.557654e-05, 5.557687e-05, 5.55762e-05, 5.557641e-05, 5.557589e-05, 
    5.557623e-05, 5.557582e-05, 5.55759e-05, 5.557566e-05, 5.557573e-05, 
    5.557542e-05, 5.557562e-05, 5.557526e-05, 5.557547e-05, 5.557543e-05, 
    5.557563e-05, 5.557681e-05, 5.557658e-05, 5.557682e-05, 5.557679e-05, 
    5.55768e-05, 5.557697e-05, 5.557706e-05, 5.557724e-05, 5.557721e-05, 
    5.557707e-05, 5.557677e-05, 5.557687e-05, 5.557662e-05, 5.557662e-05, 
    5.557634e-05, 5.557646e-05, 5.557598e-05, 5.557612e-05, 5.557572e-05, 
    5.557582e-05, 5.557573e-05, 5.557575e-05, 5.557573e-05, 5.557587e-05, 
    5.557581e-05, 5.557594e-05, 5.557644e-05, 5.557629e-05, 5.557673e-05, 
    5.5577e-05, 5.557717e-05, 5.55773e-05, 5.557728e-05, 5.557725e-05, 
    5.557707e-05, 5.557691e-05, 5.557679e-05, 5.55767e-05, 5.557662e-05, 
    5.557638e-05, 5.557625e-05, 5.557595e-05, 5.557601e-05, 5.557592e-05, 
    5.557583e-05, 5.557569e-05, 5.557571e-05, 5.557565e-05, 5.557592e-05, 
    5.557574e-05, 5.557603e-05, 5.557595e-05, 5.55766e-05, 5.557685e-05, 
    5.557695e-05, 5.557705e-05, 5.557727e-05, 5.557711e-05, 5.557717e-05, 
    5.557703e-05, 5.557694e-05, 5.557698e-05, 5.55767e-05, 5.557681e-05, 
    5.557624e-05, 5.557649e-05, 5.557584e-05, 5.557599e-05, 5.557581e-05, 
    5.55759e-05, 5.557574e-05, 5.557589e-05, 5.557563e-05, 5.557557e-05, 
    5.557561e-05, 5.557546e-05, 5.557589e-05, 5.557573e-05, 5.557698e-05, 
    5.557698e-05, 5.557694e-05, 5.557709e-05, 5.55771e-05, 5.557724e-05, 
    5.557712e-05, 5.557707e-05, 5.557693e-05, 5.557685e-05, 5.557678e-05, 
    5.557661e-05, 5.557643e-05, 5.557617e-05, 5.557599e-05, 5.557586e-05, 
    5.557594e-05, 5.557587e-05, 5.557595e-05, 5.557598e-05, 5.557559e-05, 
    5.557581e-05, 5.557548e-05, 5.55755e-05, 5.557565e-05, 5.55755e-05, 
    5.557697e-05, 5.557701e-05, 5.557716e-05, 5.557705e-05, 5.557726e-05, 
    5.557714e-05, 5.557707e-05, 5.557681e-05, 5.557675e-05, 5.55767e-05, 
    5.557659e-05, 5.557646e-05, 5.557622e-05, 5.557602e-05, 5.557583e-05, 
    5.557584e-05, 5.557583e-05, 5.557579e-05, 5.55759e-05, 5.557578e-05, 
    5.557576e-05, 5.557581e-05, 5.55755e-05, 5.557559e-05, 5.55755e-05, 
    5.557556e-05, 5.5577e-05, 5.557693e-05, 5.557697e-05, 5.557689e-05, 
    5.557694e-05, 5.557672e-05, 5.557665e-05, 5.557633e-05, 5.557646e-05, 
    5.557625e-05, 5.557644e-05, 5.557641e-05, 5.557625e-05, 5.557643e-05, 
    5.557603e-05, 5.55763e-05, 5.557579e-05, 5.557606e-05, 5.557578e-05, 
    5.557583e-05, 5.557574e-05, 5.557566e-05, 5.557557e-05, 5.557538e-05, 
    5.557543e-05, 5.557527e-05, 5.557682e-05, 5.557673e-05, 5.557674e-05, 
    5.557664e-05, 5.557657e-05, 5.557641e-05, 5.557616e-05, 5.557626e-05, 
    5.557608e-05, 5.557605e-05, 5.557631e-05, 5.557615e-05, 5.557667e-05, 
    5.557658e-05, 5.557663e-05, 5.557681e-05, 5.557623e-05, 5.557653e-05, 
    5.557598e-05, 5.557614e-05, 5.557567e-05, 5.557591e-05, 5.557545e-05, 
    5.557525e-05, 5.557507e-05, 5.557486e-05, 5.557668e-05, 5.557674e-05, 
    5.557663e-05, 5.557647e-05, 5.557633e-05, 5.557613e-05, 5.557611e-05, 
    5.557608e-05, 5.557598e-05, 5.557591e-05, 5.557607e-05, 5.557589e-05, 
    5.557656e-05, 5.557621e-05, 5.557677e-05, 5.55766e-05, 5.557648e-05, 
    5.557653e-05, 5.557627e-05, 5.557621e-05, 5.557595e-05, 5.557608e-05, 
    5.55753e-05, 5.557565e-05, 5.557469e-05, 5.557496e-05, 5.557676e-05, 
    5.557668e-05, 5.557638e-05, 5.557652e-05, 5.557612e-05, 5.557602e-05, 
    5.557594e-05, 5.557584e-05, 5.557583e-05, 5.557577e-05, 5.557587e-05, 
    5.557577e-05, 5.557613e-05, 5.557597e-05, 5.557642e-05, 5.557631e-05, 
    5.557636e-05, 5.557641e-05, 5.557624e-05, 5.557606e-05, 5.557606e-05, 
    5.5576e-05, 5.557584e-05, 5.557612e-05, 5.557526e-05, 5.557579e-05, 
    5.557658e-05, 5.557642e-05, 5.55764e-05, 5.557646e-05, 5.557603e-05, 
    5.557619e-05, 5.557577e-05, 5.557588e-05, 5.55757e-05, 5.557579e-05, 
    5.55758e-05, 5.557592e-05, 5.557599e-05, 5.557618e-05, 5.557633e-05, 
    5.557645e-05, 5.557642e-05, 5.557629e-05, 5.557605e-05, 5.557583e-05, 
    5.557588e-05, 5.557571e-05, 5.557615e-05, 5.557597e-05, 5.557604e-05, 
    5.557585e-05, 5.557626e-05, 5.557591e-05, 5.557635e-05, 5.557631e-05, 
    5.557619e-05, 5.557595e-05, 5.55759e-05, 5.557585e-05, 5.557588e-05, 
    5.557605e-05, 5.557607e-05, 5.557619e-05, 5.557623e-05, 5.557632e-05, 
    5.557639e-05, 5.557632e-05, 5.557625e-05, 5.557605e-05, 5.557586e-05, 
    5.557566e-05, 5.557561e-05, 5.557538e-05, 5.557557e-05, 5.557526e-05, 
    5.557552e-05, 5.557506e-05, 5.557589e-05, 5.557553e-05, 5.557618e-05, 
    5.557611e-05, 5.557599e-05, 5.557569e-05, 5.557585e-05, 5.557567e-05, 
    5.557607e-05, 5.557629e-05, 5.557634e-05, 5.557645e-05, 5.557634e-05, 
    5.557635e-05, 5.557625e-05, 5.557628e-05, 5.557604e-05, 5.557617e-05, 
    5.55758e-05, 5.557567e-05, 5.557529e-05, 5.557506e-05, 5.557482e-05, 
    5.557472e-05, 5.557469e-05, 5.557467e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.797766e-13, 7.81914e-13, 7.814988e-13, 7.832214e-13, 7.822662e-13, 
    7.833939e-13, 7.802104e-13, 7.819985e-13, 7.808573e-13, 7.799695e-13, 
    7.865604e-13, 7.832983e-13, 7.89948e-13, 7.878701e-13, 7.930878e-13, 
    7.896243e-13, 7.937857e-13, 7.929887e-13, 7.953886e-13, 7.947014e-13, 
    7.977667e-13, 7.957057e-13, 7.993555e-13, 7.972752e-13, 7.976004e-13, 
    7.956376e-13, 7.839559e-13, 7.861543e-13, 7.838254e-13, 7.84139e-13, 
    7.839985e-13, 7.822857e-13, 7.814217e-13, 7.796137e-13, 7.799421e-13, 
    7.812703e-13, 7.842801e-13, 7.832593e-13, 7.858328e-13, 7.857747e-13, 
    7.886364e-13, 7.873465e-13, 7.921523e-13, 7.907875e-13, 7.947301e-13, 
    7.93739e-13, 7.946834e-13, 7.943972e-13, 7.946871e-13, 7.932335e-13, 
    7.938564e-13, 7.925772e-13, 7.87588e-13, 7.89055e-13, 7.846768e-13, 
    7.820397e-13, 7.802887e-13, 7.790449e-13, 7.792208e-13, 7.795558e-13, 
    7.812781e-13, 7.82897e-13, 7.8413e-13, 7.849543e-13, 7.857664e-13, 
    7.882209e-13, 7.895208e-13, 7.924278e-13, 7.919041e-13, 7.927918e-13, 
    7.936404e-13, 7.950637e-13, 7.948296e-13, 7.954563e-13, 7.927688e-13, 
    7.945551e-13, 7.916056e-13, 7.924126e-13, 7.859845e-13, 7.835349e-13, 
    7.824907e-13, 7.815785e-13, 7.793559e-13, 7.808908e-13, 7.802858e-13, 
    7.817255e-13, 7.826396e-13, 7.821877e-13, 7.849768e-13, 7.838927e-13, 
    7.895978e-13, 7.871419e-13, 7.935415e-13, 7.920117e-13, 7.939081e-13, 
    7.929407e-13, 7.945978e-13, 7.931065e-13, 7.956897e-13, 7.962516e-13, 
    7.958676e-13, 7.973432e-13, 7.930237e-13, 7.946832e-13, 7.821749e-13, 
    7.822486e-13, 7.825923e-13, 7.810814e-13, 7.80989e-13, 7.796045e-13, 
    7.808368e-13, 7.813611e-13, 7.826928e-13, 7.834798e-13, 7.842278e-13, 
    7.858718e-13, 7.877062e-13, 7.9027e-13, 7.921108e-13, 7.933439e-13, 
    7.925881e-13, 7.932553e-13, 7.925093e-13, 7.921596e-13, 7.960409e-13, 
    7.93862e-13, 7.97131e-13, 7.969503e-13, 7.954712e-13, 7.969707e-13, 
    7.823004e-13, 7.818762e-13, 7.80402e-13, 7.815558e-13, 7.794538e-13, 
    7.806302e-13, 7.813063e-13, 7.839148e-13, 7.844883e-13, 7.85019e-13, 
    7.860677e-13, 7.874125e-13, 7.897699e-13, 7.918197e-13, 7.936899e-13, 
    7.93553e-13, 7.936012e-13, 7.940185e-13, 7.929843e-13, 7.941883e-13, 
    7.943901e-13, 7.938621e-13, 7.969261e-13, 7.960512e-13, 7.969465e-13, 
    7.963769e-13, 7.820142e-13, 7.82728e-13, 7.823422e-13, 7.830675e-13, 
    7.825564e-13, 7.848275e-13, 7.855081e-13, 7.886911e-13, 7.873859e-13, 
    7.894635e-13, 7.875973e-13, 7.879279e-13, 7.895302e-13, 7.876983e-13, 
    7.917063e-13, 7.889887e-13, 7.940348e-13, 7.913224e-13, 7.942045e-13, 
    7.936819e-13, 7.945475e-13, 7.953222e-13, 7.962971e-13, 7.980939e-13, 
    7.976781e-13, 7.991804e-13, 7.837921e-13, 7.847171e-13, 7.846362e-13, 
    7.856043e-13, 7.863199e-13, 7.87871e-13, 7.903562e-13, 7.894221e-13, 
    7.911372e-13, 7.914812e-13, 7.888757e-13, 7.904753e-13, 7.853364e-13, 
    7.861668e-13, 7.856728e-13, 7.838648e-13, 7.896367e-13, 7.866758e-13, 
    7.921411e-13, 7.905392e-13, 7.952117e-13, 7.928885e-13, 7.97449e-13, 
    7.993946e-13, 8.012265e-13, 8.033629e-13, 7.852224e-13, 7.84594e-13, 
    7.857195e-13, 7.872751e-13, 7.887191e-13, 7.906369e-13, 7.908333e-13, 
    7.911922e-13, 7.921223e-13, 7.929038e-13, 7.913052e-13, 7.930997e-13, 
    7.863584e-13, 7.898938e-13, 7.843559e-13, 7.86024e-13, 7.871837e-13, 
    7.866755e-13, 7.893154e-13, 7.899371e-13, 7.924614e-13, 7.911571e-13, 
    7.989141e-13, 7.954852e-13, 8.049898e-13, 8.023373e-13, 7.843742e-13, 
    7.852205e-13, 7.881629e-13, 7.867634e-13, 7.907651e-13, 7.917489e-13, 
    7.925489e-13, 7.935703e-13, 7.936809e-13, 7.942859e-13, 7.932944e-13, 
    7.942469e-13, 7.906409e-13, 7.922531e-13, 7.878273e-13, 7.889049e-13, 
    7.884094e-13, 7.878654e-13, 7.895439e-13, 7.913302e-13, 7.913692e-13, 
    7.919415e-13, 7.935523e-13, 7.907813e-13, 7.993548e-13, 7.940622e-13, 
    7.861429e-13, 7.877705e-13, 7.880039e-13, 7.873734e-13, 7.916503e-13, 
    7.901013e-13, 7.942713e-13, 7.931451e-13, 7.949903e-13, 7.940735e-13, 
    7.939385e-13, 7.927607e-13, 7.920269e-13, 7.901722e-13, 7.886624e-13, 
    7.874649e-13, 7.877435e-13, 7.890587e-13, 7.914396e-13, 7.936906e-13, 
    7.931975e-13, 7.948501e-13, 7.904751e-13, 7.923101e-13, 7.916008e-13, 
    7.934501e-13, 7.893971e-13, 7.928464e-13, 7.885144e-13, 7.888947e-13, 
    7.900706e-13, 7.92434e-13, 7.929578e-13, 7.935155e-13, 7.931715e-13, 
    7.915002e-13, 7.912266e-13, 7.900422e-13, 7.897146e-13, 7.888119e-13, 
    7.880639e-13, 7.887472e-13, 7.894643e-13, 7.915013e-13, 7.933351e-13, 
    7.953331e-13, 7.958222e-13, 7.981522e-13, 7.962546e-13, 7.993841e-13, 
    7.96722e-13, 8.013292e-13, 7.930474e-13, 7.966452e-13, 7.901243e-13, 
    7.908279e-13, 7.92099e-13, 7.950137e-13, 7.934414e-13, 7.952805e-13, 
    7.91216e-13, 7.891037e-13, 7.885579e-13, 7.875376e-13, 7.885812e-13, 
    7.884964e-13, 7.894946e-13, 7.891739e-13, 7.915689e-13, 7.902827e-13, 
    7.939349e-13, 7.952662e-13, 7.990227e-13, 8.013221e-13, 8.036617e-13, 
    8.046933e-13, 8.050073e-13, 8.051386e-13 ;

 LITR2C =
  1.939613e-05, 1.939611e-05, 1.939611e-05, 1.93961e-05, 1.939611e-05, 
    1.93961e-05, 1.939612e-05, 1.939611e-05, 1.939612e-05, 1.939613e-05, 
    1.939607e-05, 1.93961e-05, 1.939603e-05, 1.939605e-05, 1.9396e-05, 
    1.939604e-05, 1.9396e-05, 1.939601e-05, 1.939598e-05, 1.939599e-05, 
    1.939596e-05, 1.939598e-05, 1.939595e-05, 1.939597e-05, 1.939596e-05, 
    1.939598e-05, 1.939609e-05, 1.939607e-05, 1.939609e-05, 1.939609e-05, 
    1.939609e-05, 1.93961e-05, 1.939611e-05, 1.939613e-05, 1.939613e-05, 
    1.939612e-05, 1.939609e-05, 1.93961e-05, 1.939607e-05, 1.939607e-05, 
    1.939605e-05, 1.939606e-05, 1.939601e-05, 1.939603e-05, 1.939599e-05, 
    1.9396e-05, 1.939599e-05, 1.939599e-05, 1.939599e-05, 1.9396e-05, 
    1.9396e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 1.939608e-05, 
    1.939611e-05, 1.939612e-05, 1.939614e-05, 1.939613e-05, 1.939613e-05, 
    1.939612e-05, 1.93961e-05, 1.939609e-05, 1.939608e-05, 1.939607e-05, 
    1.939605e-05, 1.939604e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 
    1.9396e-05, 1.939599e-05, 1.939599e-05, 1.939598e-05, 1.939601e-05, 
    1.939599e-05, 1.939602e-05, 1.939601e-05, 1.939607e-05, 1.939609e-05, 
    1.93961e-05, 1.939611e-05, 1.939613e-05, 1.939612e-05, 1.939612e-05, 
    1.939611e-05, 1.93961e-05, 1.939611e-05, 1.939608e-05, 1.939609e-05, 
    1.939604e-05, 1.939606e-05, 1.9396e-05, 1.939601e-05, 1.9396e-05, 
    1.939601e-05, 1.939599e-05, 1.9396e-05, 1.939598e-05, 1.939597e-05, 
    1.939598e-05, 1.939597e-05, 1.939601e-05, 1.939599e-05, 1.939611e-05, 
    1.939611e-05, 1.93961e-05, 1.939612e-05, 1.939612e-05, 1.939613e-05, 
    1.939612e-05, 1.939611e-05, 1.93961e-05, 1.939609e-05, 1.939609e-05, 
    1.939607e-05, 1.939605e-05, 1.939603e-05, 1.939601e-05, 1.9396e-05, 
    1.939601e-05, 1.9396e-05, 1.939601e-05, 1.939601e-05, 1.939598e-05, 
    1.9396e-05, 1.939597e-05, 1.939597e-05, 1.939598e-05, 1.939597e-05, 
    1.93961e-05, 1.939611e-05, 1.939612e-05, 1.939611e-05, 1.939613e-05, 
    1.939612e-05, 1.939611e-05, 1.939609e-05, 1.939608e-05, 1.939608e-05, 
    1.939607e-05, 1.939606e-05, 1.939603e-05, 1.939602e-05, 1.9396e-05, 
    1.9396e-05, 1.9396e-05, 1.9396e-05, 1.939601e-05, 1.939599e-05, 
    1.939599e-05, 1.9396e-05, 1.939597e-05, 1.939598e-05, 1.939597e-05, 
    1.939597e-05, 1.939611e-05, 1.93961e-05, 1.93961e-05, 1.93961e-05, 
    1.93961e-05, 1.939608e-05, 1.939608e-05, 1.939605e-05, 1.939606e-05, 
    1.939604e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 
    1.939602e-05, 1.939604e-05, 1.9396e-05, 1.939602e-05, 1.939599e-05, 
    1.9396e-05, 1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 
    1.939596e-05, 1.939595e-05, 1.939609e-05, 1.939608e-05, 1.939608e-05, 
    1.939608e-05, 1.939607e-05, 1.939605e-05, 1.939603e-05, 1.939604e-05, 
    1.939602e-05, 1.939602e-05, 1.939604e-05, 1.939603e-05, 1.939608e-05, 
    1.939607e-05, 1.939607e-05, 1.939609e-05, 1.939604e-05, 1.939606e-05, 
    1.939601e-05, 1.939603e-05, 1.939599e-05, 1.939601e-05, 1.939596e-05, 
    1.939595e-05, 1.939593e-05, 1.939591e-05, 1.939608e-05, 1.939608e-05, 
    1.939607e-05, 1.939606e-05, 1.939605e-05, 1.939603e-05, 1.939603e-05, 
    1.939602e-05, 1.939601e-05, 1.939601e-05, 1.939602e-05, 1.9396e-05, 
    1.939607e-05, 1.939603e-05, 1.939609e-05, 1.939607e-05, 1.939606e-05, 
    1.939606e-05, 1.939604e-05, 1.939603e-05, 1.939601e-05, 1.939602e-05, 
    1.939595e-05, 1.939598e-05, 1.939589e-05, 1.939592e-05, 1.939609e-05, 
    1.939608e-05, 1.939605e-05, 1.939606e-05, 1.939603e-05, 1.939602e-05, 
    1.939601e-05, 1.9396e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939603e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 
    1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939602e-05, 1.939602e-05, 
    1.939601e-05, 1.9396e-05, 1.939603e-05, 1.939595e-05, 1.939599e-05, 
    1.939607e-05, 1.939605e-05, 1.939605e-05, 1.939606e-05, 1.939602e-05, 
    1.939603e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.9396e-05, 1.939601e-05, 1.939601e-05, 1.939603e-05, 1.939605e-05, 
    1.939606e-05, 1.939605e-05, 1.939604e-05, 1.939602e-05, 1.9396e-05, 
    1.9396e-05, 1.939599e-05, 1.939603e-05, 1.939601e-05, 1.939602e-05, 
    1.9396e-05, 1.939604e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 
    1.939603e-05, 1.939601e-05, 1.939601e-05, 1.9396e-05, 1.9396e-05, 
    1.939602e-05, 1.939602e-05, 1.939603e-05, 1.939604e-05, 1.939604e-05, 
    1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939602e-05, 1.9396e-05, 
    1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 1.939595e-05, 
    1.939597e-05, 1.939593e-05, 1.939601e-05, 1.939597e-05, 1.939603e-05, 
    1.939603e-05, 1.939601e-05, 1.939599e-05, 1.9396e-05, 1.939598e-05, 
    1.939602e-05, 1.939604e-05, 1.939605e-05, 1.939606e-05, 1.939605e-05, 
    1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939602e-05, 1.939603e-05, 
    1.9396e-05, 1.939598e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 
    1.93959e-05, 1.939589e-05, 1.939589e-05 ;

 LITR2C_TO_SOIL1C =
  1.187434e-13, 1.190692e-13, 1.190059e-13, 1.192685e-13, 1.191229e-13, 
    1.192948e-13, 1.188095e-13, 1.190821e-13, 1.189081e-13, 1.187728e-13, 
    1.197775e-13, 1.192802e-13, 1.202939e-13, 1.199771e-13, 1.207725e-13, 
    1.202445e-13, 1.208789e-13, 1.207574e-13, 1.211232e-13, 1.210185e-13, 
    1.214857e-13, 1.211716e-13, 1.217279e-13, 1.214108e-13, 1.214604e-13, 
    1.211612e-13, 1.193805e-13, 1.197156e-13, 1.193606e-13, 1.194084e-13, 
    1.193869e-13, 1.191259e-13, 1.189942e-13, 1.187186e-13, 1.187686e-13, 
    1.189711e-13, 1.194299e-13, 1.192743e-13, 1.196666e-13, 1.196577e-13, 
    1.200939e-13, 1.198973e-13, 1.206299e-13, 1.204218e-13, 1.210228e-13, 
    1.208718e-13, 1.210157e-13, 1.209721e-13, 1.210163e-13, 1.207947e-13, 
    1.208896e-13, 1.206946e-13, 1.199341e-13, 1.201577e-13, 1.194903e-13, 
    1.190884e-13, 1.188214e-13, 1.186319e-13, 1.186587e-13, 1.187097e-13, 
    1.189723e-13, 1.19219e-13, 1.19407e-13, 1.195326e-13, 1.196564e-13, 
    1.200306e-13, 1.202287e-13, 1.206719e-13, 1.20592e-13, 1.207274e-13, 
    1.208567e-13, 1.210737e-13, 1.21038e-13, 1.211335e-13, 1.207239e-13, 
    1.209961e-13, 1.205465e-13, 1.206695e-13, 1.196897e-13, 1.193163e-13, 
    1.191571e-13, 1.190181e-13, 1.186793e-13, 1.189132e-13, 1.18821e-13, 
    1.190405e-13, 1.191798e-13, 1.191109e-13, 1.195361e-13, 1.193708e-13, 
    1.202405e-13, 1.198661e-13, 1.208416e-13, 1.206084e-13, 1.208975e-13, 
    1.207501e-13, 1.210027e-13, 1.207753e-13, 1.211691e-13, 1.212548e-13, 
    1.211962e-13, 1.214212e-13, 1.207627e-13, 1.210157e-13, 1.19109e-13, 
    1.191202e-13, 1.191726e-13, 1.189423e-13, 1.189282e-13, 1.187172e-13, 
    1.18905e-13, 1.189849e-13, 1.191879e-13, 1.193079e-13, 1.194219e-13, 
    1.196725e-13, 1.199521e-13, 1.20343e-13, 1.206236e-13, 1.208115e-13, 
    1.206963e-13, 1.20798e-13, 1.206843e-13, 1.20631e-13, 1.212227e-13, 
    1.208905e-13, 1.213888e-13, 1.213613e-13, 1.211358e-13, 1.213644e-13, 
    1.191281e-13, 1.190634e-13, 1.188387e-13, 1.190146e-13, 1.186942e-13, 
    1.188735e-13, 1.189766e-13, 1.193742e-13, 1.194616e-13, 1.195425e-13, 
    1.197024e-13, 1.199074e-13, 1.202667e-13, 1.205792e-13, 1.208643e-13, 
    1.208434e-13, 1.208507e-13, 1.209144e-13, 1.207567e-13, 1.209402e-13, 
    1.20971e-13, 1.208905e-13, 1.213576e-13, 1.212242e-13, 1.213607e-13, 
    1.212739e-13, 1.190845e-13, 1.191933e-13, 1.191345e-13, 1.19245e-13, 
    1.191671e-13, 1.195133e-13, 1.196171e-13, 1.201023e-13, 1.199033e-13, 
    1.2022e-13, 1.199355e-13, 1.199859e-13, 1.202302e-13, 1.199509e-13, 
    1.205619e-13, 1.201476e-13, 1.209168e-13, 1.205034e-13, 1.209427e-13, 
    1.20863e-13, 1.20995e-13, 1.211131e-13, 1.212617e-13, 1.215356e-13, 
    1.214722e-13, 1.217012e-13, 1.193555e-13, 1.194965e-13, 1.194842e-13, 
    1.196317e-13, 1.197408e-13, 1.199772e-13, 1.203561e-13, 1.202137e-13, 
    1.204751e-13, 1.205276e-13, 1.201304e-13, 1.203742e-13, 1.195909e-13, 
    1.197175e-13, 1.196422e-13, 1.193666e-13, 1.202464e-13, 1.197951e-13, 
    1.206282e-13, 1.20384e-13, 1.210962e-13, 1.207421e-13, 1.214373e-13, 
    1.217339e-13, 1.220131e-13, 1.223388e-13, 1.195735e-13, 1.194777e-13, 
    1.196493e-13, 1.198864e-13, 1.201065e-13, 1.203989e-13, 1.204288e-13, 
    1.204835e-13, 1.206253e-13, 1.207444e-13, 1.205008e-13, 1.207743e-13, 
    1.197467e-13, 1.202856e-13, 1.194414e-13, 1.196957e-13, 1.198725e-13, 
    1.19795e-13, 1.201974e-13, 1.202922e-13, 1.20677e-13, 1.204782e-13, 
    1.216606e-13, 1.211379e-13, 1.225868e-13, 1.221825e-13, 1.194442e-13, 
    1.195732e-13, 1.200217e-13, 1.198084e-13, 1.204184e-13, 1.205684e-13, 
    1.206903e-13, 1.20846e-13, 1.208629e-13, 1.209551e-13, 1.20804e-13, 
    1.209492e-13, 1.203995e-13, 1.206452e-13, 1.199706e-13, 1.201349e-13, 
    1.200593e-13, 1.199764e-13, 1.202323e-13, 1.205046e-13, 1.205105e-13, 
    1.205977e-13, 1.208433e-13, 1.204209e-13, 1.217278e-13, 1.20921e-13, 
    1.197138e-13, 1.199619e-13, 1.199975e-13, 1.199014e-13, 1.205533e-13, 
    1.203172e-13, 1.209529e-13, 1.207812e-13, 1.210625e-13, 1.209227e-13, 
    1.209022e-13, 1.207226e-13, 1.206108e-13, 1.20328e-13, 1.200979e-13, 
    1.199153e-13, 1.199578e-13, 1.201583e-13, 1.205212e-13, 1.208644e-13, 
    1.207892e-13, 1.210411e-13, 1.203742e-13, 1.206539e-13, 1.205458e-13, 
    1.208277e-13, 1.202099e-13, 1.207357e-13, 1.200753e-13, 1.201333e-13, 
    1.203125e-13, 1.206728e-13, 1.207527e-13, 1.208377e-13, 1.207852e-13, 
    1.205305e-13, 1.204888e-13, 1.203082e-13, 1.202583e-13, 1.201207e-13, 
    1.200067e-13, 1.201108e-13, 1.202201e-13, 1.205306e-13, 1.208102e-13, 
    1.211148e-13, 1.211893e-13, 1.215445e-13, 1.212552e-13, 1.217323e-13, 
    1.213265e-13, 1.220288e-13, 1.207663e-13, 1.213148e-13, 1.203207e-13, 
    1.20428e-13, 1.206217e-13, 1.210661e-13, 1.208264e-13, 1.211067e-13, 
    1.204871e-13, 1.201652e-13, 1.20082e-13, 1.199264e-13, 1.200855e-13, 
    1.200726e-13, 1.202247e-13, 1.201759e-13, 1.205409e-13, 1.203449e-13, 
    1.209016e-13, 1.211045e-13, 1.216772e-13, 1.220277e-13, 1.223844e-13, 
    1.225416e-13, 1.225895e-13, 1.226095e-13 ;

 LITR2C_vr =
  0.001107539, 0.001107538, 0.001107538, 0.001107537, 0.001107538, 
    0.001107537, 0.001107539, 0.001107538, 0.001107538, 0.001107539, 
    0.001107535, 0.001107537, 0.001107534, 0.001107535, 0.001107532, 
    0.001107534, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.001107531, 0.001107529, 0.00110753, 0.00110753, 
    0.001107531, 0.001107537, 0.001107536, 0.001107537, 0.001107537, 
    0.001107537, 0.001107538, 0.001107538, 0.001107539, 0.001107539, 
    0.001107538, 0.001107537, 0.001107537, 0.001107536, 0.001107536, 
    0.001107534, 0.001107535, 0.001107532, 0.001107533, 0.001107531, 
    0.001107532, 0.001107531, 0.001107531, 0.001107531, 0.001107532, 
    0.001107531, 0.001107532, 0.001107535, 0.001107534, 0.001107536, 
    0.001107538, 0.001107539, 0.001107539, 0.001107539, 0.001107539, 
    0.001107538, 0.001107537, 0.001107537, 0.001107536, 0.001107536, 
    0.001107535, 0.001107534, 0.001107532, 0.001107533, 0.001107532, 
    0.001107532, 0.001107531, 0.001107531, 0.001107531, 0.001107532, 
    0.001107531, 0.001107533, 0.001107532, 0.001107536, 0.001107537, 
    0.001107538, 0.001107538, 0.001107539, 0.001107538, 0.001107539, 
    0.001107538, 0.001107537, 0.001107538, 0.001107536, 0.001107537, 
    0.001107534, 0.001107535, 0.001107532, 0.001107533, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.00110753, 
    0.00110753, 0.00110753, 0.001107532, 0.001107531, 0.001107538, 
    0.001107538, 0.001107537, 0.001107538, 0.001107538, 0.001107539, 
    0.001107538, 0.001107538, 0.001107537, 0.001107537, 0.001107537, 
    0.001107536, 0.001107535, 0.001107533, 0.001107532, 0.001107532, 
    0.001107532, 0.001107532, 0.001107532, 0.001107532, 0.00110753, 
    0.001107531, 0.00110753, 0.00110753, 0.001107531, 0.00110753, 
    0.001107538, 0.001107538, 0.001107539, 0.001107538, 0.001107539, 
    0.001107538, 0.001107538, 0.001107537, 0.001107536, 0.001107536, 
    0.001107536, 0.001107535, 0.001107534, 0.001107533, 0.001107532, 
    0.001107532, 0.001107532, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.00110753, 0.00110753, 0.00110753, 
    0.001107538, 0.001107537, 0.001107538, 0.001107537, 0.001107538, 
    0.001107536, 0.001107536, 0.001107534, 0.001107535, 0.001107534, 
    0.001107535, 0.001107535, 0.001107534, 0.001107535, 0.001107533, 
    0.001107534, 0.001107531, 0.001107533, 0.001107531, 0.001107532, 
    0.001107531, 0.001107531, 0.00110753, 0.001107529, 0.00110753, 
    0.001107529, 0.001107537, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107535, 0.001107533, 0.001107534, 0.001107533, 
    0.001107533, 0.001107534, 0.001107533, 0.001107536, 0.001107536, 
    0.001107536, 0.001107537, 0.001107534, 0.001107535, 0.001107532, 
    0.001107533, 0.001107531, 0.001107532, 0.00110753, 0.001107529, 
    0.001107528, 0.001107526, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107533, 
    0.001107532, 0.001107532, 0.001107533, 0.001107532, 0.001107535, 
    0.001107534, 0.001107536, 0.001107536, 0.001107535, 0.001107535, 
    0.001107534, 0.001107534, 0.001107532, 0.001107533, 0.001107529, 
    0.001107531, 0.001107526, 0.001107527, 0.001107536, 0.001107536, 
    0.001107535, 0.001107535, 0.001107533, 0.001107533, 0.001107532, 
    0.001107532, 0.001107532, 0.001107531, 0.001107532, 0.001107531, 
    0.001107533, 0.001107532, 0.001107535, 0.001107534, 0.001107534, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107533, 
    0.001107532, 0.001107533, 0.001107529, 0.001107531, 0.001107536, 
    0.001107535, 0.001107535, 0.001107535, 0.001107533, 0.001107533, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.001107531, 
    0.001107532, 0.001107532, 0.001107533, 0.001107534, 0.001107535, 
    0.001107535, 0.001107534, 0.001107533, 0.001107532, 0.001107532, 
    0.001107531, 0.001107533, 0.001107532, 0.001107533, 0.001107532, 
    0.001107534, 0.001107532, 0.001107534, 0.001107534, 0.001107533, 
    0.001107532, 0.001107532, 0.001107532, 0.001107532, 0.001107533, 
    0.001107533, 0.001107534, 0.001107534, 0.001107534, 0.001107535, 
    0.001107534, 0.001107534, 0.001107533, 0.001107532, 0.001107531, 
    0.00110753, 0.001107529, 0.00110753, 0.001107529, 0.00110753, 
    0.001107528, 0.001107532, 0.00110753, 0.001107533, 0.001107533, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.001107533, 
    0.001107534, 0.001107534, 0.001107535, 0.001107534, 0.001107534, 
    0.001107534, 0.001107534, 0.001107533, 0.001107533, 0.001107531, 
    0.001107531, 0.001107529, 0.001107528, 0.001107526, 0.001107526, 
    0.001107526, 0.001107526,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684282e-07, 2.684279e-07, 2.684279e-07, 2.684277e-07, 2.684278e-07, 
    2.684277e-07, 2.684281e-07, 2.684279e-07, 2.68428e-07, 2.684281e-07, 
    2.684273e-07, 2.684277e-07, 2.684268e-07, 2.684271e-07, 2.684264e-07, 
    2.684269e-07, 2.684264e-07, 2.684264e-07, 2.684261e-07, 2.684262e-07, 
    2.684259e-07, 2.684261e-07, 2.684256e-07, 2.684259e-07, 2.684259e-07, 
    2.684261e-07, 2.684276e-07, 2.684273e-07, 2.684276e-07, 2.684276e-07, 
    2.684276e-07, 2.684278e-07, 2.68428e-07, 2.684282e-07, 2.684281e-07, 
    2.68428e-07, 2.684276e-07, 2.684277e-07, 2.684274e-07, 2.684274e-07, 
    2.68427e-07, 2.684272e-07, 2.684266e-07, 2.684267e-07, 2.684262e-07, 
    2.684264e-07, 2.684262e-07, 2.684263e-07, 2.684262e-07, 2.684264e-07, 
    2.684263e-07, 2.684265e-07, 2.684272e-07, 2.68427e-07, 2.684275e-07, 
    2.684279e-07, 2.684281e-07, 2.684282e-07, 2.684282e-07, 2.684282e-07, 
    2.68428e-07, 2.684278e-07, 2.684276e-07, 2.684275e-07, 2.684274e-07, 
    2.684271e-07, 2.684269e-07, 2.684265e-07, 2.684266e-07, 2.684265e-07, 
    2.684264e-07, 2.684262e-07, 2.684262e-07, 2.684261e-07, 2.684265e-07, 
    2.684262e-07, 2.684266e-07, 2.684265e-07, 2.684274e-07, 2.684277e-07, 
    2.684278e-07, 2.684279e-07, 2.684282e-07, 2.68428e-07, 2.684281e-07, 
    2.684279e-07, 2.684278e-07, 2.684278e-07, 2.684275e-07, 2.684276e-07, 
    2.684269e-07, 2.684272e-07, 2.684264e-07, 2.684266e-07, 2.684263e-07, 
    2.684265e-07, 2.684262e-07, 2.684264e-07, 2.684261e-07, 2.68426e-07, 
    2.684261e-07, 2.684259e-07, 2.684264e-07, 2.684262e-07, 2.684278e-07, 
    2.684278e-07, 2.684278e-07, 2.68428e-07, 2.68428e-07, 2.684282e-07, 
    2.68428e-07, 2.68428e-07, 2.684278e-07, 2.684277e-07, 2.684276e-07, 
    2.684274e-07, 2.684271e-07, 2.684268e-07, 2.684266e-07, 2.684264e-07, 
    2.684265e-07, 2.684264e-07, 2.684265e-07, 2.684266e-07, 2.684261e-07, 
    2.684263e-07, 2.684259e-07, 2.684259e-07, 2.684261e-07, 2.684259e-07, 
    2.684278e-07, 2.684279e-07, 2.684281e-07, 2.684279e-07, 2.684282e-07, 
    2.68428e-07, 2.68428e-07, 2.684276e-07, 2.684276e-07, 2.684275e-07, 
    2.684274e-07, 2.684272e-07, 2.684269e-07, 2.684266e-07, 2.684264e-07, 
    2.684264e-07, 2.684264e-07, 2.684263e-07, 2.684264e-07, 2.684263e-07, 
    2.684263e-07, 2.684263e-07, 2.684259e-07, 2.68426e-07, 2.684259e-07, 
    2.68426e-07, 2.684279e-07, 2.684278e-07, 2.684278e-07, 2.684277e-07, 
    2.684278e-07, 2.684275e-07, 2.684274e-07, 2.68427e-07, 2.684272e-07, 
    2.684269e-07, 2.684272e-07, 2.684271e-07, 2.684269e-07, 2.684271e-07, 
    2.684266e-07, 2.68427e-07, 2.684263e-07, 2.684267e-07, 2.684263e-07, 
    2.684264e-07, 2.684262e-07, 2.684262e-07, 2.68426e-07, 2.684258e-07, 
    2.684259e-07, 2.684257e-07, 2.684276e-07, 2.684275e-07, 2.684275e-07, 
    2.684274e-07, 2.684273e-07, 2.684271e-07, 2.684268e-07, 2.684269e-07, 
    2.684267e-07, 2.684266e-07, 2.68427e-07, 2.684268e-07, 2.684274e-07, 
    2.684273e-07, 2.684274e-07, 2.684276e-07, 2.684269e-07, 2.684273e-07, 
    2.684266e-07, 2.684268e-07, 2.684262e-07, 2.684265e-07, 2.684259e-07, 
    2.684256e-07, 2.684254e-07, 2.684251e-07, 2.684274e-07, 2.684275e-07, 
    2.684274e-07, 2.684272e-07, 2.68427e-07, 2.684268e-07, 2.684267e-07, 
    2.684267e-07, 2.684266e-07, 2.684265e-07, 2.684267e-07, 2.684264e-07, 
    2.684273e-07, 2.684268e-07, 2.684276e-07, 2.684274e-07, 2.684272e-07, 
    2.684273e-07, 2.684269e-07, 2.684268e-07, 2.684265e-07, 2.684267e-07, 
    2.684257e-07, 2.684261e-07, 2.684249e-07, 2.684253e-07, 2.684276e-07, 
    2.684274e-07, 2.684271e-07, 2.684272e-07, 2.684267e-07, 2.684266e-07, 
    2.684265e-07, 2.684264e-07, 2.684264e-07, 2.684263e-07, 2.684264e-07, 
    2.684263e-07, 2.684268e-07, 2.684266e-07, 2.684271e-07, 2.68427e-07, 
    2.68427e-07, 2.684271e-07, 2.684269e-07, 2.684267e-07, 2.684267e-07, 
    2.684266e-07, 2.684264e-07, 2.684267e-07, 2.684257e-07, 2.684263e-07, 
    2.684273e-07, 2.684271e-07, 2.684271e-07, 2.684272e-07, 2.684266e-07, 
    2.684268e-07, 2.684263e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 
    2.684263e-07, 2.684265e-07, 2.684266e-07, 2.684268e-07, 2.68427e-07, 
    2.684272e-07, 2.684271e-07, 2.68427e-07, 2.684266e-07, 2.684264e-07, 
    2.684264e-07, 2.684262e-07, 2.684268e-07, 2.684265e-07, 2.684266e-07, 
    2.684264e-07, 2.684269e-07, 2.684265e-07, 2.68427e-07, 2.68427e-07, 
    2.684268e-07, 2.684265e-07, 2.684264e-07, 2.684264e-07, 2.684264e-07, 
    2.684266e-07, 2.684267e-07, 2.684268e-07, 2.684269e-07, 2.68427e-07, 
    2.684271e-07, 2.68427e-07, 2.684269e-07, 2.684266e-07, 2.684264e-07, 
    2.684262e-07, 2.684261e-07, 2.684258e-07, 2.68426e-07, 2.684256e-07, 
    2.68426e-07, 2.684254e-07, 2.684264e-07, 2.68426e-07, 2.684268e-07, 
    2.684267e-07, 2.684266e-07, 2.684262e-07, 2.684264e-07, 2.684262e-07, 
    2.684267e-07, 2.68427e-07, 2.68427e-07, 2.684272e-07, 2.68427e-07, 
    2.68427e-07, 2.684269e-07, 2.68427e-07, 2.684266e-07, 2.684268e-07, 
    2.684263e-07, 2.684262e-07, 2.684257e-07, 2.684254e-07, 2.684251e-07, 
    2.684249e-07, 2.684249e-07, 2.684249e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -2.695996e-26, 9.313441e-26, -1.960724e-26, 1.053889e-25, -6.127264e-26, 
    5.391992e-26, 1.519561e-25, -1.127417e-25, -1.29898e-25, -2.941087e-26, 
    -2.08327e-25, 1.151926e-25, 2.450905e-26, -2.450906e-27, 9.068351e-26, 
    1.936215e-25, 2.401887e-25, 4.901811e-27, 2.450905e-26, -1.764652e-25, 
    9.803622e-26, -8.82326e-26, 4.166539e-26, -3.186177e-25, -2.450906e-27, 
    7.597807e-26, -6.617445e-26, 5.146902e-26, -1.102908e-25, 2.794032e-25, 
    1.151926e-25, -1.078398e-25, 3.088141e-25, 1.421525e-25, -6.372354e-26, 
    6.862535e-26, 2.499924e-25, 5.882173e-26, -1.397016e-25, 2.279342e-25, 
    1.053889e-25, 1.691125e-25, 2.058761e-25, 2.745014e-25, -1.838179e-25, 
    8.82326e-26, -7.107626e-26, -1.715634e-25, -1.470543e-25, 1.004871e-25, 
    -9.803622e-27, 8.82326e-26, 1.470543e-26, -9.068351e-26, -4.901811e-27, 
    -6.862535e-26, 1.911706e-25, 1.960724e-26, 1.530638e-41, -2.450905e-26, 
    2.450905e-26, -2.499924e-25, 7.352717e-27, 1.960724e-25, 4.901811e-26, 
    -3.186177e-26, 5.882173e-26, -2.377378e-25, -6.127264e-26, -1.715634e-25, 
    -3.921449e-26, 7.352717e-26, 2.941087e-26, -2.941087e-26, 2.695996e-25, 
    -1.176435e-25, -1.078398e-25, 1.053889e-25, -2.695996e-26, 3.921449e-26, 
    1.519561e-25, -7.352717e-26, 2.279342e-25, 1.004871e-25, -7.352717e-26, 
    1.249962e-25, 7.352717e-26, 3.676358e-26, -1.446034e-25, 2.426396e-25, 
    4.65672e-26, -7.352717e-26, -4.65672e-26, 1.02938e-25, -1.225453e-25, 
    -1.519561e-25, -1.715634e-26, 1.495052e-25, -4.043994e-25, -3.431268e-26, 
    -4.901811e-26, 1.911706e-25, -9.313441e-26, 7.597807e-26, 2.181306e-25, 
    -2.009742e-25, -9.558531e-26, 1.421525e-25, -8.087988e-26, 5.146902e-26, 
    1.446034e-25, -8.333079e-26, 1.127417e-25, -1.519561e-25, -9.803622e-26, 
    -3.431268e-26, -8.333079e-26, -2.450906e-27, 1.127417e-25, 5.391992e-26, 
    1.519561e-25, -6.617445e-26, 2.426396e-25, 2.254833e-25, 1.225453e-25, 
    5.637083e-26, -6.372354e-26, -1.29898e-25, -1.078398e-25, -1.004871e-25, 
    -1.691125e-25, -2.205815e-26, -1.862688e-25, -6.372354e-26, -4.65672e-26, 
    4.65672e-26, 3.308722e-25, 1.127417e-25, -4.65672e-26, -3.431268e-26, 
    3.921449e-26, -1.81367e-25, -1.02938e-25, -1.225453e-26, -3.676358e-26, 
    -4.65672e-26, -9.068351e-26, -8.087988e-26, 2.08327e-25, 5.391992e-26, 
    -4.65672e-26, 6.127264e-26, -2.450906e-27, -2.695996e-25, -1.642107e-25, 
    0, -1.985233e-25, 2.818541e-25, -2.132288e-25, -2.475414e-25, 
    1.29898e-25, 3.921449e-26, -9.558531e-26, -3.431268e-26, 9.068351e-26, 
    -6.127264e-26, 3.431268e-26, 7.842898e-26, 1.200944e-25, -5.391992e-26, 
    -7.352717e-27, -1.715634e-26, 1.274471e-25, -6.372354e-26, 8.087988e-26, 
    6.372354e-26, -1.078398e-25, 2.941087e-26, -1.078398e-25, -1.740143e-25, 
    1.249962e-25, -3.431268e-26, -1.004871e-25, 1.715634e-26, 2.377378e-25, 
    -3.186177e-26, 2.205815e-26, -1.053889e-25, -4.65672e-26, -4.901811e-27, 
    1.715634e-26, 1.666616e-25, -1.225453e-26, 1.838179e-25, 1.715634e-25, 
    1.127417e-25, -9.803622e-27, 2.843051e-25, -1.936215e-25, -6.862535e-26, 
    2.450905e-26, 1.274471e-25, 1.02938e-25, -2.107779e-25, 1.02938e-25, 
    4.65672e-26, -6.862535e-26, 1.372507e-25, -9.558531e-26, 1.02938e-25, 
    -8.578169e-26, -1.200944e-25, -4.41163e-26, 2.230324e-25, -8.578169e-26, 
    1.56858e-25, -2.254833e-25, -1.470543e-26, -3.921449e-26, 2.794032e-25, 
    8.333079e-26, -6.372354e-26, 3.088141e-25, 1.225453e-26, 2.59796e-25, 
    -1.078398e-25, 3.431268e-26, 1.249962e-25, 6.127264e-26, -5.391992e-26, 
    -1.740143e-25, 1.887197e-25, 1.54407e-25, 1.81367e-25, 1.715634e-26, 
    -6.372354e-26, -2.230324e-25, -1.470543e-26, 1.54407e-25, -1.397016e-25, 
    -1.323489e-25, -2.720505e-25, -2.08327e-25, 4.41163e-26, 2.695996e-26, 
    1.421525e-25, 1.960724e-25, -8.087988e-26, 6.372354e-26, 2.941087e-26, 
    -1.470543e-26, 3.186177e-26, 1.347998e-25, -9.803622e-26, 1.446034e-25, 
    -1.421525e-25, 1.642107e-25, 5.391992e-26, 9.558531e-26, 5.882173e-26, 
    -2.107779e-25, 3.308722e-25, 2.450906e-27, -1.176435e-25, -2.058761e-25, 
    5.391992e-26, 8.087988e-26, -5.882173e-26, 2.941087e-26, 1.200944e-25, 
    8.087988e-26, -1.960724e-26, 7.352717e-26, -2.450905e-26, 1.960724e-26, 
    -7.597807e-26, -1.593089e-25, -5.146902e-26, 3.921449e-26, -1.102908e-25, 
    1.470543e-26, 8.82326e-26, -1.470543e-26, -9.803622e-26, -7.352717e-26, 
    -1.740143e-25, 1.29898e-25, 1.004871e-25, -9.558531e-26, -7.597807e-26, 
    2.107779e-25, 1.323489e-25, 1.740143e-25, 7.352717e-27, 6.617445e-26, 
    1.372507e-25, 7.842898e-26, 6.617445e-26, 3.921449e-26, 1.642107e-25, 
    -1.495052e-25, -1.911706e-25, 2.818541e-25, -8.333079e-26, 1.715634e-25, 
    1.530638e-41, -3.431268e-26, 7.597807e-26, -1.127417e-25, -8.087988e-26, 
    -1.54407e-25, 1.323489e-25, -2.941087e-26, -4.65672e-26, 2.009742e-25, 
    1.715634e-26, -3.872431e-25, 1.740143e-25, -6.862535e-26, 1.56858e-25, 
    1.004871e-25, -4.65672e-26, 8.82326e-26, 7.597807e-26, -8.333079e-26, 
    -7.597807e-26, 1.56858e-25, -5.146902e-26, -4.166539e-26, 8.82326e-26, 
    -2.205815e-26, -3.088141e-25, -7.107626e-26, 2.230324e-25, 4.41163e-26, 
    -1.715634e-26, -1.666616e-25, -4.65672e-26,
  2.676268e-32, 2.676265e-32, 2.676266e-32, 2.676263e-32, 2.676265e-32, 
    2.676263e-32, 2.676267e-32, 2.676265e-32, 2.676267e-32, 2.676268e-32, 
    2.676259e-32, 2.676263e-32, 2.676255e-32, 2.676257e-32, 2.676251e-32, 
    2.676255e-32, 2.67625e-32, 2.676251e-32, 2.676248e-32, 2.676249e-32, 
    2.676244e-32, 2.676247e-32, 2.676242e-32, 2.676245e-32, 2.676245e-32, 
    2.676247e-32, 2.676262e-32, 2.67626e-32, 2.676263e-32, 2.676262e-32, 
    2.676262e-32, 2.676265e-32, 2.676266e-32, 2.676268e-32, 2.676268e-32, 
    2.676266e-32, 2.676262e-32, 2.676263e-32, 2.67626e-32, 2.67626e-32, 
    2.676257e-32, 2.676258e-32, 2.676252e-32, 2.676254e-32, 2.676249e-32, 
    2.67625e-32, 2.676249e-32, 2.676249e-32, 2.676249e-32, 2.67625e-32, 
    2.67625e-32, 2.676251e-32, 2.676258e-32, 2.676256e-32, 2.676262e-32, 
    2.676265e-32, 2.676267e-32, 2.676269e-32, 2.676269e-32, 2.676268e-32, 
    2.676266e-32, 2.676264e-32, 2.676262e-32, 2.676261e-32, 2.67626e-32, 
    2.676257e-32, 2.676255e-32, 2.676252e-32, 2.676252e-32, 2.676251e-32, 
    2.67625e-32, 2.676248e-32, 2.676248e-32, 2.676248e-32, 2.676251e-32, 
    2.676249e-32, 2.676253e-32, 2.676252e-32, 2.67626e-32, 2.676263e-32, 
    2.676264e-32, 2.676266e-32, 2.676268e-32, 2.676267e-32, 2.676267e-32, 
    2.676265e-32, 2.676264e-32, 2.676265e-32, 2.676261e-32, 2.676262e-32, 
    2.676255e-32, 2.676258e-32, 2.67625e-32, 2.676252e-32, 2.676249e-32, 
    2.676251e-32, 2.676249e-32, 2.676251e-32, 2.676247e-32, 2.676247e-32, 
    2.676247e-32, 2.676245e-32, 2.676251e-32, 2.676249e-32, 2.676265e-32, 
    2.676265e-32, 2.676264e-32, 2.676266e-32, 2.676266e-32, 2.676268e-32, 
    2.676267e-32, 2.676266e-32, 2.676264e-32, 2.676263e-32, 2.676262e-32, 
    2.67626e-32, 2.676258e-32, 2.676254e-32, 2.676252e-32, 2.67625e-32, 
    2.676251e-32, 2.67625e-32, 2.676252e-32, 2.676252e-32, 2.676247e-32, 
    2.67625e-32, 2.676245e-32, 2.676246e-32, 2.676248e-32, 2.676246e-32, 
    2.676264e-32, 2.676265e-32, 2.676267e-32, 2.676266e-32, 2.676268e-32, 
    2.676267e-32, 2.676266e-32, 2.676262e-32, 2.676262e-32, 2.676261e-32, 
    2.67626e-32, 2.676258e-32, 2.676255e-32, 2.676252e-32, 2.67625e-32, 
    2.67625e-32, 2.67625e-32, 2.676249e-32, 2.676251e-32, 2.676249e-32, 
    2.676249e-32, 2.67625e-32, 2.676246e-32, 2.676247e-32, 2.676246e-32, 
    2.676247e-32, 2.676265e-32, 2.676264e-32, 2.676264e-32, 2.676264e-32, 
    2.676264e-32, 2.676261e-32, 2.67626e-32, 2.676256e-32, 2.676258e-32, 
    2.676255e-32, 2.676258e-32, 2.676257e-32, 2.676255e-32, 2.676258e-32, 
    2.676252e-32, 2.676256e-32, 2.676249e-32, 2.676253e-32, 2.676249e-32, 
    2.67625e-32, 2.676249e-32, 2.676248e-32, 2.676247e-32, 2.676244e-32, 
    2.676245e-32, 2.676243e-32, 2.676263e-32, 2.676262e-32, 2.676262e-32, 
    2.67626e-32, 2.676259e-32, 2.676257e-32, 2.676254e-32, 2.676255e-32, 
    2.676253e-32, 2.676253e-32, 2.676256e-32, 2.676254e-32, 2.676261e-32, 
    2.676259e-32, 2.67626e-32, 2.676263e-32, 2.676255e-32, 2.676259e-32, 
    2.676252e-32, 2.676254e-32, 2.676248e-32, 2.676251e-32, 2.676245e-32, 
    2.676242e-32, 2.67624e-32, 2.676237e-32, 2.676261e-32, 2.676262e-32, 
    2.67626e-32, 2.676258e-32, 2.676256e-32, 2.676254e-32, 2.676254e-32, 
    2.676253e-32, 2.676252e-32, 2.676251e-32, 2.676253e-32, 2.676251e-32, 
    2.676259e-32, 2.676255e-32, 2.676262e-32, 2.67626e-32, 2.676258e-32, 
    2.676259e-32, 2.676256e-32, 2.676255e-32, 2.676252e-32, 2.676253e-32, 
    2.676243e-32, 2.676248e-32, 2.676235e-32, 2.676239e-32, 2.676262e-32, 
    2.676261e-32, 2.676257e-32, 2.676259e-32, 2.676254e-32, 2.676252e-32, 
    2.676251e-32, 2.67625e-32, 2.67625e-32, 2.676249e-32, 2.67625e-32, 
    2.676249e-32, 2.676254e-32, 2.676252e-32, 2.676257e-32, 2.676256e-32, 
    2.676257e-32, 2.676257e-32, 2.676255e-32, 2.676253e-32, 2.676253e-32, 
    2.676252e-32, 2.67625e-32, 2.676254e-32, 2.676243e-32, 2.676249e-32, 
    2.67626e-32, 2.676257e-32, 2.676257e-32, 2.676258e-32, 2.676252e-32, 
    2.676254e-32, 2.676249e-32, 2.676251e-32, 2.676248e-32, 2.676249e-32, 
    2.676249e-32, 2.676251e-32, 2.676252e-32, 2.676254e-32, 2.676257e-32, 
    2.676258e-32, 2.676258e-32, 2.676256e-32, 2.676253e-32, 2.67625e-32, 
    2.676251e-32, 2.676248e-32, 2.676254e-32, 2.676252e-32, 2.676253e-32, 
    2.67625e-32, 2.676255e-32, 2.676251e-32, 2.676257e-32, 2.676256e-32, 
    2.676254e-32, 2.676252e-32, 2.676251e-32, 2.67625e-32, 2.676251e-32, 
    2.676253e-32, 2.676253e-32, 2.676254e-32, 2.676255e-32, 2.676256e-32, 
    2.676257e-32, 2.676256e-32, 2.676255e-32, 2.676253e-32, 2.67625e-32, 
    2.676248e-32, 2.676247e-32, 2.676244e-32, 2.676247e-32, 2.676242e-32, 
    2.676246e-32, 2.67624e-32, 2.676251e-32, 2.676246e-32, 2.676254e-32, 
    2.676254e-32, 2.676252e-32, 2.676248e-32, 2.67625e-32, 2.676248e-32, 
    2.676253e-32, 2.676256e-32, 2.676257e-32, 2.676258e-32, 2.676257e-32, 
    2.676257e-32, 2.676255e-32, 2.676256e-32, 2.676253e-32, 2.676254e-32, 
    2.676249e-32, 2.676248e-32, 2.676243e-32, 2.67624e-32, 2.676237e-32, 
    2.676236e-32, 2.676235e-32, 2.676235e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.286642e-15, 3.29566e-15, 3.293909e-15, 3.301177e-15, 3.297147e-15, 
    3.301904e-15, 3.288473e-15, 3.296017e-15, 3.291202e-15, 3.287456e-15, 
    3.315265e-15, 3.301501e-15, 3.329557e-15, 3.32079e-15, 3.342805e-15, 
    3.328192e-15, 3.345749e-15, 3.342387e-15, 3.352513e-15, 3.349613e-15, 
    3.362547e-15, 3.353851e-15, 3.36925e-15, 3.360472e-15, 3.361845e-15, 
    3.353563e-15, 3.304276e-15, 3.313551e-15, 3.303725e-15, 3.305048e-15, 
    3.304455e-15, 3.297229e-15, 3.293583e-15, 3.285955e-15, 3.287341e-15, 
    3.292945e-15, 3.305643e-15, 3.301336e-15, 3.312194e-15, 3.311949e-15, 
    3.324023e-15, 3.318581e-15, 3.338858e-15, 3.333099e-15, 3.349734e-15, 
    3.345553e-15, 3.349537e-15, 3.348329e-15, 3.349553e-15, 3.34342e-15, 
    3.346048e-15, 3.34065e-15, 3.3196e-15, 3.32579e-15, 3.307317e-15, 
    3.296191e-15, 3.288803e-15, 3.283555e-15, 3.284297e-15, 3.285711e-15, 
    3.292977e-15, 3.299808e-15, 3.30501e-15, 3.308488e-15, 3.311914e-15, 
    3.32227e-15, 3.327755e-15, 3.34002e-15, 3.337811e-15, 3.341556e-15, 
    3.345137e-15, 3.351142e-15, 3.350154e-15, 3.352798e-15, 3.341459e-15, 
    3.348995e-15, 3.336551e-15, 3.339956e-15, 3.312834e-15, 3.302499e-15, 
    3.298094e-15, 3.294245e-15, 3.284868e-15, 3.291344e-15, 3.288791e-15, 
    3.294865e-15, 3.298722e-15, 3.296815e-15, 3.308583e-15, 3.304009e-15, 
    3.32808e-15, 3.317718e-15, 3.344719e-15, 3.338264e-15, 3.346266e-15, 
    3.342184e-15, 3.349176e-15, 3.342884e-15, 3.353783e-15, 3.356154e-15, 
    3.354534e-15, 3.360759e-15, 3.342535e-15, 3.349536e-15, 3.296761e-15, 
    3.297072e-15, 3.298522e-15, 3.292147e-15, 3.291758e-15, 3.285917e-15, 
    3.291115e-15, 3.293328e-15, 3.298946e-15, 3.302267e-15, 3.305423e-15, 
    3.312359e-15, 3.320099e-15, 3.330916e-15, 3.338683e-15, 3.343885e-15, 
    3.340696e-15, 3.343512e-15, 3.340364e-15, 3.338889e-15, 3.355265e-15, 
    3.346072e-15, 3.359864e-15, 3.359102e-15, 3.352861e-15, 3.359188e-15, 
    3.297291e-15, 3.295501e-15, 3.289281e-15, 3.294149e-15, 3.28528e-15, 
    3.290244e-15, 3.293096e-15, 3.304102e-15, 3.306521e-15, 3.308761e-15, 
    3.313185e-15, 3.31886e-15, 3.328806e-15, 3.337454e-15, 3.345345e-15, 
    3.344768e-15, 3.344971e-15, 3.346732e-15, 3.342368e-15, 3.347448e-15, 
    3.348299e-15, 3.346072e-15, 3.359e-15, 3.355308e-15, 3.359086e-15, 
    3.356682e-15, 3.296083e-15, 3.299095e-15, 3.297467e-15, 3.300527e-15, 
    3.298371e-15, 3.307953e-15, 3.310824e-15, 3.324254e-15, 3.318747e-15, 
    3.327513e-15, 3.319639e-15, 3.321034e-15, 3.327794e-15, 3.320065e-15, 
    3.336976e-15, 3.32551e-15, 3.3468e-15, 3.335356e-15, 3.347517e-15, 
    3.345311e-15, 3.348964e-15, 3.352232e-15, 3.356345e-15, 3.363927e-15, 
    3.362172e-15, 3.368511e-15, 3.303584e-15, 3.307487e-15, 3.307146e-15, 
    3.31123e-15, 3.31425e-15, 3.320794e-15, 3.33128e-15, 3.327338e-15, 
    3.334575e-15, 3.336026e-15, 3.325033e-15, 3.331782e-15, 3.3101e-15, 
    3.313604e-15, 3.311519e-15, 3.303891e-15, 3.328244e-15, 3.315751e-15, 
    3.338811e-15, 3.332052e-15, 3.351766e-15, 3.341964e-15, 3.361206e-15, 
    3.369415e-15, 3.377145e-15, 3.386158e-15, 3.309619e-15, 3.306968e-15, 
    3.311716e-15, 3.31828e-15, 3.324372e-15, 3.332464e-15, 3.333292e-15, 
    3.334807e-15, 3.338731e-15, 3.342028e-15, 3.335283e-15, 3.342855e-15, 
    3.314412e-15, 3.329328e-15, 3.305963e-15, 3.313001e-15, 3.317894e-15, 
    3.31575e-15, 3.326888e-15, 3.329511e-15, 3.340162e-15, 3.334659e-15, 
    3.367388e-15, 3.35292e-15, 3.393023e-15, 3.381831e-15, 3.306041e-15, 
    3.309611e-15, 3.322026e-15, 3.316121e-15, 3.333005e-15, 3.337156e-15, 
    3.340531e-15, 3.344841e-15, 3.345307e-15, 3.34786e-15, 3.343676e-15, 
    3.347695e-15, 3.332481e-15, 3.339283e-15, 3.32061e-15, 3.325156e-15, 
    3.323066e-15, 3.32077e-15, 3.327852e-15, 3.335389e-15, 3.335553e-15, 
    3.337968e-15, 3.344765e-15, 3.333073e-15, 3.369247e-15, 3.346916e-15, 
    3.313503e-15, 3.32037e-15, 3.321355e-15, 3.318694e-15, 3.33674e-15, 
    3.330204e-15, 3.347798e-15, 3.343047e-15, 3.350832e-15, 3.346964e-15, 
    3.346394e-15, 3.341425e-15, 3.338329e-15, 3.330503e-15, 3.324133e-15, 
    3.319081e-15, 3.320256e-15, 3.325805e-15, 3.335851e-15, 3.345348e-15, 
    3.343268e-15, 3.35024e-15, 3.331781e-15, 3.339524e-15, 3.336531e-15, 
    3.344333e-15, 3.327233e-15, 3.341786e-15, 3.323508e-15, 3.325113e-15, 
    3.330074e-15, 3.340046e-15, 3.342256e-15, 3.344609e-15, 3.343158e-15, 
    3.336106e-15, 3.334952e-15, 3.329955e-15, 3.328573e-15, 3.324764e-15, 
    3.321608e-15, 3.324491e-15, 3.327516e-15, 3.336111e-15, 3.343848e-15, 
    3.352278e-15, 3.354342e-15, 3.364173e-15, 3.356166e-15, 3.369371e-15, 
    3.358138e-15, 3.377578e-15, 3.342634e-15, 3.357815e-15, 3.330301e-15, 
    3.333269e-15, 3.338633e-15, 3.350931e-15, 3.344297e-15, 3.352056e-15, 
    3.334907e-15, 3.325995e-15, 3.323692e-15, 3.319387e-15, 3.32379e-15, 
    3.323432e-15, 3.327644e-15, 3.326291e-15, 3.336396e-15, 3.330969e-15, 
    3.346379e-15, 3.351996e-15, 3.367846e-15, 3.377548e-15, 3.387419e-15, 
    3.391772e-15, 3.393097e-15, 3.393651e-15 ;

 LITR2N_vr =
  1.532753e-05, 1.532751e-05, 1.532751e-05, 1.53275e-05, 1.532751e-05, 
    1.53275e-05, 1.532752e-05, 1.532751e-05, 1.532752e-05, 1.532752e-05, 
    1.532748e-05, 1.53275e-05, 1.532745e-05, 1.532747e-05, 1.532743e-05, 
    1.532745e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.532742e-05, 
    1.532739e-05, 1.532741e-05, 1.532738e-05, 1.53274e-05, 1.532739e-05, 
    1.532741e-05, 1.532749e-05, 1.532748e-05, 1.53275e-05, 1.532749e-05, 
    1.532749e-05, 1.532751e-05, 1.532751e-05, 1.532753e-05, 1.532752e-05, 
    1.532751e-05, 1.532749e-05, 1.53275e-05, 1.532748e-05, 1.532748e-05, 
    1.532746e-05, 1.532747e-05, 1.532743e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 
    1.532742e-05, 1.532743e-05, 1.532747e-05, 1.532746e-05, 1.532749e-05, 
    1.532751e-05, 1.532752e-05, 1.532753e-05, 1.532753e-05, 1.532753e-05, 
    1.532751e-05, 1.53275e-05, 1.532749e-05, 1.532749e-05, 1.532748e-05, 
    1.532746e-05, 1.532745e-05, 1.532743e-05, 1.532744e-05, 1.532743e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532741e-05, 1.532743e-05, 
    1.532742e-05, 1.532744e-05, 1.532743e-05, 1.532748e-05, 1.53275e-05, 
    1.532751e-05, 1.532751e-05, 1.532753e-05, 1.532752e-05, 1.532752e-05, 
    1.532751e-05, 1.53275e-05, 1.532751e-05, 1.532749e-05, 1.532749e-05, 
    1.532745e-05, 1.532747e-05, 1.532742e-05, 1.532744e-05, 1.532742e-05, 
    1.532743e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.53274e-05, 
    1.532741e-05, 1.53274e-05, 1.532743e-05, 1.532742e-05, 1.532751e-05, 
    1.532751e-05, 1.532751e-05, 1.532752e-05, 1.532752e-05, 1.532753e-05, 
    1.532752e-05, 1.532751e-05, 1.53275e-05, 1.53275e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532743e-05, 1.532743e-05, 1.532743e-05, 1.53274e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532741e-05, 1.53274e-05, 
    1.532751e-05, 1.532751e-05, 1.532752e-05, 1.532751e-05, 1.532753e-05, 
    1.532752e-05, 1.532751e-05, 1.532749e-05, 1.532749e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532751e-05, 1.53275e-05, 1.532751e-05, 1.53275e-05, 
    1.532751e-05, 1.532749e-05, 1.532748e-05, 1.532746e-05, 1.532747e-05, 
    1.532745e-05, 1.532747e-05, 1.532747e-05, 1.532745e-05, 1.532747e-05, 
    1.532744e-05, 1.532746e-05, 1.532742e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.53275e-05, 1.532749e-05, 1.532749e-05, 
    1.532748e-05, 1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532745e-05, 
    1.532744e-05, 1.532744e-05, 1.532746e-05, 1.532745e-05, 1.532749e-05, 
    1.532748e-05, 1.532748e-05, 1.53275e-05, 1.532745e-05, 1.532747e-05, 
    1.532743e-05, 1.532745e-05, 1.532741e-05, 1.532743e-05, 1.53274e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532749e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532746e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532743e-05, 1.532743e-05, 1.532744e-05, 1.532743e-05, 
    1.532748e-05, 1.532745e-05, 1.532749e-05, 1.532748e-05, 1.532747e-05, 
    1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532743e-05, 1.532744e-05, 
    1.532738e-05, 1.532741e-05, 1.532734e-05, 1.532736e-05, 1.532749e-05, 
    1.532749e-05, 1.532746e-05, 1.532747e-05, 1.532744e-05, 1.532744e-05, 
    1.532743e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 
    1.532742e-05, 1.532744e-05, 1.532743e-05, 1.532747e-05, 1.532746e-05, 
    1.532746e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532742e-05, 1.532744e-05, 1.532738e-05, 1.532742e-05, 
    1.532748e-05, 1.532747e-05, 1.532747e-05, 1.532747e-05, 1.532744e-05, 
    1.532745e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.532742e-05, 
    1.532742e-05, 1.532743e-05, 1.532744e-05, 1.532745e-05, 1.532746e-05, 
    1.532747e-05, 1.532747e-05, 1.532746e-05, 1.532744e-05, 1.532742e-05, 
    1.532743e-05, 1.532741e-05, 1.532745e-05, 1.532743e-05, 1.532744e-05, 
    1.532742e-05, 1.532745e-05, 1.532743e-05, 1.532746e-05, 1.532746e-05, 
    1.532745e-05, 1.532743e-05, 1.532743e-05, 1.532742e-05, 1.532743e-05, 
    1.532744e-05, 1.532744e-05, 1.532745e-05, 1.532745e-05, 1.532746e-05, 
    1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532744e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 1.532738e-05, 
    1.53274e-05, 1.532737e-05, 1.532743e-05, 1.53274e-05, 1.532745e-05, 
    1.532744e-05, 1.532743e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 
    1.532744e-05, 1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532746e-05, 
    1.532746e-05, 1.532745e-05, 1.532746e-05, 1.532744e-05, 1.532745e-05, 
    1.532742e-05, 1.532741e-05, 1.532738e-05, 1.532737e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532734e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.187434e-13, 1.190692e-13, 1.190059e-13, 1.192685e-13, 1.191229e-13, 
    1.192948e-13, 1.188095e-13, 1.190821e-13, 1.189081e-13, 1.187728e-13, 
    1.197775e-13, 1.192802e-13, 1.202939e-13, 1.199771e-13, 1.207725e-13, 
    1.202445e-13, 1.208789e-13, 1.207574e-13, 1.211232e-13, 1.210185e-13, 
    1.214857e-13, 1.211716e-13, 1.217279e-13, 1.214108e-13, 1.214604e-13, 
    1.211612e-13, 1.193805e-13, 1.197156e-13, 1.193606e-13, 1.194084e-13, 
    1.193869e-13, 1.191259e-13, 1.189942e-13, 1.187186e-13, 1.187686e-13, 
    1.189711e-13, 1.194299e-13, 1.192743e-13, 1.196666e-13, 1.196577e-13, 
    1.200939e-13, 1.198973e-13, 1.206299e-13, 1.204218e-13, 1.210228e-13, 
    1.208718e-13, 1.210157e-13, 1.209721e-13, 1.210163e-13, 1.207947e-13, 
    1.208896e-13, 1.206946e-13, 1.199341e-13, 1.201577e-13, 1.194903e-13, 
    1.190884e-13, 1.188214e-13, 1.186319e-13, 1.186587e-13, 1.187097e-13, 
    1.189723e-13, 1.19219e-13, 1.19407e-13, 1.195326e-13, 1.196564e-13, 
    1.200306e-13, 1.202287e-13, 1.206719e-13, 1.20592e-13, 1.207274e-13, 
    1.208567e-13, 1.210737e-13, 1.21038e-13, 1.211335e-13, 1.207239e-13, 
    1.209961e-13, 1.205465e-13, 1.206695e-13, 1.196897e-13, 1.193163e-13, 
    1.191571e-13, 1.190181e-13, 1.186793e-13, 1.189132e-13, 1.18821e-13, 
    1.190405e-13, 1.191798e-13, 1.191109e-13, 1.195361e-13, 1.193708e-13, 
    1.202405e-13, 1.198661e-13, 1.208416e-13, 1.206084e-13, 1.208975e-13, 
    1.207501e-13, 1.210027e-13, 1.207753e-13, 1.211691e-13, 1.212548e-13, 
    1.211962e-13, 1.214212e-13, 1.207627e-13, 1.210157e-13, 1.19109e-13, 
    1.191202e-13, 1.191726e-13, 1.189423e-13, 1.189282e-13, 1.187172e-13, 
    1.18905e-13, 1.189849e-13, 1.191879e-13, 1.193079e-13, 1.194219e-13, 
    1.196725e-13, 1.199521e-13, 1.20343e-13, 1.206236e-13, 1.208115e-13, 
    1.206963e-13, 1.20798e-13, 1.206843e-13, 1.20631e-13, 1.212227e-13, 
    1.208905e-13, 1.213888e-13, 1.213613e-13, 1.211358e-13, 1.213644e-13, 
    1.191281e-13, 1.190634e-13, 1.188387e-13, 1.190146e-13, 1.186942e-13, 
    1.188735e-13, 1.189766e-13, 1.193742e-13, 1.194616e-13, 1.195425e-13, 
    1.197024e-13, 1.199074e-13, 1.202667e-13, 1.205792e-13, 1.208643e-13, 
    1.208434e-13, 1.208507e-13, 1.209144e-13, 1.207567e-13, 1.209402e-13, 
    1.20971e-13, 1.208905e-13, 1.213576e-13, 1.212242e-13, 1.213607e-13, 
    1.212739e-13, 1.190845e-13, 1.191933e-13, 1.191345e-13, 1.19245e-13, 
    1.191671e-13, 1.195133e-13, 1.196171e-13, 1.201023e-13, 1.199033e-13, 
    1.2022e-13, 1.199355e-13, 1.199859e-13, 1.202302e-13, 1.199509e-13, 
    1.205619e-13, 1.201476e-13, 1.209168e-13, 1.205034e-13, 1.209427e-13, 
    1.20863e-13, 1.20995e-13, 1.211131e-13, 1.212617e-13, 1.215356e-13, 
    1.214722e-13, 1.217012e-13, 1.193555e-13, 1.194965e-13, 1.194842e-13, 
    1.196317e-13, 1.197408e-13, 1.199772e-13, 1.203561e-13, 1.202137e-13, 
    1.204751e-13, 1.205276e-13, 1.201304e-13, 1.203742e-13, 1.195909e-13, 
    1.197175e-13, 1.196422e-13, 1.193666e-13, 1.202464e-13, 1.197951e-13, 
    1.206282e-13, 1.20384e-13, 1.210962e-13, 1.207421e-13, 1.214373e-13, 
    1.217339e-13, 1.220131e-13, 1.223388e-13, 1.195735e-13, 1.194777e-13, 
    1.196493e-13, 1.198864e-13, 1.201065e-13, 1.203989e-13, 1.204288e-13, 
    1.204835e-13, 1.206253e-13, 1.207444e-13, 1.205008e-13, 1.207743e-13, 
    1.197467e-13, 1.202856e-13, 1.194414e-13, 1.196957e-13, 1.198725e-13, 
    1.19795e-13, 1.201974e-13, 1.202922e-13, 1.20677e-13, 1.204782e-13, 
    1.216606e-13, 1.211379e-13, 1.225868e-13, 1.221825e-13, 1.194442e-13, 
    1.195732e-13, 1.200217e-13, 1.198084e-13, 1.204184e-13, 1.205684e-13, 
    1.206903e-13, 1.20846e-13, 1.208629e-13, 1.209551e-13, 1.20804e-13, 
    1.209492e-13, 1.203995e-13, 1.206452e-13, 1.199706e-13, 1.201349e-13, 
    1.200593e-13, 1.199764e-13, 1.202323e-13, 1.205046e-13, 1.205105e-13, 
    1.205977e-13, 1.208433e-13, 1.204209e-13, 1.217278e-13, 1.20921e-13, 
    1.197138e-13, 1.199619e-13, 1.199975e-13, 1.199014e-13, 1.205533e-13, 
    1.203172e-13, 1.209529e-13, 1.207812e-13, 1.210625e-13, 1.209227e-13, 
    1.209022e-13, 1.207226e-13, 1.206108e-13, 1.20328e-13, 1.200979e-13, 
    1.199153e-13, 1.199578e-13, 1.201583e-13, 1.205212e-13, 1.208644e-13, 
    1.207892e-13, 1.210411e-13, 1.203742e-13, 1.206539e-13, 1.205458e-13, 
    1.208277e-13, 1.202099e-13, 1.207357e-13, 1.200753e-13, 1.201333e-13, 
    1.203125e-13, 1.206728e-13, 1.207527e-13, 1.208377e-13, 1.207852e-13, 
    1.205305e-13, 1.204888e-13, 1.203082e-13, 1.202583e-13, 1.201207e-13, 
    1.200067e-13, 1.201108e-13, 1.202201e-13, 1.205306e-13, 1.208102e-13, 
    1.211148e-13, 1.211893e-13, 1.215445e-13, 1.212552e-13, 1.217323e-13, 
    1.213265e-13, 1.220288e-13, 1.207663e-13, 1.213148e-13, 1.203207e-13, 
    1.20428e-13, 1.206217e-13, 1.210661e-13, 1.208264e-13, 1.211067e-13, 
    1.204871e-13, 1.201652e-13, 1.20082e-13, 1.199264e-13, 1.200855e-13, 
    1.200726e-13, 1.202247e-13, 1.201759e-13, 1.205409e-13, 1.203449e-13, 
    1.209016e-13, 1.211045e-13, 1.216772e-13, 1.220277e-13, 1.223844e-13, 
    1.225416e-13, 1.225895e-13, 1.226095e-13 ;

 LITR3C =
  9.698061e-06, 9.698051e-06, 9.698053e-06, 9.698046e-06, 9.698049e-06, 
    9.698045e-06, 9.698059e-06, 9.698051e-06, 9.698057e-06, 9.69806e-06, 
    9.698029e-06, 9.698045e-06, 9.698014e-06, 9.698024e-06, 9.697999e-06, 
    9.698016e-06, 9.697997e-06, 9.698e-06, 9.697988e-06, 9.697992e-06, 
    9.697977e-06, 9.697987e-06, 9.69797e-06, 9.69798e-06, 9.697978e-06, 
    9.697987e-06, 9.698042e-06, 9.698032e-06, 9.698042e-06, 9.698041e-06, 
    9.698042e-06, 9.698049e-06, 9.698054e-06, 9.698062e-06, 9.69806e-06, 
    9.698054e-06, 9.69804e-06, 9.698045e-06, 9.698033e-06, 9.698033e-06, 
    9.69802e-06, 9.698026e-06, 9.698004e-06, 9.69801e-06, 9.697992e-06, 
    9.697997e-06, 9.697992e-06, 9.697993e-06, 9.697992e-06, 9.697998e-06, 
    9.697996e-06, 9.698002e-06, 9.698025e-06, 9.698018e-06, 9.698038e-06, 
    9.698051e-06, 9.698058e-06, 9.698065e-06, 9.698064e-06, 9.698062e-06, 
    9.698054e-06, 9.698047e-06, 9.698041e-06, 9.698038e-06, 9.698034e-06, 
    9.698022e-06, 9.698016e-06, 9.698003e-06, 9.698005e-06, 9.698001e-06, 
    9.697997e-06, 9.69799e-06, 9.697991e-06, 9.697988e-06, 9.698001e-06, 
    9.697993e-06, 9.698007e-06, 9.698003e-06, 9.698032e-06, 9.698044e-06, 
    9.698048e-06, 9.698053e-06, 9.698063e-06, 9.698056e-06, 9.698058e-06, 
    9.698052e-06, 9.698048e-06, 9.69805e-06, 9.698038e-06, 9.698042e-06, 
    9.698016e-06, 9.698027e-06, 9.697997e-06, 9.698005e-06, 9.697996e-06, 
    9.698e-06, 9.697992e-06, 9.697999e-06, 9.697987e-06, 9.697985e-06, 
    9.697987e-06, 9.697979e-06, 9.697999e-06, 9.697992e-06, 9.69805e-06, 
    9.698049e-06, 9.698048e-06, 9.698055e-06, 9.698056e-06, 9.698062e-06, 
    9.698057e-06, 9.698054e-06, 9.698048e-06, 9.698044e-06, 9.69804e-06, 
    9.698033e-06, 9.698025e-06, 9.698013e-06, 9.698004e-06, 9.697998e-06, 
    9.698002e-06, 9.697998e-06, 9.698002e-06, 9.698004e-06, 9.697986e-06, 
    9.697996e-06, 9.697981e-06, 9.697981e-06, 9.697988e-06, 9.697981e-06, 
    9.698049e-06, 9.698051e-06, 9.698058e-06, 9.698053e-06, 9.698063e-06, 
    9.698058e-06, 9.698054e-06, 9.698042e-06, 9.698039e-06, 9.698037e-06, 
    9.698032e-06, 9.698026e-06, 9.698015e-06, 9.698006e-06, 9.697997e-06, 
    9.697997e-06, 9.697997e-06, 9.697995e-06, 9.698e-06, 9.697995e-06, 
    9.697994e-06, 9.697996e-06, 9.697982e-06, 9.697986e-06, 9.697981e-06, 
    9.697984e-06, 9.698051e-06, 9.698048e-06, 9.698049e-06, 9.698046e-06, 
    9.698048e-06, 9.698038e-06, 9.698035e-06, 9.69802e-06, 9.698026e-06, 
    9.698017e-06, 9.698025e-06, 9.698023e-06, 9.698016e-06, 9.698025e-06, 
    9.698006e-06, 9.698018e-06, 9.697995e-06, 9.698007e-06, 9.697994e-06, 
    9.697997e-06, 9.697993e-06, 9.697989e-06, 9.697985e-06, 9.697977e-06, 
    9.697978e-06, 9.697971e-06, 9.698043e-06, 9.698038e-06, 9.698038e-06, 
    9.698034e-06, 9.698031e-06, 9.698024e-06, 9.698012e-06, 9.698017e-06, 
    9.698008e-06, 9.698007e-06, 9.698019e-06, 9.698011e-06, 9.698036e-06, 
    9.698031e-06, 9.698034e-06, 9.698042e-06, 9.698016e-06, 9.698029e-06, 
    9.698004e-06, 9.698011e-06, 9.697989e-06, 9.698e-06, 9.697979e-06, 
    9.69797e-06, 9.697962e-06, 9.697952e-06, 9.698036e-06, 9.698039e-06, 
    9.698034e-06, 9.698027e-06, 9.698019e-06, 9.698011e-06, 9.69801e-06, 
    9.698008e-06, 9.698004e-06, 9.698e-06, 9.698007e-06, 9.697999e-06, 
    9.69803e-06, 9.698014e-06, 9.69804e-06, 9.698032e-06, 9.698027e-06, 
    9.698029e-06, 9.698017e-06, 9.698014e-06, 9.698002e-06, 9.698008e-06, 
    9.697972e-06, 9.697988e-06, 9.697944e-06, 9.697957e-06, 9.69804e-06, 
    9.698036e-06, 9.698022e-06, 9.698028e-06, 9.69801e-06, 9.698006e-06, 
    9.698002e-06, 9.697997e-06, 9.697997e-06, 9.697994e-06, 9.697998e-06, 
    9.697994e-06, 9.698011e-06, 9.698003e-06, 9.698024e-06, 9.698019e-06, 
    9.698021e-06, 9.698024e-06, 9.698016e-06, 9.698007e-06, 9.698007e-06, 
    9.698005e-06, 9.697997e-06, 9.69801e-06, 9.69797e-06, 9.697995e-06, 
    9.698032e-06, 9.698024e-06, 9.698023e-06, 9.698026e-06, 9.698006e-06, 
    9.698013e-06, 9.697994e-06, 9.697999e-06, 9.69799e-06, 9.697995e-06, 
    9.697996e-06, 9.698001e-06, 9.698005e-06, 9.698013e-06, 9.69802e-06, 
    9.698026e-06, 9.698024e-06, 9.698018e-06, 9.698007e-06, 9.697997e-06, 
    9.697999e-06, 9.697991e-06, 9.698011e-06, 9.698003e-06, 9.698007e-06, 
    9.697997e-06, 9.698017e-06, 9.698e-06, 9.69802e-06, 9.698019e-06, 
    9.698014e-06, 9.698002e-06, 9.698e-06, 9.697997e-06, 9.697999e-06, 
    9.698007e-06, 9.698008e-06, 9.698014e-06, 9.698015e-06, 9.698019e-06, 
    9.698023e-06, 9.698019e-06, 9.698017e-06, 9.698007e-06, 9.697998e-06, 
    9.697989e-06, 9.697987e-06, 9.697976e-06, 9.697985e-06, 9.69797e-06, 
    9.697983e-06, 9.697961e-06, 9.697999e-06, 9.697983e-06, 9.698013e-06, 
    9.69801e-06, 9.698004e-06, 9.69799e-06, 9.697997e-06, 9.697989e-06, 
    9.698008e-06, 9.698017e-06, 9.69802e-06, 9.698025e-06, 9.69802e-06, 
    9.698021e-06, 9.698016e-06, 9.698017e-06, 9.698007e-06, 9.698012e-06, 
    9.697996e-06, 9.697989e-06, 9.697972e-06, 9.697961e-06, 9.69795e-06, 
    9.697946e-06, 9.697944e-06, 9.697944e-06 ;

 LITR3C_TO_SOIL2C =
  5.937168e-14, 5.953458e-14, 5.950294e-14, 5.963423e-14, 5.956143e-14, 
    5.964737e-14, 5.940474e-14, 5.954102e-14, 5.945405e-14, 5.938638e-14, 
    5.988872e-14, 5.964009e-14, 6.014692e-14, 5.998854e-14, 6.038622e-14, 
    6.012224e-14, 6.043942e-14, 6.037867e-14, 6.056159e-14, 6.050921e-14, 
    6.074285e-14, 6.058576e-14, 6.086395e-14, 6.070538e-14, 6.073017e-14, 
    6.058057e-14, 5.969021e-14, 5.985777e-14, 5.968026e-14, 5.970417e-14, 
    5.969345e-14, 5.956292e-14, 5.949706e-14, 5.935926e-14, 5.938429e-14, 
    5.948552e-14, 5.971492e-14, 5.963712e-14, 5.983326e-14, 5.982884e-14, 
    6.004694e-14, 5.994863e-14, 6.031493e-14, 6.02109e-14, 6.05114e-14, 
    6.043586e-14, 6.050784e-14, 6.048603e-14, 6.050812e-14, 6.039733e-14, 
    6.044481e-14, 6.03473e-14, 5.996704e-14, 6.007885e-14, 5.974516e-14, 
    5.954417e-14, 5.941071e-14, 5.931591e-14, 5.932932e-14, 5.935485e-14, 
    5.948611e-14, 5.960951e-14, 5.970348e-14, 5.976631e-14, 5.982819e-14, 
    6.001527e-14, 6.011436e-14, 6.033592e-14, 6.029601e-14, 6.036366e-14, 
    6.042835e-14, 6.053683e-14, 6.051899e-14, 6.056675e-14, 6.036191e-14, 
    6.049805e-14, 6.027325e-14, 6.033476e-14, 5.984482e-14, 5.965812e-14, 
    5.957854e-14, 5.950901e-14, 5.933962e-14, 5.94566e-14, 5.941049e-14, 
    5.952022e-14, 5.958989e-14, 5.955544e-14, 5.976802e-14, 5.96854e-14, 
    6.012022e-14, 5.993304e-14, 6.04208e-14, 6.030421e-14, 6.044875e-14, 
    6.037501e-14, 6.050132e-14, 6.038765e-14, 6.058454e-14, 6.062737e-14, 
    6.05981e-14, 6.071056e-14, 6.038134e-14, 6.050782e-14, 5.955447e-14, 
    5.956008e-14, 5.958627e-14, 5.947113e-14, 5.946408e-14, 5.935856e-14, 
    5.945248e-14, 5.949244e-14, 5.959394e-14, 5.965392e-14, 5.971093e-14, 
    5.983624e-14, 5.997605e-14, 6.017146e-14, 6.031176e-14, 6.040574e-14, 
    6.034813e-14, 6.039899e-14, 6.034213e-14, 6.031548e-14, 6.061131e-14, 
    6.044523e-14, 6.069439e-14, 6.068062e-14, 6.056788e-14, 6.068217e-14, 
    5.956403e-14, 5.95317e-14, 5.941935e-14, 5.950728e-14, 5.934707e-14, 
    5.943674e-14, 5.948826e-14, 5.968708e-14, 5.973078e-14, 5.977124e-14, 
    5.985117e-14, 5.995366e-14, 6.013334e-14, 6.028958e-14, 6.043211e-14, 
    6.042168e-14, 6.042535e-14, 6.045716e-14, 6.037833e-14, 6.04701e-14, 
    6.048548e-14, 6.044524e-14, 6.067878e-14, 6.061209e-14, 6.068033e-14, 
    6.063691e-14, 5.954221e-14, 5.959662e-14, 5.956723e-14, 5.962249e-14, 
    5.958354e-14, 5.975664e-14, 5.980852e-14, 6.005111e-14, 5.995164e-14, 
    6.010999e-14, 5.996774e-14, 5.999294e-14, 6.011507e-14, 5.997545e-14, 
    6.028092e-14, 6.007379e-14, 6.04584e-14, 6.025166e-14, 6.047134e-14, 
    6.04315e-14, 6.049748e-14, 6.055653e-14, 6.063083e-14, 6.076778e-14, 
    6.073609e-14, 6.08506e-14, 5.967773e-14, 5.974823e-14, 5.974206e-14, 
    5.981585e-14, 5.987039e-14, 5.998861e-14, 6.017802e-14, 6.010683e-14, 
    6.023755e-14, 6.026378e-14, 6.006519e-14, 6.018711e-14, 5.979543e-14, 
    5.985872e-14, 5.982106e-14, 5.968327e-14, 6.012318e-14, 5.989751e-14, 
    6.031407e-14, 6.019197e-14, 6.05481e-14, 6.037104e-14, 6.071863e-14, 
    6.086692e-14, 6.100656e-14, 6.116939e-14, 5.978674e-14, 5.973884e-14, 
    5.982463e-14, 5.994319e-14, 6.005325e-14, 6.019942e-14, 6.021439e-14, 
    6.024174e-14, 6.031264e-14, 6.03722e-14, 6.025035e-14, 6.038713e-14, 
    5.987332e-14, 6.014278e-14, 5.972069e-14, 5.984783e-14, 5.993623e-14, 
    5.989749e-14, 6.00987e-14, 6.014608e-14, 6.033848e-14, 6.023907e-14, 
    6.08303e-14, 6.056895e-14, 6.129339e-14, 6.109121e-14, 5.972209e-14, 
    5.978659e-14, 6.001085e-14, 5.990419e-14, 6.020919e-14, 6.028418e-14, 
    6.034515e-14, 6.0423e-14, 6.043143e-14, 6.047754e-14, 6.040197e-14, 
    6.047457e-14, 6.019973e-14, 6.03226e-14, 5.998528e-14, 6.006741e-14, 
    6.002965e-14, 5.998818e-14, 6.011612e-14, 6.025227e-14, 6.025523e-14, 
    6.029886e-14, 6.042162e-14, 6.021043e-14, 6.086389e-14, 6.046049e-14, 
    5.98569e-14, 5.998095e-14, 5.999874e-14, 5.995068e-14, 6.027666e-14, 
    6.01586e-14, 6.047642e-14, 6.03906e-14, 6.053122e-14, 6.046135e-14, 
    6.045107e-14, 6.03613e-14, 6.030536e-14, 6.0164e-14, 6.004892e-14, 
    5.995766e-14, 5.997889e-14, 6.007913e-14, 6.02606e-14, 6.043216e-14, 
    6.039459e-14, 6.052054e-14, 6.018708e-14, 6.032695e-14, 6.027289e-14, 
    6.041384e-14, 6.010492e-14, 6.036783e-14, 6.003765e-14, 6.006663e-14, 
    6.015625e-14, 6.033639e-14, 6.037631e-14, 6.041882e-14, 6.03926e-14, 
    6.026522e-14, 6.024437e-14, 6.015409e-14, 6.012913e-14, 6.006032e-14, 
    6.000331e-14, 6.005539e-14, 6.011005e-14, 6.02653e-14, 6.040507e-14, 
    6.055736e-14, 6.059464e-14, 6.077223e-14, 6.062759e-14, 6.086612e-14, 
    6.066322e-14, 6.101438e-14, 6.038314e-14, 6.065737e-14, 6.016035e-14, 
    6.021397e-14, 6.031086e-14, 6.053301e-14, 6.041317e-14, 6.055335e-14, 
    6.024356e-14, 6.008256e-14, 6.004096e-14, 5.99632e-14, 6.004274e-14, 
    6.003627e-14, 6.011236e-14, 6.008791e-14, 6.027045e-14, 6.017242e-14, 
    6.045079e-14, 6.055226e-14, 6.083858e-14, 6.101384e-14, 6.119216e-14, 
    6.12708e-14, 6.129473e-14, 6.130473e-14 ;

 LITR3C_vr =
  0.0005537693, 0.0005537688, 0.0005537689, 0.0005537684, 0.0005537687, 
    0.0005537684, 0.0005537692, 0.0005537687, 0.0005537691, 0.0005537693, 
    0.0005537675, 0.0005537684, 0.0005537666, 0.0005537672, 0.0005537658, 
    0.0005537667, 0.0005537656, 0.0005537658, 0.0005537652, 0.0005537653, 
    0.0005537646, 0.0005537651, 0.0005537641, 0.0005537647, 0.0005537646, 
    0.0005537651, 0.0005537682, 0.0005537676, 0.0005537682, 0.0005537682, 
    0.0005537682, 0.0005537687, 0.0005537689, 0.0005537694, 0.0005537693, 
    0.0005537689, 0.0005537681, 0.0005537684, 0.0005537677, 0.0005537677, 
    0.000553767, 0.0005537673, 0.000553766, 0.0005537664, 0.0005537653, 
    0.0005537656, 0.0005537654, 0.0005537655, 0.0005537654, 0.0005537657, 
    0.0005537656, 0.0005537659, 0.0005537673, 0.0005537668, 0.000553768, 
    0.0005537687, 0.0005537692, 0.0005537695, 0.0005537695, 0.0005537694, 
    0.0005537689, 0.0005537685, 0.0005537682, 0.000553768, 0.0005537677, 
    0.0005537671, 0.0005537667, 0.000553766, 0.0005537661, 0.0005537659, 
    0.0005537656, 0.0005537653, 0.0005537653, 0.0005537652, 0.0005537659, 
    0.0005537654, 0.0005537662, 0.000553766, 0.0005537677, 0.0005537683, 
    0.0005537686, 0.0005537688, 0.0005537694, 0.000553769, 0.0005537692, 
    0.0005537688, 0.0005537685, 0.0005537687, 0.000553768, 0.0005537682, 
    0.0005537667, 0.0005537674, 0.0005537657, 0.0005537661, 0.0005537656, 
    0.0005537658, 0.0005537654, 0.0005537658, 0.0005537651, 0.0005537649, 
    0.000553765, 0.0005537646, 0.0005537658, 0.0005537654, 0.0005537687, 
    0.0005537687, 0.0005537686, 0.0005537689, 0.000553769, 0.0005537694, 
    0.0005537691, 0.0005537689, 0.0005537685, 0.0005537684, 0.0005537681, 
    0.0005537677, 0.0005537672, 0.0005537666, 0.000553766, 0.0005537657, 
    0.0005537659, 0.0005537657, 0.0005537659, 0.000553766, 0.000553765, 
    0.0005537656, 0.0005537647, 0.0005537648, 0.0005537652, 0.0005537648, 
    0.0005537687, 0.0005537688, 0.0005537692, 0.0005537688, 0.0005537694, 
    0.0005537691, 0.0005537689, 0.0005537682, 0.0005537681, 0.000553768, 
    0.0005537677, 0.0005537673, 0.0005537667, 0.0005537661, 0.0005537656, 
    0.0005537657, 0.0005537656, 0.0005537656, 0.0005537658, 0.0005537655, 
    0.0005537655, 0.0005537656, 0.0005537648, 0.000553765, 0.0005537648, 
    0.0005537649, 0.0005537687, 0.0005537685, 0.0005537687, 0.0005537684, 
    0.0005537686, 0.000553768, 0.0005537678, 0.000553767, 0.0005537673, 
    0.0005537667, 0.0005537673, 0.0005537671, 0.0005537667, 0.0005537672, 
    0.0005537661, 0.0005537668, 0.0005537656, 0.0005537663, 0.0005537655, 
    0.0005537656, 0.0005537654, 0.0005537652, 0.0005537649, 0.0005537645, 
    0.0005537646, 0.0005537642, 0.0005537682, 0.000553768, 0.000553768, 
    0.0005537678, 0.0005537676, 0.0005537672, 0.0005537665, 0.0005537668, 
    0.0005537663, 0.0005537662, 0.0005537669, 0.0005537665, 0.0005537678, 
    0.0005537676, 0.0005537678, 0.0005537682, 0.0005537667, 0.0005537675, 
    0.000553766, 0.0005537664, 0.0005537652, 0.0005537659, 0.0005537646, 
    0.0005537641, 0.0005537636, 0.0005537631, 0.0005537679, 0.000553768, 
    0.0005537677, 0.0005537673, 0.000553767, 0.0005537664, 0.0005537664, 
    0.0005537663, 0.000553766, 0.0005537659, 0.0005537663, 0.0005537658, 
    0.0005537675, 0.0005537666, 0.0005537681, 0.0005537677, 0.0005537674, 
    0.0005537675, 0.0005537668, 0.0005537666, 0.000553766, 0.0005537663, 
    0.0005537642, 0.0005537652, 0.0005537627, 0.0005537634, 0.0005537681, 
    0.0005537679, 0.0005537671, 0.0005537675, 0.0005537664, 0.0005537661, 
    0.0005537659, 0.0005537657, 0.0005537656, 0.0005537655, 0.0005537657, 
    0.0005537655, 0.0005537664, 0.000553766, 0.0005537672, 0.0005537669, 
    0.000553767, 0.0005537672, 0.0005537667, 0.0005537663, 0.0005537663, 
    0.0005537661, 0.0005537657, 0.0005537664, 0.0005537641, 0.0005537655, 
    0.0005537676, 0.0005537672, 0.0005537671, 0.0005537673, 0.0005537661, 
    0.0005537666, 0.0005537655, 0.0005537658, 0.0005537653, 0.0005537655, 
    0.0005537656, 0.0005537659, 0.0005537661, 0.0005537666, 0.000553767, 
    0.0005537673, 0.0005537672, 0.0005537668, 0.0005537662, 0.0005537656, 
    0.0005537657, 0.0005537653, 0.0005537665, 0.000553766, 0.0005537662, 
    0.0005537657, 0.0005537668, 0.0005537659, 0.000553767, 0.0005537669, 
    0.0005537666, 0.000553766, 0.0005537658, 0.0005537657, 0.0005537657, 
    0.0005537662, 0.0005537663, 0.0005537666, 0.0005537667, 0.0005537669, 
    0.0005537671, 0.000553767, 0.0005537667, 0.0005537662, 0.0005537657, 
    0.0005537652, 0.000553765, 0.0005537645, 0.0005537649, 0.0005537641, 
    0.0005537648, 0.0005537636, 0.0005537658, 0.0005537649, 0.0005537666, 
    0.0005537664, 0.000553766, 0.0005537653, 0.0005537657, 0.0005537652, 
    0.0005537663, 0.0005537668, 0.000553767, 0.0005537673, 0.000553767, 
    0.000553767, 0.0005537667, 0.0005537668, 0.0005537662, 0.0005537666, 
    0.0005537656, 0.0005537652, 0.0005537642, 0.0005537636, 0.000553763, 
    0.0005537627, 0.0005537627, 0.0005537626,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342141e-07, 1.342139e-07, 1.34214e-07, 1.342138e-07, 1.342139e-07, 
    1.342138e-07, 1.34214e-07, 1.342139e-07, 1.34214e-07, 1.342141e-07, 
    1.342136e-07, 1.342138e-07, 1.342134e-07, 1.342136e-07, 1.342132e-07, 
    1.342134e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.342129e-07, 1.342131e-07, 1.342128e-07, 1.34213e-07, 1.342129e-07, 
    1.342131e-07, 1.342138e-07, 1.342137e-07, 1.342138e-07, 1.342138e-07, 
    1.342138e-07, 1.342139e-07, 1.34214e-07, 1.342141e-07, 1.342141e-07, 
    1.34214e-07, 1.342138e-07, 1.342138e-07, 1.342137e-07, 1.342137e-07, 
    1.342135e-07, 1.342136e-07, 1.342133e-07, 1.342134e-07, 1.342131e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342133e-07, 1.342136e-07, 1.342135e-07, 1.342138e-07, 
    1.342139e-07, 1.34214e-07, 1.342141e-07, 1.342141e-07, 1.342141e-07, 
    1.34214e-07, 1.342139e-07, 1.342138e-07, 1.342137e-07, 1.342137e-07, 
    1.342135e-07, 1.342135e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342133e-07, 1.342133e-07, 1.342137e-07, 1.342138e-07, 
    1.342139e-07, 1.34214e-07, 1.342141e-07, 1.34214e-07, 1.34214e-07, 
    1.342139e-07, 1.342139e-07, 1.342139e-07, 1.342137e-07, 1.342138e-07, 
    1.342134e-07, 1.342136e-07, 1.342132e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 1.342139e-07, 
    1.342139e-07, 1.342139e-07, 1.34214e-07, 1.34214e-07, 1.342141e-07, 
    1.34214e-07, 1.34214e-07, 1.342139e-07, 1.342138e-07, 1.342138e-07, 
    1.342137e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342133e-07, 1.342132e-07, 1.342133e-07, 1.342133e-07, 1.34213e-07, 
    1.342132e-07, 1.34213e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 
    1.342139e-07, 1.342139e-07, 1.34214e-07, 1.34214e-07, 1.342141e-07, 
    1.34214e-07, 1.34214e-07, 1.342138e-07, 1.342138e-07, 1.342137e-07, 
    1.342137e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342132e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342139e-07, 1.342139e-07, 1.342139e-07, 1.342139e-07, 
    1.342139e-07, 1.342137e-07, 1.342137e-07, 1.342135e-07, 1.342136e-07, 
    1.342135e-07, 1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342136e-07, 
    1.342133e-07, 1.342135e-07, 1.342132e-07, 1.342133e-07, 1.342131e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342138e-07, 1.342137e-07, 1.342138e-07, 
    1.342137e-07, 1.342136e-07, 1.342136e-07, 1.342134e-07, 1.342135e-07, 
    1.342133e-07, 1.342133e-07, 1.342135e-07, 1.342134e-07, 1.342137e-07, 
    1.342137e-07, 1.342137e-07, 1.342138e-07, 1.342134e-07, 1.342136e-07, 
    1.342133e-07, 1.342134e-07, 1.342131e-07, 1.342132e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342137e-07, 1.342138e-07, 
    1.342137e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342132e-07, 1.342133e-07, 1.342132e-07, 
    1.342136e-07, 1.342134e-07, 1.342138e-07, 1.342137e-07, 1.342136e-07, 
    1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342128e-07, 1.342131e-07, 1.342125e-07, 1.342126e-07, 1.342138e-07, 
    1.342137e-07, 1.342135e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342134e-07, 1.342133e-07, 1.342136e-07, 1.342135e-07, 
    1.342135e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.342134e-07, 1.342128e-07, 1.342132e-07, 
    1.342137e-07, 1.342136e-07, 1.342135e-07, 1.342136e-07, 1.342133e-07, 
    1.342134e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342132e-07, 1.342133e-07, 1.342134e-07, 1.342135e-07, 
    1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342132e-07, 1.342135e-07, 1.342132e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342135e-07, 1.342133e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 
    1.34213e-07, 1.342127e-07, 1.342132e-07, 1.34213e-07, 1.342134e-07, 
    1.342134e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 
    1.342133e-07, 1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342135e-07, 1.342133e-07, 1.342134e-07, 
    1.342132e-07, 1.342131e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342124e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  5.024356e-26, -1.838179e-26, -1.102908e-26, 2.450905e-26, 4.901811e-26, 
    6.372354e-26, 8.210533e-26, 1.470543e-26, 8.455624e-26, 4.41163e-26, 
    7.352717e-27, 1.519561e-25, 3.798904e-26, -4.901811e-26, -7.965443e-26, 
    -4.166539e-26, -1.960724e-26, -1.225453e-26, 7.352717e-27, -8.578169e-27, 
    -1.225453e-27, 5.391992e-26, -8.333079e-26, -9.803622e-27, -8.700715e-26, 
    4.166539e-26, 3.431268e-26, 9.803622e-27, 5.024356e-26, -1.151926e-25, 
    -6.249809e-26, 8.087988e-26, 1.347998e-26, -1.347998e-26, 2.205815e-26, 
    5.391992e-26, 9.803622e-26, -2.695996e-26, 1.960724e-26, 9.926167e-26, 
    5.637083e-26, -7.230172e-26, -8.578169e-26, -4.289085e-26, -6.249809e-26, 
    -7.352717e-26, 6.98508e-26, -4.779266e-26, -5.391992e-26, 4.534175e-26, 
    -9.803622e-26, 4.65672e-26, 6.004719e-26, -6.127264e-27, -2.818541e-26, 
    -8.700715e-26, 1.372507e-25, -1.470543e-26, -4.901811e-26, -2.205815e-26, 
    -2.941087e-26, 4.901811e-27, -5.882173e-26, -8.578169e-26, -7.352717e-27, 
    8.578169e-27, 3.553813e-26, -8.578169e-27, 1.213198e-25, 2.695996e-26, 
    6.004719e-26, 5.391992e-26, -1.151926e-25, -5.269447e-26, -6.4949e-26, 
    4.901811e-27, 5.024356e-26, 1.470543e-26, 1.470543e-26, 7.652491e-42, 
    -2.32836e-26, 2.450906e-27, -7.107626e-26, 6.4949e-26, 8.700715e-26, 
    -4.901811e-26, 3.431268e-26, 8.578169e-27, -9.190896e-26, 0, 
    -2.695996e-26, 7.352717e-26, -6.862535e-26, 2.695996e-26, -3.826946e-42, 
    -6.862535e-26, -1.225453e-26, 6.73999e-26, 4.043994e-26, 7.597807e-26, 
    5.514538e-26, 1.470543e-25, -4.534175e-26, -2.573451e-26, 5.391992e-26, 
    4.166539e-26, 7.720352e-26, -6.372354e-26, -6.862535e-26, 9.926167e-26, 
    -3.798904e-26, -5.024356e-26, -1.593089e-26, 5.514538e-26, -3.676358e-27, 
    -5.759628e-26, 3.676358e-27, 6.004719e-26, 2.941087e-26, -3.798904e-26, 
    5.882173e-26, -2.205815e-26, 1.102908e-25, 1.274471e-25, 6.862535e-26, 
    -1.041635e-25, -8.210533e-26, -2.695996e-26, -4.779266e-26, 2.450906e-27, 
    -4.166539e-26, 6.617445e-26, -2.941087e-26, -6.004719e-26, -3.431268e-26, 
    2.818541e-26, -3.186177e-26, -1.323489e-25, -1.605343e-25, 6.127264e-27, 
    1.531816e-25, -1.960724e-26, 3.186177e-26, 4.901811e-27, -6.127264e-26, 
    5.146902e-26, -2.450906e-27, -3.676358e-26, 1.225453e-26, 2.08327e-26, 
    -1.041635e-25, 1.470543e-26, 1.715634e-26, -1.347998e-26, -8.945805e-26, 
    8.945805e-26, 1.593089e-26, 2.205815e-26, -5.882173e-26, 1.102908e-26, 
    8.700715e-26, 4.166539e-26, 2.08327e-26, 1.102908e-26, 5.146902e-26, 
    -6.127264e-26, 6.127264e-26, 8.333079e-26, -7.720352e-26, -9.068351e-26, 
    -6.617445e-26, -5.391992e-26, -3.431268e-26, -4.65672e-26, 3.921449e-26, 
    1.017126e-25, -6.004719e-26, 2.818541e-26, -5.269447e-26, 2.32836e-26, 
    7.107626e-26, 4.779266e-26, 8.578169e-26, -5.514538e-26, 9.313441e-26, 
    1.200944e-25, -4.41163e-26, 6.127264e-26, 3.553813e-26, 3.798904e-26, 
    1.115162e-25, -1.715634e-26, -3.186177e-26, -6.862535e-26, 2.32836e-26, 
    -4.901811e-27, 8.578169e-26, 2.941087e-26, 1.200944e-25, -1.360253e-25, 
    -1.102908e-26, -4.534175e-26, 1.115162e-25, -2.695996e-26, 2.08327e-26, 
    -5.514538e-26, -6.127264e-26, -3.676358e-26, -1.213198e-25, 
    -7.107626e-26, 3.186177e-26, 1.470543e-25, 3.063632e-26, -1.593089e-26, 
    3.676358e-26, -1.115162e-25, 5.882173e-26, -1.347998e-25, -1.470543e-25, 
    5.024356e-26, -9.803622e-26, 1.715634e-26, 9.803622e-27, -4.043994e-26, 
    7.352717e-27, -4.289085e-26, 1.16418e-25, 7.965443e-26, 5.882173e-26, 
    -4.901811e-26, -1.225453e-26, 4.779266e-26, -1.715634e-26, 6.249809e-26, 
    -1.02938e-25, 1.102908e-26, -4.41163e-26, 1.347998e-26, 3.921449e-26, 
    -1.593089e-26, 1.347998e-26, 1.200944e-25, -6.617445e-26, 1.078398e-25, 
    -1.715634e-26, -1.470543e-26, 6.127264e-26, 1.593089e-26, -6.004719e-26, 
    6.004719e-26, -6.127264e-27, -6.862535e-26, -2.08327e-26, -4.289085e-26, 
    -2.08327e-26, -6.617445e-26, 1.225453e-27, 8.578169e-27, -4.901811e-26, 
    8.578169e-27, -2.573451e-26, -2.32836e-26, -2.818541e-26, -2.450905e-26, 
    1.017126e-25, -1.715634e-26, -4.901811e-26, 3.186177e-26, 3.798904e-26, 
    5.759628e-26, 5.146902e-26, 3.063632e-26, -8.210533e-26, -2.695996e-26, 
    -4.901811e-26, 7.842898e-26, 1.188689e-25, 3.063632e-26, -2.32836e-26, 
    1.43378e-25, -6.249809e-26, 1.225453e-27, 6.127264e-26, -5.759628e-26, 
    5.514538e-26, 4.043994e-26, -6.249809e-26, 1.960724e-26, 6.862535e-26, 
    -8.455624e-26, -9.803622e-27, -4.289085e-26, 8.82326e-26, 2.32836e-26, 
    1.347998e-26, 8.087988e-26, 3.553813e-26, 1.090653e-25, 1.127417e-25, 
    -9.068351e-26, -5.514538e-26, -6.862535e-26, 4.901811e-26, 1.960724e-26, 
    4.901811e-26, 4.65672e-26, 2.573451e-26, 2.450905e-26, -5.024356e-26, 
    4.41163e-26, -4.901811e-26, -8.087988e-26, 3.798904e-26, -3.676358e-27, 
    -1.323489e-25, -7.597807e-26, -8.578169e-26, 2.450906e-27, -4.901811e-26, 
    -4.289085e-26, -7.352717e-27, 7.842898e-26, -5.391992e-26, -8.210533e-26, 
    1.225453e-27, -1.225453e-27, 3.798904e-26, -5.882173e-26, -3.921449e-26, 
    1.225453e-26, -1.176435e-25, 8.578169e-26, -9.681077e-26, -1.225453e-27, 
    -5.146902e-26, -9.681077e-26, -1.642107e-25, 1.225453e-25,
  1.338134e-32, 1.338133e-32, 1.338133e-32, 1.338132e-32, 1.338132e-32, 
    1.338131e-32, 1.338134e-32, 1.338132e-32, 1.338133e-32, 1.338134e-32, 
    1.338129e-32, 1.338132e-32, 1.338127e-32, 1.338129e-32, 1.338125e-32, 
    1.338128e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338122e-32, 1.338124e-32, 1.338121e-32, 1.338123e-32, 1.338122e-32, 
    1.338124e-32, 1.338131e-32, 1.33813e-32, 1.338131e-32, 1.338131e-32, 
    1.338131e-32, 1.338132e-32, 1.338133e-32, 1.338134e-32, 1.338134e-32, 
    1.338133e-32, 1.338131e-32, 1.338132e-32, 1.33813e-32, 1.33813e-32, 
    1.338128e-32, 1.338129e-32, 1.338126e-32, 1.338127e-32, 1.338124e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338126e-32, 1.338129e-32, 1.338128e-32, 1.338131e-32, 
    1.338132e-32, 1.338134e-32, 1.338134e-32, 1.338134e-32, 1.338134e-32, 
    1.338133e-32, 1.338132e-32, 1.338131e-32, 1.33813e-32, 1.33813e-32, 
    1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338126e-32, 1.338126e-32, 1.33813e-32, 1.338131e-32, 
    1.338132e-32, 1.338133e-32, 1.338134e-32, 1.338133e-32, 1.338134e-32, 
    1.338133e-32, 1.338132e-32, 1.338132e-32, 1.33813e-32, 1.338131e-32, 
    1.338128e-32, 1.338129e-32, 1.338125e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338123e-32, 
    1.338123e-32, 1.338123e-32, 1.338125e-32, 1.338124e-32, 1.338132e-32, 
    1.338132e-32, 1.338132e-32, 1.338133e-32, 1.338133e-32, 1.338134e-32, 
    1.338133e-32, 1.338133e-32, 1.338132e-32, 1.338131e-32, 1.338131e-32, 
    1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338126e-32, 1.338125e-32, 1.338126e-32, 1.338126e-32, 1.338123e-32, 
    1.338125e-32, 1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 
    1.338132e-32, 1.338133e-32, 1.338133e-32, 1.338133e-32, 1.338134e-32, 
    1.338133e-32, 1.338133e-32, 1.338131e-32, 1.338131e-32, 1.33813e-32, 
    1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338125e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338132e-32, 1.338132e-32, 1.338132e-32, 1.338132e-32, 
    1.338132e-32, 1.338131e-32, 1.33813e-32, 1.338128e-32, 1.338129e-32, 
    1.338128e-32, 1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338129e-32, 
    1.338126e-32, 1.338128e-32, 1.338125e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338131e-32, 1.338131e-32, 1.338131e-32, 
    1.33813e-32, 1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338128e-32, 
    1.338126e-32, 1.338126e-32, 1.338128e-32, 1.338127e-32, 1.33813e-32, 
    1.33813e-32, 1.33813e-32, 1.338131e-32, 1.338128e-32, 1.338129e-32, 
    1.338126e-32, 1.338127e-32, 1.338124e-32, 1.338125e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.33813e-32, 1.338131e-32, 
    1.33813e-32, 1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338127e-32, 
    1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338126e-32, 1.338125e-32, 
    1.33813e-32, 1.338127e-32, 1.338131e-32, 1.33813e-32, 1.338129e-32, 
    1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338121e-32, 1.338124e-32, 1.338118e-32, 1.338119e-32, 1.338131e-32, 
    1.33813e-32, 1.338128e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338127e-32, 1.338126e-32, 1.338129e-32, 1.338128e-32, 
    1.338128e-32, 1.338129e-32, 1.338128e-32, 1.338126e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338127e-32, 1.338121e-32, 1.338125e-32, 
    1.33813e-32, 1.338129e-32, 1.338129e-32, 1.338129e-32, 1.338126e-32, 
    1.338127e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338126e-32, 1.338127e-32, 1.338128e-32, 
    1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338125e-32, 1.338128e-32, 1.338125e-32, 1.338128e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 1.338128e-32, 
    1.338129e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338123e-32, 1.338121e-32, 
    1.338123e-32, 1.33812e-32, 1.338125e-32, 1.338123e-32, 1.338127e-32, 
    1.338127e-32, 1.338126e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 
    1.338126e-32, 1.338128e-32, 1.338128e-32, 1.338129e-32, 1.338128e-32, 
    1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338127e-32, 
    1.338125e-32, 1.338124e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338118e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.643321e-15, 1.64783e-15, 1.646954e-15, 1.650588e-15, 1.648573e-15, 
    1.650952e-15, 1.644236e-15, 1.648008e-15, 1.645601e-15, 1.643728e-15, 
    1.657632e-15, 1.650751e-15, 1.664779e-15, 1.660395e-15, 1.671402e-15, 
    1.664096e-15, 1.672875e-15, 1.671193e-15, 1.676256e-15, 1.674806e-15, 
    1.681273e-15, 1.676925e-15, 1.684625e-15, 1.680236e-15, 1.680922e-15, 
    1.676781e-15, 1.652138e-15, 1.656775e-15, 1.651862e-15, 1.652524e-15, 
    1.652228e-15, 1.648614e-15, 1.646792e-15, 1.642977e-15, 1.64367e-15, 
    1.646472e-15, 1.652822e-15, 1.650668e-15, 1.656097e-15, 1.655975e-15, 
    1.662012e-15, 1.65929e-15, 1.669429e-15, 1.66655e-15, 1.674867e-15, 
    1.672776e-15, 1.674768e-15, 1.674165e-15, 1.674776e-15, 1.67171e-15, 
    1.673024e-15, 1.670325e-15, 1.6598e-15, 1.662895e-15, 1.653659e-15, 
    1.648095e-15, 1.644401e-15, 1.641778e-15, 1.642149e-15, 1.642856e-15, 
    1.646489e-15, 1.649904e-15, 1.652505e-15, 1.654244e-15, 1.655957e-15, 
    1.661135e-15, 1.663877e-15, 1.67001e-15, 1.668905e-15, 1.670778e-15, 
    1.672568e-15, 1.675571e-15, 1.675077e-15, 1.676399e-15, 1.67073e-15, 
    1.674498e-15, 1.668275e-15, 1.669978e-15, 1.656417e-15, 1.651249e-15, 
    1.649047e-15, 1.647122e-15, 1.642434e-15, 1.645672e-15, 1.644395e-15, 
    1.647433e-15, 1.649361e-15, 1.648408e-15, 1.654291e-15, 1.652004e-15, 
    1.66404e-15, 1.658859e-15, 1.672359e-15, 1.669132e-15, 1.673133e-15, 
    1.671092e-15, 1.674588e-15, 1.671442e-15, 1.676891e-15, 1.678077e-15, 
    1.677267e-15, 1.68038e-15, 1.671267e-15, 1.674768e-15, 1.648381e-15, 
    1.648536e-15, 1.649261e-15, 1.646074e-15, 1.645879e-15, 1.642958e-15, 
    1.645558e-15, 1.646664e-15, 1.649473e-15, 1.651133e-15, 1.652711e-15, 
    1.656179e-15, 1.660049e-15, 1.665458e-15, 1.669341e-15, 1.671943e-15, 
    1.670348e-15, 1.671756e-15, 1.670182e-15, 1.669444e-15, 1.677632e-15, 
    1.673036e-15, 1.679932e-15, 1.679551e-15, 1.67643e-15, 1.679594e-15, 
    1.648645e-15, 1.64775e-15, 1.644641e-15, 1.647074e-15, 1.64264e-15, 
    1.645122e-15, 1.646548e-15, 1.652051e-15, 1.653261e-15, 1.65438e-15, 
    1.656593e-15, 1.65943e-15, 1.664403e-15, 1.668727e-15, 1.672673e-15, 
    1.672384e-15, 1.672485e-15, 1.673366e-15, 1.671184e-15, 1.673724e-15, 
    1.67415e-15, 1.673036e-15, 1.6795e-15, 1.677654e-15, 1.679543e-15, 
    1.678341e-15, 1.648042e-15, 1.649547e-15, 1.648734e-15, 1.650263e-15, 
    1.649185e-15, 1.653976e-15, 1.655412e-15, 1.662127e-15, 1.659374e-15, 
    1.663757e-15, 1.659819e-15, 1.660517e-15, 1.663897e-15, 1.660033e-15, 
    1.668488e-15, 1.662755e-15, 1.6734e-15, 1.667678e-15, 1.673758e-15, 
    1.672656e-15, 1.674482e-15, 1.676116e-15, 1.678173e-15, 1.681963e-15, 
    1.681086e-15, 1.684256e-15, 1.651792e-15, 1.653744e-15, 1.653573e-15, 
    1.655615e-15, 1.657125e-15, 1.660397e-15, 1.66564e-15, 1.663669e-15, 
    1.667287e-15, 1.668013e-15, 1.662516e-15, 1.665891e-15, 1.65505e-15, 
    1.656802e-15, 1.65576e-15, 1.651945e-15, 1.664122e-15, 1.657875e-15, 
    1.669405e-15, 1.666026e-15, 1.675883e-15, 1.670982e-15, 1.680603e-15, 
    1.684707e-15, 1.688572e-15, 1.693079e-15, 1.654809e-15, 1.653484e-15, 
    1.655858e-15, 1.65914e-15, 1.662186e-15, 1.666232e-15, 1.666646e-15, 
    1.667403e-15, 1.669365e-15, 1.671014e-15, 1.667642e-15, 1.671427e-15, 
    1.657206e-15, 1.664664e-15, 1.652981e-15, 1.6565e-15, 1.658947e-15, 
    1.657875e-15, 1.663444e-15, 1.664755e-15, 1.670081e-15, 1.667329e-15, 
    1.683694e-15, 1.67646e-15, 1.696511e-15, 1.690915e-15, 1.65302e-15, 
    1.654805e-15, 1.661013e-15, 1.65806e-15, 1.666502e-15, 1.668578e-15, 
    1.670265e-15, 1.67242e-15, 1.672654e-15, 1.67393e-15, 1.671838e-15, 
    1.673848e-15, 1.66624e-15, 1.669641e-15, 1.660305e-15, 1.662578e-15, 
    1.661533e-15, 1.660385e-15, 1.663926e-15, 1.667694e-15, 1.667777e-15, 
    1.668984e-15, 1.672382e-15, 1.666536e-15, 1.684623e-15, 1.673458e-15, 
    1.656751e-15, 1.660185e-15, 1.660677e-15, 1.659347e-15, 1.66837e-15, 
    1.665102e-15, 1.673899e-15, 1.671523e-15, 1.675416e-15, 1.673482e-15, 
    1.673197e-15, 1.670712e-15, 1.669164e-15, 1.665252e-15, 1.662066e-15, 
    1.65954e-15, 1.660128e-15, 1.662902e-15, 1.667925e-15, 1.672674e-15, 
    1.671634e-15, 1.67512e-15, 1.665891e-15, 1.669762e-15, 1.668265e-15, 
    1.672167e-15, 1.663616e-15, 1.670893e-15, 1.661754e-15, 1.662556e-15, 
    1.665037e-15, 1.670023e-15, 1.671128e-15, 1.672305e-15, 1.671579e-15, 
    1.668053e-15, 1.667476e-15, 1.664977e-15, 1.664286e-15, 1.662382e-15, 
    1.660804e-15, 1.662245e-15, 1.663758e-15, 1.668055e-15, 1.671924e-15, 
    1.676139e-15, 1.677171e-15, 1.682086e-15, 1.678083e-15, 1.684685e-15, 
    1.679069e-15, 1.688789e-15, 1.671317e-15, 1.678907e-15, 1.665151e-15, 
    1.666635e-15, 1.669316e-15, 1.675465e-15, 1.672148e-15, 1.676028e-15, 
    1.667453e-15, 1.662997e-15, 1.661846e-15, 1.659694e-15, 1.661895e-15, 
    1.661716e-15, 1.663822e-15, 1.663145e-15, 1.668198e-15, 1.665485e-15, 
    1.673189e-15, 1.675998e-15, 1.683923e-15, 1.688774e-15, 1.69371e-15, 
    1.695886e-15, 1.696548e-15, 1.696825e-15 ;

 LITR3N_vr =
  7.663763e-06, 7.663754e-06, 7.663756e-06, 7.66375e-06, 7.663753e-06, 
    7.663749e-06, 7.663761e-06, 7.663754e-06, 7.663758e-06, 7.663762e-06, 
    7.663737e-06, 7.663749e-06, 7.663725e-06, 7.663733e-06, 7.663713e-06, 
    7.663726e-06, 7.663711e-06, 7.663713e-06, 7.663705e-06, 7.663707e-06, 
    7.663696e-06, 7.663703e-06, 7.663691e-06, 7.663698e-06, 7.663697e-06, 
    7.663704e-06, 7.663747e-06, 7.663739e-06, 7.663747e-06, 7.663746e-06, 
    7.663747e-06, 7.663753e-06, 7.663756e-06, 7.663763e-06, 7.663762e-06, 
    7.663757e-06, 7.663745e-06, 7.66375e-06, 7.66374e-06, 7.66374e-06, 
    7.66373e-06, 7.663734e-06, 7.663717e-06, 7.663722e-06, 7.663707e-06, 
    7.663711e-06, 7.663707e-06, 7.663709e-06, 7.663707e-06, 7.663712e-06, 
    7.663711e-06, 7.663715e-06, 7.663733e-06, 7.663728e-06, 7.663744e-06, 
    7.663754e-06, 7.663761e-06, 7.663765e-06, 7.663764e-06, 7.663763e-06, 
    7.663757e-06, 7.663751e-06, 7.663746e-06, 7.663743e-06, 7.66374e-06, 
    7.663732e-06, 7.663726e-06, 7.663716e-06, 7.663718e-06, 7.663714e-06, 
    7.663712e-06, 7.663706e-06, 7.663707e-06, 7.663704e-06, 7.663714e-06, 
    7.663708e-06, 7.663719e-06, 7.663716e-06, 7.66374e-06, 7.663748e-06, 
    7.663753e-06, 7.663755e-06, 7.663763e-06, 7.663758e-06, 7.663761e-06, 
    7.663755e-06, 7.663752e-06, 7.663753e-06, 7.663743e-06, 7.663747e-06, 
    7.663726e-06, 7.663735e-06, 7.663712e-06, 7.663717e-06, 7.663711e-06, 
    7.663714e-06, 7.663708e-06, 7.663713e-06, 7.663703e-06, 7.663702e-06, 
    7.663703e-06, 7.663698e-06, 7.663713e-06, 7.663707e-06, 7.663753e-06, 
    7.663753e-06, 7.663752e-06, 7.663757e-06, 7.663758e-06, 7.663763e-06, 
    7.663758e-06, 7.663756e-06, 7.663752e-06, 7.663749e-06, 7.663746e-06, 
    7.66374e-06, 7.663733e-06, 7.663723e-06, 7.663717e-06, 7.663712e-06, 
    7.663715e-06, 7.663712e-06, 7.663715e-06, 7.663717e-06, 7.663702e-06, 
    7.663711e-06, 7.663699e-06, 7.663699e-06, 7.663704e-06, 7.663699e-06, 
    7.663753e-06, 7.663754e-06, 7.66376e-06, 7.663755e-06, 7.663763e-06, 
    7.663759e-06, 7.663756e-06, 7.663747e-06, 7.663745e-06, 7.663743e-06, 
    7.663739e-06, 7.663734e-06, 7.663725e-06, 7.663718e-06, 7.663711e-06, 
    7.663712e-06, 7.663712e-06, 7.66371e-06, 7.663713e-06, 7.663709e-06, 
    7.663709e-06, 7.663711e-06, 7.663699e-06, 7.663702e-06, 7.663699e-06, 
    7.663702e-06, 7.663754e-06, 7.663752e-06, 7.663753e-06, 7.66375e-06, 
    7.663752e-06, 7.663743e-06, 7.663742e-06, 7.66373e-06, 7.663734e-06, 
    7.663727e-06, 7.663733e-06, 7.663733e-06, 7.663726e-06, 7.663733e-06, 
    7.663718e-06, 7.663728e-06, 7.66371e-06, 7.66372e-06, 7.663709e-06, 
    7.663712e-06, 7.663708e-06, 7.663705e-06, 7.663702e-06, 7.663695e-06, 
    7.663696e-06, 7.663691e-06, 7.663747e-06, 7.663744e-06, 7.663744e-06, 
    7.663741e-06, 7.663738e-06, 7.663733e-06, 7.663723e-06, 7.663727e-06, 
    7.663721e-06, 7.663719e-06, 7.663729e-06, 7.663722e-06, 7.663742e-06, 
    7.663739e-06, 7.663741e-06, 7.663747e-06, 7.663726e-06, 7.663737e-06, 
    7.663717e-06, 7.663722e-06, 7.663705e-06, 7.663714e-06, 7.663697e-06, 
    7.66369e-06, 7.663683e-06, 7.663675e-06, 7.663743e-06, 7.663744e-06, 
    7.663741e-06, 7.663734e-06, 7.66373e-06, 7.663722e-06, 7.663722e-06, 
    7.663721e-06, 7.663717e-06, 7.663714e-06, 7.66372e-06, 7.663713e-06, 
    7.663738e-06, 7.663725e-06, 7.663745e-06, 7.663739e-06, 7.663735e-06, 
    7.663737e-06, 7.663727e-06, 7.663725e-06, 7.663715e-06, 7.663721e-06, 
    7.663692e-06, 7.663704e-06, 7.66367e-06, 7.66368e-06, 7.663745e-06, 
    7.663743e-06, 7.663732e-06, 7.663736e-06, 7.663722e-06, 7.663718e-06, 
    7.663715e-06, 7.663712e-06, 7.663712e-06, 7.663709e-06, 7.663712e-06, 
    7.663709e-06, 7.663722e-06, 7.663716e-06, 7.663733e-06, 7.663729e-06, 
    7.663731e-06, 7.663733e-06, 7.663726e-06, 7.66372e-06, 7.66372e-06, 
    7.663718e-06, 7.663712e-06, 7.663722e-06, 7.663691e-06, 7.66371e-06, 
    7.663739e-06, 7.663733e-06, 7.663732e-06, 7.663734e-06, 7.663719e-06, 
    7.663724e-06, 7.663709e-06, 7.663713e-06, 7.663706e-06, 7.66371e-06, 
    7.66371e-06, 7.663714e-06, 7.663717e-06, 7.663724e-06, 7.66373e-06, 
    7.663734e-06, 7.663733e-06, 7.663728e-06, 7.66372e-06, 7.663711e-06, 
    7.663712e-06, 7.663707e-06, 7.663722e-06, 7.663716e-06, 7.663719e-06, 
    7.663712e-06, 7.663727e-06, 7.663714e-06, 7.66373e-06, 7.663729e-06, 
    7.663724e-06, 7.663716e-06, 7.663713e-06, 7.663712e-06, 7.663713e-06, 
    7.663719e-06, 7.66372e-06, 7.663724e-06, 7.663726e-06, 7.663729e-06, 
    7.663732e-06, 7.663729e-06, 7.663727e-06, 7.663719e-06, 7.663712e-06, 
    7.663705e-06, 7.663703e-06, 7.663694e-06, 7.663702e-06, 7.66369e-06, 
    7.6637e-06, 7.663683e-06, 7.663713e-06, 7.663701e-06, 7.663724e-06, 
    7.663722e-06, 7.663717e-06, 7.663706e-06, 7.663712e-06, 7.663705e-06, 
    7.66372e-06, 7.663728e-06, 7.66373e-06, 7.663733e-06, 7.66373e-06, 
    7.66373e-06, 7.663726e-06, 7.663728e-06, 7.663719e-06, 7.663723e-06, 
    7.66371e-06, 7.663705e-06, 7.663692e-06, 7.663683e-06, 7.663674e-06, 
    7.663671e-06, 7.66367e-06, 7.663669e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.937168e-14, 5.953458e-14, 5.950294e-14, 5.963423e-14, 5.956143e-14, 
    5.964737e-14, 5.940474e-14, 5.954102e-14, 5.945405e-14, 5.938638e-14, 
    5.988872e-14, 5.964009e-14, 6.014692e-14, 5.998854e-14, 6.038622e-14, 
    6.012224e-14, 6.043942e-14, 6.037867e-14, 6.056159e-14, 6.050921e-14, 
    6.074285e-14, 6.058576e-14, 6.086395e-14, 6.070538e-14, 6.073017e-14, 
    6.058057e-14, 5.969021e-14, 5.985777e-14, 5.968026e-14, 5.970417e-14, 
    5.969345e-14, 5.956292e-14, 5.949706e-14, 5.935926e-14, 5.938429e-14, 
    5.948552e-14, 5.971492e-14, 5.963712e-14, 5.983326e-14, 5.982884e-14, 
    6.004694e-14, 5.994863e-14, 6.031493e-14, 6.02109e-14, 6.05114e-14, 
    6.043586e-14, 6.050784e-14, 6.048603e-14, 6.050812e-14, 6.039733e-14, 
    6.044481e-14, 6.03473e-14, 5.996704e-14, 6.007885e-14, 5.974516e-14, 
    5.954417e-14, 5.941071e-14, 5.931591e-14, 5.932932e-14, 5.935485e-14, 
    5.948611e-14, 5.960951e-14, 5.970348e-14, 5.976631e-14, 5.982819e-14, 
    6.001527e-14, 6.011436e-14, 6.033592e-14, 6.029601e-14, 6.036366e-14, 
    6.042835e-14, 6.053683e-14, 6.051899e-14, 6.056675e-14, 6.036191e-14, 
    6.049805e-14, 6.027325e-14, 6.033476e-14, 5.984482e-14, 5.965812e-14, 
    5.957854e-14, 5.950901e-14, 5.933962e-14, 5.94566e-14, 5.941049e-14, 
    5.952022e-14, 5.958989e-14, 5.955544e-14, 5.976802e-14, 5.96854e-14, 
    6.012022e-14, 5.993304e-14, 6.04208e-14, 6.030421e-14, 6.044875e-14, 
    6.037501e-14, 6.050132e-14, 6.038765e-14, 6.058454e-14, 6.062737e-14, 
    6.05981e-14, 6.071056e-14, 6.038134e-14, 6.050782e-14, 5.955447e-14, 
    5.956008e-14, 5.958627e-14, 5.947113e-14, 5.946408e-14, 5.935856e-14, 
    5.945248e-14, 5.949244e-14, 5.959394e-14, 5.965392e-14, 5.971093e-14, 
    5.983624e-14, 5.997605e-14, 6.017146e-14, 6.031176e-14, 6.040574e-14, 
    6.034813e-14, 6.039899e-14, 6.034213e-14, 6.031548e-14, 6.061131e-14, 
    6.044523e-14, 6.069439e-14, 6.068062e-14, 6.056788e-14, 6.068217e-14, 
    5.956403e-14, 5.95317e-14, 5.941935e-14, 5.950728e-14, 5.934707e-14, 
    5.943674e-14, 5.948826e-14, 5.968708e-14, 5.973078e-14, 5.977124e-14, 
    5.985117e-14, 5.995366e-14, 6.013334e-14, 6.028958e-14, 6.043211e-14, 
    6.042168e-14, 6.042535e-14, 6.045716e-14, 6.037833e-14, 6.04701e-14, 
    6.048548e-14, 6.044524e-14, 6.067878e-14, 6.061209e-14, 6.068033e-14, 
    6.063691e-14, 5.954221e-14, 5.959662e-14, 5.956723e-14, 5.962249e-14, 
    5.958354e-14, 5.975664e-14, 5.980852e-14, 6.005111e-14, 5.995164e-14, 
    6.010999e-14, 5.996774e-14, 5.999294e-14, 6.011507e-14, 5.997545e-14, 
    6.028092e-14, 6.007379e-14, 6.04584e-14, 6.025166e-14, 6.047134e-14, 
    6.04315e-14, 6.049748e-14, 6.055653e-14, 6.063083e-14, 6.076778e-14, 
    6.073609e-14, 6.08506e-14, 5.967773e-14, 5.974823e-14, 5.974206e-14, 
    5.981585e-14, 5.987039e-14, 5.998861e-14, 6.017802e-14, 6.010683e-14, 
    6.023755e-14, 6.026378e-14, 6.006519e-14, 6.018711e-14, 5.979543e-14, 
    5.985872e-14, 5.982106e-14, 5.968327e-14, 6.012318e-14, 5.989751e-14, 
    6.031407e-14, 6.019197e-14, 6.05481e-14, 6.037104e-14, 6.071863e-14, 
    6.086692e-14, 6.100656e-14, 6.116939e-14, 5.978674e-14, 5.973884e-14, 
    5.982463e-14, 5.994319e-14, 6.005325e-14, 6.019942e-14, 6.021439e-14, 
    6.024174e-14, 6.031264e-14, 6.03722e-14, 6.025035e-14, 6.038713e-14, 
    5.987332e-14, 6.014278e-14, 5.972069e-14, 5.984783e-14, 5.993623e-14, 
    5.989749e-14, 6.00987e-14, 6.014608e-14, 6.033848e-14, 6.023907e-14, 
    6.08303e-14, 6.056895e-14, 6.129339e-14, 6.109121e-14, 5.972209e-14, 
    5.978659e-14, 6.001085e-14, 5.990419e-14, 6.020919e-14, 6.028418e-14, 
    6.034515e-14, 6.0423e-14, 6.043143e-14, 6.047754e-14, 6.040197e-14, 
    6.047457e-14, 6.019973e-14, 6.03226e-14, 5.998528e-14, 6.006741e-14, 
    6.002965e-14, 5.998818e-14, 6.011612e-14, 6.025227e-14, 6.025523e-14, 
    6.029886e-14, 6.042162e-14, 6.021043e-14, 6.086389e-14, 6.046049e-14, 
    5.98569e-14, 5.998095e-14, 5.999874e-14, 5.995068e-14, 6.027666e-14, 
    6.01586e-14, 6.047642e-14, 6.03906e-14, 6.053122e-14, 6.046135e-14, 
    6.045107e-14, 6.03613e-14, 6.030536e-14, 6.0164e-14, 6.004892e-14, 
    5.995766e-14, 5.997889e-14, 6.007913e-14, 6.02606e-14, 6.043216e-14, 
    6.039459e-14, 6.052054e-14, 6.018708e-14, 6.032695e-14, 6.027289e-14, 
    6.041384e-14, 6.010492e-14, 6.036783e-14, 6.003765e-14, 6.006663e-14, 
    6.015625e-14, 6.033639e-14, 6.037631e-14, 6.041882e-14, 6.03926e-14, 
    6.026522e-14, 6.024437e-14, 6.015409e-14, 6.012913e-14, 6.006032e-14, 
    6.000331e-14, 6.005539e-14, 6.011005e-14, 6.02653e-14, 6.040507e-14, 
    6.055736e-14, 6.059464e-14, 6.077223e-14, 6.062759e-14, 6.086612e-14, 
    6.066322e-14, 6.101438e-14, 6.038314e-14, 6.065737e-14, 6.016035e-14, 
    6.021397e-14, 6.031086e-14, 6.053301e-14, 6.041317e-14, 6.055335e-14, 
    6.024356e-14, 6.008256e-14, 6.004096e-14, 5.99632e-14, 6.004274e-14, 
    6.003627e-14, 6.011236e-14, 6.008791e-14, 6.027045e-14, 6.017242e-14, 
    6.045079e-14, 6.055226e-14, 6.083858e-14, 6.101384e-14, 6.119216e-14, 
    6.12708e-14, 6.129473e-14, 6.130473e-14 ;

 LITTERC =
  5.976299e-05, 5.976284e-05, 5.976287e-05, 5.976275e-05, 5.976282e-05, 
    5.976274e-05, 5.976296e-05, 5.976284e-05, 5.976292e-05, 5.976298e-05, 
    5.976252e-05, 5.976275e-05, 5.976229e-05, 5.976243e-05, 5.976207e-05, 
    5.976231e-05, 5.976202e-05, 5.976207e-05, 5.976191e-05, 5.976195e-05, 
    5.976174e-05, 5.976189e-05, 5.976163e-05, 5.976178e-05, 5.976175e-05, 
    5.976189e-05, 5.97627e-05, 5.976255e-05, 5.976271e-05, 5.976269e-05, 
    5.97627e-05, 5.976282e-05, 5.976288e-05, 5.9763e-05, 5.976298e-05, 
    5.976289e-05, 5.976268e-05, 5.976275e-05, 5.976257e-05, 5.976257e-05, 
    5.976238e-05, 5.976246e-05, 5.976213e-05, 5.976223e-05, 5.976195e-05, 
    5.976202e-05, 5.976195e-05, 5.976198e-05, 5.976195e-05, 5.976206e-05, 
    5.976201e-05, 5.97621e-05, 5.976245e-05, 5.976235e-05, 5.976265e-05, 
    5.976284e-05, 5.976296e-05, 5.976304e-05, 5.976303e-05, 5.976301e-05, 
    5.976289e-05, 5.976277e-05, 5.976269e-05, 5.976263e-05, 5.976258e-05, 
    5.976241e-05, 5.976231e-05, 5.976211e-05, 5.976215e-05, 5.976209e-05, 
    5.976203e-05, 5.976193e-05, 5.976195e-05, 5.97619e-05, 5.976209e-05, 
    5.976197e-05, 5.976217e-05, 5.976211e-05, 5.976256e-05, 5.976273e-05, 
    5.97628e-05, 5.976286e-05, 5.976302e-05, 5.976291e-05, 5.976296e-05, 
    5.976286e-05, 5.976279e-05, 5.976282e-05, 5.976263e-05, 5.97627e-05, 
    5.976231e-05, 5.976248e-05, 5.976203e-05, 5.976214e-05, 5.976201e-05, 
    5.976208e-05, 5.976196e-05, 5.976207e-05, 5.976189e-05, 5.976185e-05, 
    5.976187e-05, 5.976177e-05, 5.976207e-05, 5.976195e-05, 5.976282e-05, 
    5.976282e-05, 5.976279e-05, 5.97629e-05, 5.976291e-05, 5.9763e-05, 
    5.976292e-05, 5.976288e-05, 5.976279e-05, 5.976273e-05, 5.976268e-05, 
    5.976257e-05, 5.976244e-05, 5.976226e-05, 5.976214e-05, 5.976205e-05, 
    5.97621e-05, 5.976206e-05, 5.976211e-05, 5.976213e-05, 5.976186e-05, 
    5.976201e-05, 5.976179e-05, 5.97618e-05, 5.97619e-05, 5.97618e-05, 
    5.976282e-05, 5.976285e-05, 5.976295e-05, 5.976287e-05, 5.976301e-05, 
    5.976293e-05, 5.976289e-05, 5.97627e-05, 5.976266e-05, 5.976263e-05, 
    5.976255e-05, 5.976246e-05, 5.97623e-05, 5.976215e-05, 5.976202e-05, 
    5.976203e-05, 5.976203e-05, 5.9762e-05, 5.976207e-05, 5.976199e-05, 
    5.976198e-05, 5.976201e-05, 5.97618e-05, 5.976186e-05, 5.97618e-05, 
    5.976184e-05, 5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976276e-05, 
    5.97628e-05, 5.976264e-05, 5.976259e-05, 5.976237e-05, 5.976246e-05, 
    5.976232e-05, 5.976245e-05, 5.976242e-05, 5.976231e-05, 5.976244e-05, 
    5.976216e-05, 5.976235e-05, 5.9762e-05, 5.976219e-05, 5.976199e-05, 
    5.976203e-05, 5.976197e-05, 5.976191e-05, 5.976185e-05, 5.976172e-05, 
    5.976175e-05, 5.976165e-05, 5.976271e-05, 5.976265e-05, 5.976265e-05, 
    5.976259e-05, 5.976254e-05, 5.976243e-05, 5.976226e-05, 5.976232e-05, 
    5.97622e-05, 5.976218e-05, 5.976236e-05, 5.976225e-05, 5.976261e-05, 
    5.976255e-05, 5.976258e-05, 5.976271e-05, 5.976231e-05, 5.976251e-05, 
    5.976213e-05, 5.976224e-05, 5.976192e-05, 5.976208e-05, 5.976177e-05, 
    5.976163e-05, 5.97615e-05, 5.976135e-05, 5.976261e-05, 5.976266e-05, 
    5.976258e-05, 5.976247e-05, 5.976237e-05, 5.976224e-05, 5.976222e-05, 
    5.97622e-05, 5.976213e-05, 5.976208e-05, 5.976219e-05, 5.976207e-05, 
    5.976253e-05, 5.976229e-05, 5.976267e-05, 5.976256e-05, 5.976247e-05, 
    5.976251e-05, 5.976233e-05, 5.976229e-05, 5.976211e-05, 5.97622e-05, 
    5.976166e-05, 5.97619e-05, 5.976124e-05, 5.976142e-05, 5.976267e-05, 
    5.976261e-05, 5.976241e-05, 5.97625e-05, 5.976223e-05, 5.976216e-05, 
    5.97621e-05, 5.976203e-05, 5.976203e-05, 5.976198e-05, 5.976205e-05, 
    5.976199e-05, 5.976224e-05, 5.976213e-05, 5.976243e-05, 5.976236e-05, 
    5.976239e-05, 5.976243e-05, 5.976231e-05, 5.976219e-05, 5.976219e-05, 
    5.976215e-05, 5.976203e-05, 5.976223e-05, 5.976163e-05, 5.9762e-05, 
    5.976255e-05, 5.976243e-05, 5.976242e-05, 5.976246e-05, 5.976217e-05, 
    5.976227e-05, 5.976198e-05, 5.976206e-05, 5.976194e-05, 5.9762e-05, 
    5.976201e-05, 5.976209e-05, 5.976214e-05, 5.976227e-05, 5.976237e-05, 
    5.976246e-05, 5.976244e-05, 5.976235e-05, 5.976218e-05, 5.976202e-05, 
    5.976206e-05, 5.976194e-05, 5.976225e-05, 5.976212e-05, 5.976217e-05, 
    5.976204e-05, 5.976232e-05, 5.976208e-05, 5.976238e-05, 5.976236e-05, 
    5.976227e-05, 5.976211e-05, 5.976207e-05, 5.976204e-05, 5.976206e-05, 
    5.976218e-05, 5.976219e-05, 5.976228e-05, 5.97623e-05, 5.976236e-05, 
    5.976242e-05, 5.976237e-05, 5.976232e-05, 5.976218e-05, 5.976205e-05, 
    5.976191e-05, 5.976188e-05, 5.976171e-05, 5.976185e-05, 5.976163e-05, 
    5.976182e-05, 5.97615e-05, 5.976207e-05, 5.976182e-05, 5.976227e-05, 
    5.976222e-05, 5.976214e-05, 5.976193e-05, 5.976204e-05, 5.976191e-05, 
    5.97622e-05, 5.976234e-05, 5.976238e-05, 5.976245e-05, 5.976238e-05, 
    5.976238e-05, 5.976231e-05, 5.976234e-05, 5.976217e-05, 5.976226e-05, 
    5.976201e-05, 5.976191e-05, 5.976166e-05, 5.97615e-05, 5.976133e-05, 
    5.976126e-05, 5.976124e-05, 5.976123e-05 ;

 LITTERC_HR =
  9.578916e-13, 9.605178e-13, 9.600076e-13, 9.621242e-13, 9.609506e-13, 
    9.62336e-13, 9.584246e-13, 9.606217e-13, 9.592195e-13, 9.581287e-13, 
    9.662267e-13, 9.622187e-13, 9.703888e-13, 9.678357e-13, 9.742465e-13, 
    9.699911e-13, 9.75104e-13, 9.741248e-13, 9.770735e-13, 9.762291e-13, 
    9.799954e-13, 9.774631e-13, 9.819474e-13, 9.793914e-13, 9.797909e-13, 
    9.773793e-13, 9.630265e-13, 9.657276e-13, 9.628662e-13, 9.632516e-13, 
    9.630789e-13, 9.609745e-13, 9.599129e-13, 9.576915e-13, 9.58095e-13, 
    9.59727e-13, 9.634249e-13, 9.621707e-13, 9.653326e-13, 9.652612e-13, 
    9.687773e-13, 9.671925e-13, 9.730971e-13, 9.714202e-13, 9.762643e-13, 
    9.750466e-13, 9.76207e-13, 9.758552e-13, 9.762115e-13, 9.744256e-13, 
    9.751908e-13, 9.736191e-13, 9.674891e-13, 9.692916e-13, 9.639123e-13, 
    9.606722e-13, 9.585208e-13, 9.569927e-13, 9.572087e-13, 9.576205e-13, 
    9.597364e-13, 9.617256e-13, 9.632404e-13, 9.642532e-13, 9.65251e-13, 
    9.682667e-13, 9.698639e-13, 9.734356e-13, 9.727922e-13, 9.738828e-13, 
    9.749255e-13, 9.766743e-13, 9.763866e-13, 9.771566e-13, 9.738547e-13, 
    9.760492e-13, 9.724254e-13, 9.734169e-13, 9.655189e-13, 9.625093e-13, 
    9.612264e-13, 9.601056e-13, 9.573748e-13, 9.592607e-13, 9.585173e-13, 
    9.602862e-13, 9.614093e-13, 9.608541e-13, 9.64281e-13, 9.629489e-13, 
    9.699585e-13, 9.669412e-13, 9.748039e-13, 9.729243e-13, 9.752544e-13, 
    9.740658e-13, 9.761018e-13, 9.742695e-13, 9.774434e-13, 9.781337e-13, 
    9.77662e-13, 9.79475e-13, 9.741678e-13, 9.762066e-13, 9.608384e-13, 
    9.609289e-13, 9.613511e-13, 9.594947e-13, 9.593813e-13, 9.576802e-13, 
    9.591942e-13, 9.598384e-13, 9.614747e-13, 9.624416e-13, 9.633607e-13, 
    9.653806e-13, 9.676344e-13, 9.707844e-13, 9.730462e-13, 9.745611e-13, 
    9.736325e-13, 9.744523e-13, 9.735357e-13, 9.731061e-13, 9.778749e-13, 
    9.751978e-13, 9.792142e-13, 9.789923e-13, 9.771748e-13, 9.790172e-13, 
    9.609926e-13, 9.604713e-13, 9.586601e-13, 9.600776e-13, 9.574949e-13, 
    9.589405e-13, 9.597711e-13, 9.629761e-13, 9.636806e-13, 9.643328e-13, 
    9.656211e-13, 9.672736e-13, 9.7017e-13, 9.726885e-13, 9.749864e-13, 
    9.748181e-13, 9.748773e-13, 9.7539e-13, 9.741193e-13, 9.755986e-13, 
    9.758466e-13, 9.751979e-13, 9.789625e-13, 9.778875e-13, 9.789875e-13, 
    9.782877e-13, 9.606409e-13, 9.615179e-13, 9.61044e-13, 9.61935e-13, 
    9.61307e-13, 9.640975e-13, 9.649336e-13, 9.688445e-13, 9.672408e-13, 
    9.697936e-13, 9.675005e-13, 9.679067e-13, 9.698754e-13, 9.676246e-13, 
    9.725491e-13, 9.692101e-13, 9.7541e-13, 9.720773e-13, 9.756186e-13, 
    9.749764e-13, 9.7604e-13, 9.769918e-13, 9.781895e-13, 9.803973e-13, 
    9.798863e-13, 9.817323e-13, 9.628253e-13, 9.639619e-13, 9.638625e-13, 
    9.650518e-13, 9.659311e-13, 9.678368e-13, 9.708903e-13, 9.697426e-13, 
    9.7185e-13, 9.722726e-13, 9.690713e-13, 9.710366e-13, 9.647228e-13, 
    9.65743e-13, 9.651361e-13, 9.629146e-13, 9.700063e-13, 9.663684e-13, 
    9.730834e-13, 9.711151e-13, 9.768561e-13, 9.740017e-13, 9.79605e-13, 
    9.819954e-13, 9.842463e-13, 9.868711e-13, 9.645827e-13, 9.638105e-13, 
    9.651934e-13, 9.671048e-13, 9.688789e-13, 9.712351e-13, 9.714765e-13, 
    9.719174e-13, 9.730602e-13, 9.740205e-13, 9.720563e-13, 9.742611e-13, 
    9.659784e-13, 9.703221e-13, 9.63518e-13, 9.655675e-13, 9.669924e-13, 
    9.66368e-13, 9.696115e-13, 9.703754e-13, 9.734769e-13, 9.718743e-13, 
    9.814051e-13, 9.771921e-13, 9.8887e-13, 9.85611e-13, 9.635406e-13, 
    9.645803e-13, 9.681955e-13, 9.664759e-13, 9.713927e-13, 9.726014e-13, 
    9.735844e-13, 9.748393e-13, 9.749752e-13, 9.757185e-13, 9.745003e-13, 
    9.756707e-13, 9.712401e-13, 9.73221e-13, 9.677831e-13, 9.691072e-13, 
    9.684984e-13, 9.6783e-13, 9.698924e-13, 9.720871e-13, 9.721349e-13, 
    9.728381e-13, 9.748172e-13, 9.714126e-13, 9.819465e-13, 9.754437e-13, 
    9.657136e-13, 9.677134e-13, 9.680001e-13, 9.672254e-13, 9.724803e-13, 
    9.705771e-13, 9.757006e-13, 9.74317e-13, 9.765839e-13, 9.754576e-13, 
    9.752918e-13, 9.738446e-13, 9.729431e-13, 9.706642e-13, 9.688092e-13, 
    9.67338e-13, 9.676801e-13, 9.692961e-13, 9.722214e-13, 9.749871e-13, 
    9.743814e-13, 9.764118e-13, 9.710364e-13, 9.73291e-13, 9.724195e-13, 
    9.746917e-13, 9.697119e-13, 9.7395e-13, 9.686273e-13, 9.690946e-13, 
    9.705394e-13, 9.734432e-13, 9.740868e-13, 9.74772e-13, 9.743494e-13, 
    9.722959e-13, 9.719598e-13, 9.705045e-13, 9.70102e-13, 9.689929e-13, 
    9.680739e-13, 9.689133e-13, 9.697944e-13, 9.722971e-13, 9.745503e-13, 
    9.770053e-13, 9.776061e-13, 9.80469e-13, 9.781374e-13, 9.819825e-13, 
    9.787117e-13, 9.843724e-13, 9.741969e-13, 9.786174e-13, 9.706054e-13, 
    9.714698e-13, 9.730316e-13, 9.766128e-13, 9.746809e-13, 9.769405e-13, 
    9.719467e-13, 9.693514e-13, 9.686808e-13, 9.674272e-13, 9.687095e-13, 
    9.686052e-13, 9.698316e-13, 9.694376e-13, 9.723803e-13, 9.707999e-13, 
    9.752873e-13, 9.76923e-13, 9.815385e-13, 9.843636e-13, 9.872382e-13, 
    9.885058e-13, 9.888916e-13, 9.890528e-13 ;

 LITTERC_LOSS =
  1.774006e-12, 1.778869e-12, 1.777925e-12, 1.781844e-12, 1.779671e-12, 
    1.782237e-12, 1.774993e-12, 1.779062e-12, 1.776465e-12, 1.774445e-12, 
    1.789442e-12, 1.782019e-12, 1.797151e-12, 1.792422e-12, 1.804295e-12, 
    1.796414e-12, 1.805883e-12, 1.80407e-12, 1.809531e-12, 1.807967e-12, 
    1.814942e-12, 1.810252e-12, 1.818557e-12, 1.813824e-12, 1.814564e-12, 
    1.810097e-12, 1.783516e-12, 1.788518e-12, 1.783219e-12, 1.783932e-12, 
    1.783613e-12, 1.779715e-12, 1.777749e-12, 1.773635e-12, 1.774382e-12, 
    1.777405e-12, 1.784253e-12, 1.781931e-12, 1.787786e-12, 1.787654e-12, 
    1.794166e-12, 1.791231e-12, 1.802167e-12, 1.799061e-12, 1.808032e-12, 
    1.805777e-12, 1.807926e-12, 1.807275e-12, 1.807934e-12, 1.804627e-12, 
    1.806044e-12, 1.803133e-12, 1.79178e-12, 1.795119e-12, 1.785156e-12, 
    1.779155e-12, 1.775171e-12, 1.772341e-12, 1.772741e-12, 1.773503e-12, 
    1.777422e-12, 1.781106e-12, 1.783912e-12, 1.785787e-12, 1.787635e-12, 
    1.793221e-12, 1.796179e-12, 1.802793e-12, 1.801602e-12, 1.803622e-12, 
    1.805553e-12, 1.808792e-12, 1.808259e-12, 1.809685e-12, 1.803569e-12, 
    1.807634e-12, 1.800922e-12, 1.802759e-12, 1.788132e-12, 1.782558e-12, 
    1.780182e-12, 1.778106e-12, 1.773049e-12, 1.776541e-12, 1.775164e-12, 
    1.778441e-12, 1.780521e-12, 1.779492e-12, 1.785839e-12, 1.783372e-12, 
    1.796354e-12, 1.790766e-12, 1.805328e-12, 1.801847e-12, 1.806162e-12, 
    1.803961e-12, 1.807731e-12, 1.804338e-12, 1.810216e-12, 1.811494e-12, 
    1.810621e-12, 1.813978e-12, 1.804149e-12, 1.807925e-12, 1.779463e-12, 
    1.779631e-12, 1.780413e-12, 1.776975e-12, 1.776765e-12, 1.773614e-12, 
    1.776418e-12, 1.777611e-12, 1.780642e-12, 1.782432e-12, 1.784134e-12, 
    1.787875e-12, 1.79205e-12, 1.797883e-12, 1.802072e-12, 1.804878e-12, 
    1.803158e-12, 1.804676e-12, 1.802979e-12, 1.802183e-12, 1.811015e-12, 
    1.806057e-12, 1.813496e-12, 1.813084e-12, 1.809718e-12, 1.813131e-12, 
    1.779749e-12, 1.778783e-12, 1.775429e-12, 1.778054e-12, 1.773271e-12, 
    1.775948e-12, 1.777486e-12, 1.783422e-12, 1.784727e-12, 1.785935e-12, 
    1.788321e-12, 1.791381e-12, 1.796745e-12, 1.80141e-12, 1.805665e-12, 
    1.805354e-12, 1.805463e-12, 1.806413e-12, 1.80406e-12, 1.806799e-12, 
    1.807259e-12, 1.806057e-12, 1.813029e-12, 1.811038e-12, 1.813076e-12, 
    1.81178e-12, 1.779097e-12, 1.780722e-12, 1.779844e-12, 1.781494e-12, 
    1.780331e-12, 1.785499e-12, 1.787048e-12, 1.794291e-12, 1.791321e-12, 
    1.796048e-12, 1.791802e-12, 1.792554e-12, 1.7962e-12, 1.792031e-12, 
    1.801152e-12, 1.794968e-12, 1.80645e-12, 1.800278e-12, 1.806836e-12, 
    1.805647e-12, 1.807617e-12, 1.80938e-12, 1.811598e-12, 1.815687e-12, 
    1.81474e-12, 1.818159e-12, 1.783143e-12, 1.785248e-12, 1.785064e-12, 
    1.787267e-12, 1.788895e-12, 1.792424e-12, 1.798079e-12, 1.795954e-12, 
    1.799857e-12, 1.80064e-12, 1.794711e-12, 1.798351e-12, 1.786657e-12, 
    1.788547e-12, 1.787423e-12, 1.783308e-12, 1.796442e-12, 1.789705e-12, 
    1.802141e-12, 1.798496e-12, 1.809128e-12, 1.803842e-12, 1.814219e-12, 
    1.818646e-12, 1.822815e-12, 1.827676e-12, 1.786398e-12, 1.784968e-12, 
    1.787529e-12, 1.791069e-12, 1.794354e-12, 1.798718e-12, 1.799165e-12, 
    1.799982e-12, 1.802098e-12, 1.803876e-12, 1.800239e-12, 1.804322e-12, 
    1.788983e-12, 1.797027e-12, 1.784426e-12, 1.788222e-12, 1.790861e-12, 
    1.789704e-12, 1.795711e-12, 1.797126e-12, 1.80287e-12, 1.799902e-12, 
    1.817553e-12, 1.80975e-12, 1.831378e-12, 1.825342e-12, 1.784468e-12, 
    1.786393e-12, 1.793089e-12, 1.789904e-12, 1.79901e-12, 1.801249e-12, 
    1.803069e-12, 1.805393e-12, 1.805645e-12, 1.807022e-12, 1.804765e-12, 
    1.806933e-12, 1.798727e-12, 1.802396e-12, 1.792325e-12, 1.794777e-12, 
    1.79365e-12, 1.792412e-12, 1.796231e-12, 1.800296e-12, 1.800384e-12, 
    1.801687e-12, 1.805352e-12, 1.799047e-12, 1.818556e-12, 1.806512e-12, 
    1.788492e-12, 1.792196e-12, 1.792727e-12, 1.791292e-12, 1.801024e-12, 
    1.7975e-12, 1.806988e-12, 1.804426e-12, 1.808624e-12, 1.806538e-12, 
    1.806231e-12, 1.803551e-12, 1.801881e-12, 1.797661e-12, 1.794225e-12, 
    1.7915e-12, 1.792134e-12, 1.795127e-12, 1.800545e-12, 1.805667e-12, 
    1.804545e-12, 1.808305e-12, 1.79835e-12, 1.802526e-12, 1.800912e-12, 
    1.80512e-12, 1.795897e-12, 1.803746e-12, 1.793888e-12, 1.794754e-12, 
    1.79743e-12, 1.802807e-12, 1.803999e-12, 1.805268e-12, 1.804486e-12, 
    1.800683e-12, 1.80006e-12, 1.797365e-12, 1.79662e-12, 1.794565e-12, 
    1.792863e-12, 1.794418e-12, 1.79605e-12, 1.800685e-12, 1.804858e-12, 
    1.809405e-12, 1.810517e-12, 1.815819e-12, 1.811501e-12, 1.818623e-12, 
    1.812565e-12, 1.823048e-12, 1.804203e-12, 1.81239e-12, 1.797552e-12, 
    1.799153e-12, 1.802045e-12, 1.808678e-12, 1.8051e-12, 1.809285e-12, 
    1.800036e-12, 1.795229e-12, 1.793987e-12, 1.791666e-12, 1.794041e-12, 
    1.793847e-12, 1.796119e-12, 1.795389e-12, 1.800839e-12, 1.797912e-12, 
    1.806223e-12, 1.809252e-12, 1.8178e-12, 1.823032e-12, 1.828356e-12, 
    1.830704e-12, 1.831418e-12, 1.831717e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.676203e-18, 1.676465e-18, 1.676415e-18, 1.676624e-18, 1.67651e-18, 
    1.676646e-18, 1.676258e-18, 1.676474e-18, 1.676337e-18, 1.67623e-18, 
    1.677024e-18, 1.676634e-18, 1.677452e-18, 1.677199e-18, 1.677842e-18, 
    1.67741e-18, 1.67793e-18, 1.677835e-18, 1.678135e-18, 1.67805e-18, 
    1.678424e-18, 1.678175e-18, 1.678627e-18, 1.678367e-18, 1.678406e-18, 
    1.678166e-18, 1.676718e-18, 1.676974e-18, 1.676701e-18, 1.676738e-18, 
    1.676723e-18, 1.676511e-18, 1.676401e-18, 1.676186e-18, 1.676226e-18, 
    1.676386e-18, 1.676755e-18, 1.676633e-18, 1.676951e-18, 1.676944e-18, 
    1.677294e-18, 1.677136e-18, 1.677731e-18, 1.677563e-18, 1.678053e-18, 
    1.677929e-18, 1.678047e-18, 1.678012e-18, 1.678047e-18, 1.677865e-18, 
    1.677943e-18, 1.677784e-18, 1.677165e-18, 1.677345e-18, 1.676805e-18, 
    1.676474e-18, 1.676267e-18, 1.676116e-18, 1.676137e-18, 1.676177e-18, 
    1.676387e-18, 1.676588e-18, 1.676741e-18, 1.676842e-18, 1.676942e-18, 
    1.677234e-18, 1.677399e-18, 1.677762e-18, 1.677701e-18, 1.677808e-18, 
    1.677917e-18, 1.678093e-18, 1.678065e-18, 1.678142e-18, 1.677808e-18, 
    1.678028e-18, 1.677665e-18, 1.677764e-18, 1.676952e-18, 1.676667e-18, 
    1.67653e-18, 1.676424e-18, 1.676153e-18, 1.67634e-18, 1.676266e-18, 
    1.676445e-18, 1.676556e-18, 1.676502e-18, 1.676845e-18, 1.676711e-18, 
    1.677409e-18, 1.677108e-18, 1.677904e-18, 1.677714e-18, 1.67795e-18, 
    1.677831e-18, 1.678035e-18, 1.677851e-18, 1.678172e-18, 1.67824e-18, 
    1.678193e-18, 1.678379e-18, 1.67784e-18, 1.678045e-18, 1.6765e-18, 
    1.676508e-18, 1.676551e-18, 1.676362e-18, 1.676352e-18, 1.676184e-18, 
    1.676335e-18, 1.676398e-18, 1.676564e-18, 1.67666e-18, 1.676751e-18, 
    1.676954e-18, 1.677177e-18, 1.677495e-18, 1.677726e-18, 1.677881e-18, 
    1.677787e-18, 1.677869e-18, 1.677777e-18, 1.677734e-18, 1.678213e-18, 
    1.677942e-18, 1.678352e-18, 1.67833e-18, 1.678143e-18, 1.678333e-18, 
    1.676515e-18, 1.676464e-18, 1.676281e-18, 1.676424e-18, 1.676166e-18, 
    1.676308e-18, 1.676389e-18, 1.67671e-18, 1.676785e-18, 1.676848e-18, 
    1.676979e-18, 1.677144e-18, 1.677433e-18, 1.677688e-18, 1.677924e-18, 
    1.677907e-18, 1.677913e-18, 1.677964e-18, 1.677835e-18, 1.677985e-18, 
    1.678008e-18, 1.677944e-18, 1.678327e-18, 1.678218e-18, 1.67833e-18, 
    1.678259e-18, 1.676481e-18, 1.676568e-18, 1.67652e-18, 1.676608e-18, 
    1.676545e-18, 1.676821e-18, 1.676904e-18, 1.677297e-18, 1.67714e-18, 
    1.677395e-18, 1.677167e-18, 1.677206e-18, 1.677396e-18, 1.67718e-18, 
    1.677671e-18, 1.677332e-18, 1.677966e-18, 1.677619e-18, 1.677987e-18, 
    1.677923e-18, 1.678031e-18, 1.678126e-18, 1.678248e-18, 1.67847e-18, 
    1.678419e-18, 1.678607e-18, 1.676699e-18, 1.67681e-18, 1.676803e-18, 
    1.676922e-18, 1.677009e-18, 1.677201e-18, 1.677507e-18, 1.677393e-18, 
    1.677606e-18, 1.677648e-18, 1.677326e-18, 1.677521e-18, 1.676886e-18, 
    1.676985e-18, 1.676929e-18, 1.676705e-18, 1.677415e-18, 1.677049e-18, 
    1.677729e-18, 1.677531e-18, 1.678112e-18, 1.677819e-18, 1.67839e-18, 
    1.678627e-18, 1.678865e-18, 1.679126e-18, 1.676874e-18, 1.676798e-18, 
    1.676937e-18, 1.677123e-18, 1.677305e-18, 1.677542e-18, 1.677569e-18, 
    1.677612e-18, 1.677729e-18, 1.677826e-18, 1.677623e-18, 1.67785e-18, 
    1.677002e-18, 1.677448e-18, 1.676766e-18, 1.676967e-18, 1.677113e-18, 
    1.677052e-18, 1.677381e-18, 1.677458e-18, 1.677767e-18, 1.677609e-18, 
    1.678566e-18, 1.678141e-18, 1.679336e-18, 1.678999e-18, 1.676771e-18, 
    1.676875e-18, 1.677234e-18, 1.677064e-18, 1.67756e-18, 1.677681e-18, 
    1.677782e-18, 1.677906e-18, 1.677922e-18, 1.677996e-18, 1.677874e-18, 
    1.677993e-18, 1.677543e-18, 1.677744e-18, 1.677197e-18, 1.677328e-18, 
    1.677269e-18, 1.677202e-18, 1.677409e-18, 1.677625e-18, 1.677635e-18, 
    1.677703e-18, 1.677887e-18, 1.677562e-18, 1.678611e-18, 1.677953e-18, 
    1.676989e-18, 1.677183e-18, 1.677217e-18, 1.677141e-18, 1.677669e-18, 
    1.677476e-18, 1.677995e-18, 1.677856e-18, 1.678086e-18, 1.677971e-18, 
    1.677954e-18, 1.677808e-18, 1.677716e-18, 1.677484e-18, 1.677297e-18, 
    1.677152e-18, 1.677186e-18, 1.677346e-18, 1.677639e-18, 1.677921e-18, 
    1.677859e-18, 1.678068e-18, 1.677524e-18, 1.677749e-18, 1.67766e-18, 
    1.677893e-18, 1.677389e-18, 1.677802e-18, 1.677282e-18, 1.677329e-18, 
    1.677473e-18, 1.677761e-18, 1.677832e-18, 1.677899e-18, 1.677859e-18, 
    1.677648e-18, 1.677616e-18, 1.67747e-18, 1.677428e-18, 1.677319e-18, 
    1.677226e-18, 1.677309e-18, 1.677396e-18, 1.67765e-18, 1.677877e-18, 
    1.678126e-18, 1.678189e-18, 1.678468e-18, 1.678234e-18, 1.678613e-18, 
    1.67828e-18, 1.678863e-18, 1.677834e-18, 1.67828e-18, 1.677481e-18, 
    1.677568e-18, 1.67772e-18, 1.678081e-18, 1.677892e-18, 1.678116e-18, 
    1.677615e-18, 1.677349e-18, 1.677287e-18, 1.67716e-18, 1.67729e-18, 
    1.67728e-18, 1.677403e-18, 1.677364e-18, 1.677659e-18, 1.6775e-18, 
    1.677952e-18, 1.678116e-18, 1.678586e-18, 1.678871e-18, 1.679171e-18, 
    1.679301e-18, 1.679341e-18, 1.679357e-18 ;

 MEG_acetic_acid =
  2.514304e-19, 2.514698e-19, 2.514623e-19, 2.514937e-19, 2.514766e-19, 
    2.514969e-19, 2.514387e-19, 2.51471e-19, 2.514506e-19, 2.514344e-19, 
    2.515537e-19, 2.514951e-19, 2.516178e-19, 2.515799e-19, 2.516763e-19, 
    2.516114e-19, 2.516896e-19, 2.516752e-19, 2.517203e-19, 2.517074e-19, 
    2.517636e-19, 2.517263e-19, 2.51794e-19, 2.517551e-19, 2.517608e-19, 
    2.517249e-19, 2.515077e-19, 2.515461e-19, 2.515052e-19, 2.515107e-19, 
    2.515084e-19, 2.514766e-19, 2.514601e-19, 2.514279e-19, 2.514339e-19, 
    2.514578e-19, 2.515132e-19, 2.514949e-19, 2.515426e-19, 2.515415e-19, 
    2.515941e-19, 2.515704e-19, 2.516596e-19, 2.516344e-19, 2.51708e-19, 
    2.516893e-19, 2.51707e-19, 2.517017e-19, 2.51707e-19, 2.516797e-19, 
    2.516914e-19, 2.516676e-19, 2.515747e-19, 2.516017e-19, 2.515208e-19, 
    2.51471e-19, 2.5144e-19, 2.514174e-19, 2.514206e-19, 2.514265e-19, 
    2.51458e-19, 2.514882e-19, 2.515111e-19, 2.515263e-19, 2.515414e-19, 
    2.51585e-19, 2.516099e-19, 2.516643e-19, 2.516551e-19, 2.516712e-19, 
    2.516875e-19, 2.51714e-19, 2.517097e-19, 2.517213e-19, 2.516713e-19, 
    2.517042e-19, 2.516498e-19, 2.516646e-19, 2.515428e-19, 2.515e-19, 
    2.514795e-19, 2.514636e-19, 2.51423e-19, 2.514509e-19, 2.514398e-19, 
    2.514667e-19, 2.514835e-19, 2.514753e-19, 2.515267e-19, 2.515066e-19, 
    2.516114e-19, 2.515662e-19, 2.516856e-19, 2.516571e-19, 2.516926e-19, 
    2.516746e-19, 2.517052e-19, 2.516776e-19, 2.517258e-19, 2.51736e-19, 
    2.517289e-19, 2.517568e-19, 2.51676e-19, 2.517067e-19, 2.51475e-19, 
    2.514763e-19, 2.514827e-19, 2.514544e-19, 2.514528e-19, 2.514276e-19, 
    2.514502e-19, 2.514597e-19, 2.514846e-19, 2.514989e-19, 2.515127e-19, 
    2.51543e-19, 2.515765e-19, 2.516242e-19, 2.516589e-19, 2.516821e-19, 
    2.51668e-19, 2.516804e-19, 2.516665e-19, 2.516601e-19, 2.51732e-19, 
    2.516913e-19, 2.517528e-19, 2.517495e-19, 2.517215e-19, 2.517499e-19, 
    2.514772e-19, 2.514696e-19, 2.514422e-19, 2.514636e-19, 2.514249e-19, 
    2.514463e-19, 2.514583e-19, 2.515065e-19, 2.515177e-19, 2.515272e-19, 
    2.515468e-19, 2.515716e-19, 2.51615e-19, 2.516532e-19, 2.516886e-19, 
    2.51686e-19, 2.516869e-19, 2.516945e-19, 2.516753e-19, 2.516977e-19, 
    2.517012e-19, 2.516916e-19, 2.51749e-19, 2.517326e-19, 2.517494e-19, 
    2.517388e-19, 2.514721e-19, 2.514851e-19, 2.514781e-19, 2.514912e-19, 
    2.514818e-19, 2.515231e-19, 2.515356e-19, 2.515945e-19, 2.51571e-19, 
    2.516092e-19, 2.51575e-19, 2.515809e-19, 2.516093e-19, 2.515771e-19, 
    2.516506e-19, 2.515997e-19, 2.516948e-19, 2.516429e-19, 2.51698e-19, 
    2.516884e-19, 2.517046e-19, 2.517188e-19, 2.517372e-19, 2.517704e-19, 
    2.517628e-19, 2.517911e-19, 2.515048e-19, 2.515214e-19, 2.515204e-19, 
    2.515382e-19, 2.515513e-19, 2.515802e-19, 2.516261e-19, 2.51609e-19, 
    2.51641e-19, 2.516472e-19, 2.51599e-19, 2.516281e-19, 2.51533e-19, 
    2.515478e-19, 2.515393e-19, 2.515058e-19, 2.516123e-19, 2.515573e-19, 
    2.516594e-19, 2.516296e-19, 2.517167e-19, 2.516729e-19, 2.517585e-19, 
    2.51794e-19, 2.518297e-19, 2.518689e-19, 2.515311e-19, 2.515197e-19, 
    2.515405e-19, 2.515684e-19, 2.515957e-19, 2.516313e-19, 2.516353e-19, 
    2.516418e-19, 2.516593e-19, 2.516738e-19, 2.516434e-19, 2.516775e-19, 
    2.515503e-19, 2.516173e-19, 2.515149e-19, 2.51545e-19, 2.51567e-19, 
    2.515579e-19, 2.516072e-19, 2.516186e-19, 2.516651e-19, 2.516413e-19, 
    2.517848e-19, 2.517211e-19, 2.519004e-19, 2.518498e-19, 2.515156e-19, 
    2.515313e-19, 2.515851e-19, 2.515596e-19, 2.51634e-19, 2.516521e-19, 
    2.516673e-19, 2.516859e-19, 2.516883e-19, 2.516994e-19, 2.516812e-19, 
    2.516989e-19, 2.516314e-19, 2.516616e-19, 2.515795e-19, 2.515992e-19, 
    2.515903e-19, 2.515802e-19, 2.516113e-19, 2.516437e-19, 2.516452e-19, 
    2.516555e-19, 2.51683e-19, 2.516343e-19, 2.517916e-19, 2.516929e-19, 
    2.515483e-19, 2.515774e-19, 2.515825e-19, 2.515711e-19, 2.516503e-19, 
    2.516214e-19, 2.516993e-19, 2.516784e-19, 2.517128e-19, 2.516956e-19, 
    2.516931e-19, 2.516712e-19, 2.516574e-19, 2.516226e-19, 2.515946e-19, 
    2.515728e-19, 2.51578e-19, 2.516019e-19, 2.516459e-19, 2.516882e-19, 
    2.516788e-19, 2.517102e-19, 2.516285e-19, 2.516623e-19, 2.51649e-19, 
    2.516839e-19, 2.516084e-19, 2.516703e-19, 2.515923e-19, 2.515993e-19, 
    2.516209e-19, 2.516641e-19, 2.516748e-19, 2.516849e-19, 2.516789e-19, 
    2.516472e-19, 2.516423e-19, 2.516206e-19, 2.516142e-19, 2.515978e-19, 
    2.515839e-19, 2.515964e-19, 2.516094e-19, 2.516475e-19, 2.516815e-19, 
    2.517189e-19, 2.517284e-19, 2.517702e-19, 2.51735e-19, 2.51792e-19, 
    2.517419e-19, 2.518295e-19, 2.516751e-19, 2.517421e-19, 2.516221e-19, 
    2.516352e-19, 2.51658e-19, 2.517122e-19, 2.516838e-19, 2.517174e-19, 
    2.516422e-19, 2.516023e-19, 2.51593e-19, 2.51574e-19, 2.515934e-19, 
    2.515919e-19, 2.516105e-19, 2.516046e-19, 2.516488e-19, 2.516251e-19, 
    2.516928e-19, 2.517173e-19, 2.517878e-19, 2.518307e-19, 2.518757e-19, 
    2.518951e-19, 2.519011e-19, 2.519036e-19 ;

 MEG_acetone =
  8.435195e-17, 8.436054e-17, 8.435891e-17, 8.436576e-17, 8.436202e-17, 
    8.436646e-17, 8.435377e-17, 8.436082e-17, 8.435636e-17, 8.435283e-17, 
    8.437885e-17, 8.436608e-17, 8.439285e-17, 8.438457e-17, 8.440562e-17, 
    8.439146e-17, 8.440851e-17, 8.440538e-17, 8.441523e-17, 8.441242e-17, 
    8.442467e-17, 8.441653e-17, 8.443132e-17, 8.442281e-17, 8.442408e-17, 
    8.441623e-17, 8.436881e-17, 8.43772e-17, 8.436827e-17, 8.436948e-17, 
    8.436897e-17, 8.436204e-17, 8.435843e-17, 8.435141e-17, 8.435272e-17, 
    8.435794e-17, 8.437003e-17, 8.436603e-17, 8.437643e-17, 8.43762e-17, 
    8.438769e-17, 8.43825e-17, 8.440198e-17, 8.439647e-17, 8.441254e-17, 
    8.440847e-17, 8.441232e-17, 8.441117e-17, 8.441233e-17, 8.440637e-17, 
    8.440892e-17, 8.440373e-17, 8.438344e-17, 8.438934e-17, 8.437167e-17, 
    8.436082e-17, 8.435405e-17, 8.434912e-17, 8.434981e-17, 8.435111e-17, 
    8.435797e-17, 8.436457e-17, 8.436956e-17, 8.437287e-17, 8.437617e-17, 
    8.43857e-17, 8.439112e-17, 8.440301e-17, 8.4401e-17, 8.440451e-17, 
    8.440807e-17, 8.441385e-17, 8.441292e-17, 8.441544e-17, 8.440452e-17, 
    8.441172e-17, 8.439983e-17, 8.440306e-17, 8.437649e-17, 8.436714e-17, 
    8.436267e-17, 8.43592e-17, 8.435033e-17, 8.435643e-17, 8.435401e-17, 
    8.435988e-17, 8.436353e-17, 8.436175e-17, 8.437297e-17, 8.436858e-17, 
    8.439144e-17, 8.438159e-17, 8.440765e-17, 8.440143e-17, 8.440917e-17, 
    8.440525e-17, 8.441192e-17, 8.440591e-17, 8.441642e-17, 8.441865e-17, 
    8.441712e-17, 8.44232e-17, 8.440556e-17, 8.441226e-17, 8.436167e-17, 
    8.436196e-17, 8.436336e-17, 8.435718e-17, 8.435683e-17, 8.435135e-17, 
    8.435628e-17, 8.435833e-17, 8.436379e-17, 8.436691e-17, 8.436991e-17, 
    8.437653e-17, 8.438384e-17, 8.439425e-17, 8.440182e-17, 8.440689e-17, 
    8.440382e-17, 8.440652e-17, 8.440348e-17, 8.440208e-17, 8.441778e-17, 
    8.44089e-17, 8.442232e-17, 8.44216e-17, 8.441548e-17, 8.442168e-17, 
    8.436217e-17, 8.43605e-17, 8.435452e-17, 8.43592e-17, 8.435076e-17, 
    8.435541e-17, 8.435804e-17, 8.436854e-17, 8.437099e-17, 8.437308e-17, 
    8.437735e-17, 8.438277e-17, 8.439224e-17, 8.440058e-17, 8.44083e-17, 
    8.440775e-17, 8.440794e-17, 8.44096e-17, 8.44054e-17, 8.44103e-17, 
    8.441107e-17, 8.440897e-17, 8.44215e-17, 8.441792e-17, 8.442158e-17, 
    8.441927e-17, 8.436106e-17, 8.436389e-17, 8.436235e-17, 8.436522e-17, 
    8.436315e-17, 8.437219e-17, 8.43749e-17, 8.438777e-17, 8.438263e-17, 
    8.439097e-17, 8.438352e-17, 8.43848e-17, 8.4391e-17, 8.438396e-17, 
    8.440001e-17, 8.438891e-17, 8.440967e-17, 8.439832e-17, 8.441037e-17, 
    8.440827e-17, 8.44118e-17, 8.441491e-17, 8.441892e-17, 8.442618e-17, 
    8.442452e-17, 8.443068e-17, 8.436818e-17, 8.437181e-17, 8.43716e-17, 
    8.437549e-17, 8.437833e-17, 8.438464e-17, 8.439466e-17, 8.439092e-17, 
    8.439791e-17, 8.439927e-17, 8.438873e-17, 8.439509e-17, 8.437433e-17, 
    8.437757e-17, 8.437572e-17, 8.436841e-17, 8.439164e-17, 8.437964e-17, 
    8.440193e-17, 8.439543e-17, 8.441445e-17, 8.440487e-17, 8.442358e-17, 
    8.443132e-17, 8.443913e-17, 8.444768e-17, 8.437392e-17, 8.437144e-17, 
    8.437598e-17, 8.438207e-17, 8.438803e-17, 8.439581e-17, 8.439666e-17, 
    8.439808e-17, 8.440192e-17, 8.440509e-17, 8.439844e-17, 8.440589e-17, 
    8.43781e-17, 8.439273e-17, 8.43704e-17, 8.437697e-17, 8.438176e-17, 
    8.437977e-17, 8.439053e-17, 8.439303e-17, 8.440317e-17, 8.439799e-17, 
    8.442931e-17, 8.441541e-17, 8.445456e-17, 8.444351e-17, 8.437054e-17, 
    8.437396e-17, 8.438572e-17, 8.438014e-17, 8.439638e-17, 8.440034e-17, 
    8.440366e-17, 8.440773e-17, 8.440824e-17, 8.441067e-17, 8.440668e-17, 
    8.441055e-17, 8.439582e-17, 8.440241e-17, 8.43845e-17, 8.438879e-17, 
    8.438686e-17, 8.438465e-17, 8.439144e-17, 8.439851e-17, 8.439884e-17, 
    8.440108e-17, 8.440708e-17, 8.439645e-17, 8.443079e-17, 8.440925e-17, 
    8.437768e-17, 8.438404e-17, 8.438515e-17, 8.438265e-17, 8.439994e-17, 
    8.439364e-17, 8.441064e-17, 8.440607e-17, 8.44136e-17, 8.440984e-17, 
    8.440928e-17, 8.44045e-17, 8.440149e-17, 8.43939e-17, 8.438779e-17, 
    8.438304e-17, 8.438416e-17, 8.438938e-17, 8.439898e-17, 8.440821e-17, 
    8.440616e-17, 8.441303e-17, 8.43952e-17, 8.440257e-17, 8.439967e-17, 
    8.440728e-17, 8.439079e-17, 8.440431e-17, 8.438728e-17, 8.438881e-17, 
    8.439353e-17, 8.440296e-17, 8.44053e-17, 8.44075e-17, 8.440618e-17, 
    8.439926e-17, 8.43982e-17, 8.439345e-17, 8.439205e-17, 8.438849e-17, 
    8.438546e-17, 8.438819e-17, 8.439101e-17, 8.439934e-17, 8.440675e-17, 
    8.441492e-17, 8.441699e-17, 8.442612e-17, 8.441845e-17, 8.443087e-17, 
    8.441994e-17, 8.443907e-17, 8.440534e-17, 8.441998e-17, 8.43938e-17, 
    8.439666e-17, 8.440163e-17, 8.441346e-17, 8.440725e-17, 8.44146e-17, 
    8.439818e-17, 8.438948e-17, 8.438744e-17, 8.438329e-17, 8.438754e-17, 
    8.43872e-17, 8.439125e-17, 8.438996e-17, 8.439961e-17, 8.439443e-17, 
    8.440922e-17, 8.441458e-17, 8.442997e-17, 8.443932e-17, 8.444915e-17, 
    8.445341e-17, 8.445472e-17, 8.445525e-17 ;

 MEG_carene_3 =
  3.259626e-17, 3.259965e-17, 3.259901e-17, 3.260172e-17, 3.260024e-17, 
    3.260199e-17, 3.259697e-17, 3.259976e-17, 3.2598e-17, 3.25966e-17, 
    3.260689e-17, 3.260184e-17, 3.261243e-17, 3.260915e-17, 3.261748e-17, 
    3.261188e-17, 3.261862e-17, 3.261738e-17, 3.262127e-17, 3.262016e-17, 
    3.262501e-17, 3.262179e-17, 3.262763e-17, 3.262427e-17, 3.262477e-17, 
    3.262167e-17, 3.260292e-17, 3.260624e-17, 3.260271e-17, 3.260319e-17, 
    3.260299e-17, 3.260025e-17, 3.259882e-17, 3.259604e-17, 3.259656e-17, 
    3.259863e-17, 3.26034e-17, 3.260182e-17, 3.260594e-17, 3.260585e-17, 
    3.261038e-17, 3.260834e-17, 3.261603e-17, 3.261386e-17, 3.262021e-17, 
    3.26186e-17, 3.262012e-17, 3.261967e-17, 3.262013e-17, 3.261777e-17, 
    3.261878e-17, 3.261673e-17, 3.260871e-17, 3.261104e-17, 3.260406e-17, 
    3.259976e-17, 3.259709e-17, 3.259513e-17, 3.259541e-17, 3.259592e-17, 
    3.259864e-17, 3.260125e-17, 3.260322e-17, 3.260453e-17, 3.260583e-17, 
    3.26096e-17, 3.261174e-17, 3.261644e-17, 3.261565e-17, 3.261704e-17, 
    3.261844e-17, 3.262073e-17, 3.262036e-17, 3.262136e-17, 3.261704e-17, 
    3.261989e-17, 3.261519e-17, 3.261646e-17, 3.260596e-17, 3.260226e-17, 
    3.260049e-17, 3.259913e-17, 3.259562e-17, 3.259803e-17, 3.259707e-17, 
    3.259939e-17, 3.260084e-17, 3.260013e-17, 3.260456e-17, 3.260283e-17, 
    3.261187e-17, 3.260798e-17, 3.261828e-17, 3.261582e-17, 3.261888e-17, 
    3.261733e-17, 3.261997e-17, 3.261759e-17, 3.262174e-17, 3.262262e-17, 
    3.262202e-17, 3.262442e-17, 3.261745e-17, 3.26201e-17, 3.26001e-17, 
    3.260021e-17, 3.260077e-17, 3.259832e-17, 3.259819e-17, 3.259602e-17, 
    3.259797e-17, 3.259878e-17, 3.260094e-17, 3.260217e-17, 3.260336e-17, 
    3.260598e-17, 3.260887e-17, 3.261298e-17, 3.261597e-17, 3.261797e-17, 
    3.261676e-17, 3.261783e-17, 3.261663e-17, 3.261608e-17, 3.262228e-17, 
    3.261877e-17, 3.262408e-17, 3.262379e-17, 3.262137e-17, 3.262382e-17, 
    3.26003e-17, 3.259964e-17, 3.259727e-17, 3.259913e-17, 3.259579e-17, 
    3.259762e-17, 3.259867e-17, 3.260282e-17, 3.260379e-17, 3.260461e-17, 
    3.26063e-17, 3.260844e-17, 3.261218e-17, 3.261548e-17, 3.261853e-17, 
    3.261832e-17, 3.261839e-17, 3.261905e-17, 3.261739e-17, 3.261932e-17, 
    3.261963e-17, 3.26188e-17, 3.262375e-17, 3.262234e-17, 3.262378e-17, 
    3.262287e-17, 3.259986e-17, 3.260098e-17, 3.260037e-17, 3.26015e-17, 
    3.260069e-17, 3.260426e-17, 3.260533e-17, 3.261042e-17, 3.260839e-17, 
    3.261168e-17, 3.260874e-17, 3.260925e-17, 3.261169e-17, 3.260891e-17, 
    3.261526e-17, 3.261087e-17, 3.261907e-17, 3.261459e-17, 3.261935e-17, 
    3.261852e-17, 3.261992e-17, 3.262114e-17, 3.262273e-17, 3.26256e-17, 
    3.262495e-17, 3.262738e-17, 3.260268e-17, 3.260411e-17, 3.260403e-17, 
    3.260556e-17, 3.260669e-17, 3.260918e-17, 3.261314e-17, 3.261167e-17, 
    3.261442e-17, 3.261496e-17, 3.26108e-17, 3.261332e-17, 3.260511e-17, 
    3.260638e-17, 3.260566e-17, 3.260276e-17, 3.261195e-17, 3.26072e-17, 
    3.261602e-17, 3.261345e-17, 3.262097e-17, 3.261718e-17, 3.262458e-17, 
    3.262763e-17, 3.263072e-17, 3.26341e-17, 3.260494e-17, 3.260396e-17, 
    3.260576e-17, 3.260816e-17, 3.261052e-17, 3.261359e-17, 3.261393e-17, 
    3.26145e-17, 3.261601e-17, 3.261726e-17, 3.261463e-17, 3.261758e-17, 
    3.26066e-17, 3.261238e-17, 3.260355e-17, 3.260615e-17, 3.260804e-17, 
    3.260725e-17, 3.261151e-17, 3.26125e-17, 3.261651e-17, 3.261446e-17, 
    3.262684e-17, 3.262134e-17, 3.263682e-17, 3.263245e-17, 3.260361e-17, 
    3.260496e-17, 3.260961e-17, 3.26074e-17, 3.261382e-17, 3.261539e-17, 
    3.26167e-17, 3.261831e-17, 3.261851e-17, 3.261947e-17, 3.26179e-17, 
    3.261942e-17, 3.26136e-17, 3.261621e-17, 3.260912e-17, 3.261082e-17, 
    3.261006e-17, 3.260918e-17, 3.261187e-17, 3.261467e-17, 3.26148e-17, 
    3.261568e-17, 3.261805e-17, 3.261385e-17, 3.262742e-17, 3.261891e-17, 
    3.260643e-17, 3.260894e-17, 3.260939e-17, 3.26084e-17, 3.261523e-17, 
    3.261274e-17, 3.261946e-17, 3.261765e-17, 3.262063e-17, 3.261914e-17, 
    3.261892e-17, 3.261704e-17, 3.261584e-17, 3.261284e-17, 3.261043e-17, 
    3.260855e-17, 3.260899e-17, 3.261106e-17, 3.261485e-17, 3.26185e-17, 
    3.261769e-17, 3.26204e-17, 3.261336e-17, 3.261627e-17, 3.261512e-17, 
    3.261813e-17, 3.261161e-17, 3.261696e-17, 3.261023e-17, 3.261083e-17, 
    3.261269e-17, 3.261642e-17, 3.261735e-17, 3.261822e-17, 3.26177e-17, 
    3.261496e-17, 3.261454e-17, 3.261266e-17, 3.261211e-17, 3.26107e-17, 
    3.26095e-17, 3.261058e-17, 3.26117e-17, 3.261499e-17, 3.261793e-17, 
    3.262115e-17, 3.262197e-17, 3.262558e-17, 3.262254e-17, 3.262746e-17, 
    3.262314e-17, 3.26307e-17, 3.261737e-17, 3.262315e-17, 3.26128e-17, 
    3.261393e-17, 3.26159e-17, 3.262057e-17, 3.261812e-17, 3.262102e-17, 
    3.261453e-17, 3.261109e-17, 3.261029e-17, 3.260865e-17, 3.261033e-17, 
    3.261019e-17, 3.261179e-17, 3.261128e-17, 3.26151e-17, 3.261305e-17, 
    3.26189e-17, 3.262102e-17, 3.26271e-17, 3.26308e-17, 3.263468e-17, 
    3.263636e-17, 3.263688e-17, 3.263709e-17 ;

 MEG_ethanol =
  1.676203e-18, 1.676465e-18, 1.676415e-18, 1.676624e-18, 1.67651e-18, 
    1.676646e-18, 1.676258e-18, 1.676474e-18, 1.676337e-18, 1.67623e-18, 
    1.677024e-18, 1.676634e-18, 1.677452e-18, 1.677199e-18, 1.677842e-18, 
    1.67741e-18, 1.67793e-18, 1.677835e-18, 1.678135e-18, 1.67805e-18, 
    1.678424e-18, 1.678175e-18, 1.678627e-18, 1.678367e-18, 1.678406e-18, 
    1.678166e-18, 1.676718e-18, 1.676974e-18, 1.676701e-18, 1.676738e-18, 
    1.676723e-18, 1.676511e-18, 1.676401e-18, 1.676186e-18, 1.676226e-18, 
    1.676386e-18, 1.676755e-18, 1.676633e-18, 1.676951e-18, 1.676944e-18, 
    1.677294e-18, 1.677136e-18, 1.677731e-18, 1.677563e-18, 1.678053e-18, 
    1.677929e-18, 1.678047e-18, 1.678012e-18, 1.678047e-18, 1.677865e-18, 
    1.677943e-18, 1.677784e-18, 1.677165e-18, 1.677345e-18, 1.676805e-18, 
    1.676474e-18, 1.676267e-18, 1.676116e-18, 1.676137e-18, 1.676177e-18, 
    1.676387e-18, 1.676588e-18, 1.676741e-18, 1.676842e-18, 1.676942e-18, 
    1.677234e-18, 1.677399e-18, 1.677762e-18, 1.677701e-18, 1.677808e-18, 
    1.677917e-18, 1.678093e-18, 1.678065e-18, 1.678142e-18, 1.677808e-18, 
    1.678028e-18, 1.677665e-18, 1.677764e-18, 1.676952e-18, 1.676667e-18, 
    1.67653e-18, 1.676424e-18, 1.676153e-18, 1.67634e-18, 1.676266e-18, 
    1.676445e-18, 1.676556e-18, 1.676502e-18, 1.676845e-18, 1.676711e-18, 
    1.677409e-18, 1.677108e-18, 1.677904e-18, 1.677714e-18, 1.67795e-18, 
    1.677831e-18, 1.678035e-18, 1.677851e-18, 1.678172e-18, 1.67824e-18, 
    1.678193e-18, 1.678379e-18, 1.67784e-18, 1.678045e-18, 1.6765e-18, 
    1.676508e-18, 1.676551e-18, 1.676362e-18, 1.676352e-18, 1.676184e-18, 
    1.676335e-18, 1.676398e-18, 1.676564e-18, 1.67666e-18, 1.676751e-18, 
    1.676954e-18, 1.677177e-18, 1.677495e-18, 1.677726e-18, 1.677881e-18, 
    1.677787e-18, 1.677869e-18, 1.677777e-18, 1.677734e-18, 1.678213e-18, 
    1.677942e-18, 1.678352e-18, 1.67833e-18, 1.678143e-18, 1.678333e-18, 
    1.676515e-18, 1.676464e-18, 1.676281e-18, 1.676424e-18, 1.676166e-18, 
    1.676308e-18, 1.676389e-18, 1.67671e-18, 1.676785e-18, 1.676848e-18, 
    1.676979e-18, 1.677144e-18, 1.677433e-18, 1.677688e-18, 1.677924e-18, 
    1.677907e-18, 1.677913e-18, 1.677964e-18, 1.677835e-18, 1.677985e-18, 
    1.678008e-18, 1.677944e-18, 1.678327e-18, 1.678218e-18, 1.67833e-18, 
    1.678259e-18, 1.676481e-18, 1.676568e-18, 1.67652e-18, 1.676608e-18, 
    1.676545e-18, 1.676821e-18, 1.676904e-18, 1.677297e-18, 1.67714e-18, 
    1.677395e-18, 1.677167e-18, 1.677206e-18, 1.677396e-18, 1.67718e-18, 
    1.677671e-18, 1.677332e-18, 1.677966e-18, 1.677619e-18, 1.677987e-18, 
    1.677923e-18, 1.678031e-18, 1.678126e-18, 1.678248e-18, 1.67847e-18, 
    1.678419e-18, 1.678607e-18, 1.676699e-18, 1.67681e-18, 1.676803e-18, 
    1.676922e-18, 1.677009e-18, 1.677201e-18, 1.677507e-18, 1.677393e-18, 
    1.677606e-18, 1.677648e-18, 1.677326e-18, 1.677521e-18, 1.676886e-18, 
    1.676985e-18, 1.676929e-18, 1.676705e-18, 1.677415e-18, 1.677049e-18, 
    1.677729e-18, 1.677531e-18, 1.678112e-18, 1.677819e-18, 1.67839e-18, 
    1.678627e-18, 1.678865e-18, 1.679126e-18, 1.676874e-18, 1.676798e-18, 
    1.676937e-18, 1.677123e-18, 1.677305e-18, 1.677542e-18, 1.677569e-18, 
    1.677612e-18, 1.677729e-18, 1.677826e-18, 1.677623e-18, 1.67785e-18, 
    1.677002e-18, 1.677448e-18, 1.676766e-18, 1.676967e-18, 1.677113e-18, 
    1.677052e-18, 1.677381e-18, 1.677458e-18, 1.677767e-18, 1.677609e-18, 
    1.678566e-18, 1.678141e-18, 1.679336e-18, 1.678999e-18, 1.676771e-18, 
    1.676875e-18, 1.677234e-18, 1.677064e-18, 1.67756e-18, 1.677681e-18, 
    1.677782e-18, 1.677906e-18, 1.677922e-18, 1.677996e-18, 1.677874e-18, 
    1.677993e-18, 1.677543e-18, 1.677744e-18, 1.677197e-18, 1.677328e-18, 
    1.677269e-18, 1.677202e-18, 1.677409e-18, 1.677625e-18, 1.677635e-18, 
    1.677703e-18, 1.677887e-18, 1.677562e-18, 1.678611e-18, 1.677953e-18, 
    1.676989e-18, 1.677183e-18, 1.677217e-18, 1.677141e-18, 1.677669e-18, 
    1.677476e-18, 1.677995e-18, 1.677856e-18, 1.678086e-18, 1.677971e-18, 
    1.677954e-18, 1.677808e-18, 1.677716e-18, 1.677484e-18, 1.677297e-18, 
    1.677152e-18, 1.677186e-18, 1.677346e-18, 1.677639e-18, 1.677921e-18, 
    1.677859e-18, 1.678068e-18, 1.677524e-18, 1.677749e-18, 1.67766e-18, 
    1.677893e-18, 1.677389e-18, 1.677802e-18, 1.677282e-18, 1.677329e-18, 
    1.677473e-18, 1.677761e-18, 1.677832e-18, 1.677899e-18, 1.677859e-18, 
    1.677648e-18, 1.677616e-18, 1.67747e-18, 1.677428e-18, 1.677319e-18, 
    1.677226e-18, 1.677309e-18, 1.677396e-18, 1.67765e-18, 1.677877e-18, 
    1.678126e-18, 1.678189e-18, 1.678468e-18, 1.678234e-18, 1.678613e-18, 
    1.67828e-18, 1.678863e-18, 1.677834e-18, 1.67828e-18, 1.677481e-18, 
    1.677568e-18, 1.67772e-18, 1.678081e-18, 1.677892e-18, 1.678116e-18, 
    1.677615e-18, 1.677349e-18, 1.677287e-18, 1.67716e-18, 1.67729e-18, 
    1.67728e-18, 1.677403e-18, 1.677364e-18, 1.677659e-18, 1.6775e-18, 
    1.677952e-18, 1.678116e-18, 1.678586e-18, 1.678871e-18, 1.679171e-18, 
    1.679301e-18, 1.679341e-18, 1.679357e-18 ;

 MEG_formaldehyde =
  3.352405e-19, 3.35293e-19, 3.352831e-19, 3.353249e-19, 3.353021e-19, 
    3.353292e-19, 3.352516e-19, 3.352947e-19, 3.352675e-19, 3.352459e-19, 
    3.354049e-19, 3.353269e-19, 3.354904e-19, 3.354398e-19, 3.355684e-19, 
    3.354819e-19, 3.355861e-19, 3.35567e-19, 3.356271e-19, 3.356099e-19, 
    3.356848e-19, 3.35635e-19, 3.357253e-19, 3.356734e-19, 3.356811e-19, 
    3.356332e-19, 3.353435e-19, 3.353948e-19, 3.353403e-19, 3.353476e-19, 
    3.353446e-19, 3.353022e-19, 3.352802e-19, 3.352372e-19, 3.352452e-19, 
    3.352771e-19, 3.35351e-19, 3.353266e-19, 3.353901e-19, 3.353887e-19, 
    3.354589e-19, 3.354272e-19, 3.355461e-19, 3.355125e-19, 3.356106e-19, 
    3.355858e-19, 3.356093e-19, 3.356023e-19, 3.356094e-19, 3.35573e-19, 
    3.355885e-19, 3.355569e-19, 3.354329e-19, 3.35469e-19, 3.35361e-19, 
    3.352947e-19, 3.352533e-19, 3.352232e-19, 3.352275e-19, 3.352354e-19, 
    3.352773e-19, 3.353176e-19, 3.353481e-19, 3.353684e-19, 3.353885e-19, 
    3.354467e-19, 3.354798e-19, 3.355524e-19, 3.355402e-19, 3.355616e-19, 
    3.355833e-19, 3.356187e-19, 3.35613e-19, 3.356284e-19, 3.355617e-19, 
    3.356057e-19, 3.35533e-19, 3.355527e-19, 3.353905e-19, 3.353333e-19, 
    3.353061e-19, 3.352848e-19, 3.352307e-19, 3.352679e-19, 3.352531e-19, 
    3.35289e-19, 3.353113e-19, 3.353004e-19, 3.353689e-19, 3.353421e-19, 
    3.354818e-19, 3.354216e-19, 3.355808e-19, 3.355428e-19, 3.355901e-19, 
    3.355661e-19, 3.356069e-19, 3.355702e-19, 3.356344e-19, 3.356479e-19, 
    3.356386e-19, 3.356758e-19, 3.355681e-19, 3.35609e-19, 3.352999e-19, 
    3.353017e-19, 3.353103e-19, 3.352725e-19, 3.352704e-19, 3.352368e-19, 
    3.35267e-19, 3.352796e-19, 3.353129e-19, 3.353319e-19, 3.353503e-19, 
    3.353907e-19, 3.354354e-19, 3.354989e-19, 3.355452e-19, 3.355761e-19, 
    3.355574e-19, 3.355739e-19, 3.355553e-19, 3.355467e-19, 3.356426e-19, 
    3.355885e-19, 3.356704e-19, 3.35666e-19, 3.356286e-19, 3.356665e-19, 
    3.35303e-19, 3.352928e-19, 3.352562e-19, 3.352848e-19, 3.352332e-19, 
    3.352617e-19, 3.352778e-19, 3.353419e-19, 3.353569e-19, 3.353697e-19, 
    3.353957e-19, 3.354288e-19, 3.354866e-19, 3.355376e-19, 3.355848e-19, 
    3.355814e-19, 3.355825e-19, 3.355927e-19, 3.35567e-19, 3.355969e-19, 
    3.356017e-19, 3.355889e-19, 3.356654e-19, 3.356436e-19, 3.356659e-19, 
    3.356517e-19, 3.352962e-19, 3.353135e-19, 3.353041e-19, 3.353216e-19, 
    3.35309e-19, 3.353642e-19, 3.353808e-19, 3.354593e-19, 3.354279e-19, 
    3.354789e-19, 3.354334e-19, 3.354413e-19, 3.354791e-19, 3.354361e-19, 
    3.355342e-19, 3.354663e-19, 3.355931e-19, 3.355238e-19, 3.355974e-19, 
    3.355845e-19, 3.356061e-19, 3.356251e-19, 3.356496e-19, 3.356939e-19, 
    3.356838e-19, 3.357214e-19, 3.353397e-19, 3.353619e-19, 3.353606e-19, 
    3.353843e-19, 3.354017e-19, 3.354403e-19, 3.355015e-19, 3.354787e-19, 
    3.355213e-19, 3.355296e-19, 3.354653e-19, 3.355041e-19, 3.353773e-19, 
    3.353971e-19, 3.353858e-19, 3.353411e-19, 3.35483e-19, 3.354097e-19, 
    3.355458e-19, 3.355062e-19, 3.356223e-19, 3.355638e-19, 3.356781e-19, 
    3.357253e-19, 3.35773e-19, 3.358252e-19, 3.353747e-19, 3.353596e-19, 
    3.353873e-19, 3.354246e-19, 3.35461e-19, 3.355085e-19, 3.355137e-19, 
    3.355224e-19, 3.355458e-19, 3.355651e-19, 3.355245e-19, 3.355701e-19, 
    3.354003e-19, 3.354897e-19, 3.353532e-19, 3.353934e-19, 3.354226e-19, 
    3.354105e-19, 3.354762e-19, 3.354915e-19, 3.355534e-19, 3.355218e-19, 
    3.357131e-19, 3.356282e-19, 3.358672e-19, 3.357998e-19, 3.353541e-19, 
    3.35375e-19, 3.354468e-19, 3.354127e-19, 3.35512e-19, 3.355362e-19, 
    3.355564e-19, 3.355813e-19, 3.355844e-19, 3.355992e-19, 3.355749e-19, 
    3.355985e-19, 3.355086e-19, 3.355488e-19, 3.354394e-19, 3.354656e-19, 
    3.354538e-19, 3.354403e-19, 3.354818e-19, 3.35525e-19, 3.35527e-19, 
    3.355406e-19, 3.355774e-19, 3.355124e-19, 3.357221e-19, 3.355906e-19, 
    3.353977e-19, 3.354366e-19, 3.354434e-19, 3.354281e-19, 3.355337e-19, 
    3.354953e-19, 3.35599e-19, 3.355712e-19, 3.356171e-19, 3.355942e-19, 
    3.355907e-19, 3.355616e-19, 3.355432e-19, 3.354968e-19, 3.354595e-19, 
    3.354304e-19, 3.354373e-19, 3.354692e-19, 3.355279e-19, 3.355842e-19, 
    3.355717e-19, 3.356136e-19, 3.355047e-19, 3.355498e-19, 3.35532e-19, 
    3.355786e-19, 3.354778e-19, 3.355604e-19, 3.354564e-19, 3.354657e-19, 
    3.354945e-19, 3.355521e-19, 3.355665e-19, 3.355799e-19, 3.355718e-19, 
    3.355296e-19, 3.355231e-19, 3.354941e-19, 3.354855e-19, 3.354637e-19, 
    3.354452e-19, 3.354619e-19, 3.354792e-19, 3.3553e-19, 3.355753e-19, 
    3.356252e-19, 3.356378e-19, 3.356936e-19, 3.356467e-19, 3.357226e-19, 
    3.356559e-19, 3.357726e-19, 3.355667e-19, 3.356561e-19, 3.354962e-19, 
    3.355136e-19, 3.35544e-19, 3.356163e-19, 3.355784e-19, 3.356232e-19, 
    3.355229e-19, 3.354698e-19, 3.354574e-19, 3.35432e-19, 3.35458e-19, 
    3.354559e-19, 3.354806e-19, 3.354727e-19, 3.355317e-19, 3.355001e-19, 
    3.355904e-19, 3.356231e-19, 3.357171e-19, 3.357742e-19, 3.358342e-19, 
    3.358602e-19, 3.358682e-19, 3.358714e-19 ;

 MEG_isoprene =
  2.294416e-19, 2.294854e-19, 2.29477e-19, 2.295119e-19, 2.294929e-19, 
    2.295155e-19, 2.294509e-19, 2.294868e-19, 2.29464e-19, 2.29446e-19, 
    2.295786e-19, 2.295136e-19, 2.296498e-19, 2.296077e-19, 2.297148e-19, 
    2.296428e-19, 2.297295e-19, 2.297136e-19, 2.297637e-19, 2.297494e-19, 
    2.298117e-19, 2.297703e-19, 2.298455e-19, 2.298023e-19, 2.298087e-19, 
    2.297688e-19, 2.295275e-19, 2.295702e-19, 2.295247e-19, 2.295309e-19, 
    2.295283e-19, 2.29493e-19, 2.294746e-19, 2.294388e-19, 2.294455e-19, 
    2.294721e-19, 2.295337e-19, 2.295133e-19, 2.295663e-19, 2.295651e-19, 
    2.296236e-19, 2.295972e-19, 2.296963e-19, 2.296682e-19, 2.2975e-19, 
    2.297293e-19, 2.297489e-19, 2.29743e-19, 2.297489e-19, 2.297186e-19, 
    2.297316e-19, 2.297052e-19, 2.296019e-19, 2.29632e-19, 2.295421e-19, 
    2.294868e-19, 2.294523e-19, 2.294272e-19, 2.294307e-19, 2.294373e-19, 
    2.294723e-19, 2.295059e-19, 2.295313e-19, 2.295482e-19, 2.295649e-19, 
    2.296134e-19, 2.29641e-19, 2.297015e-19, 2.296913e-19, 2.297091e-19, 
    2.297273e-19, 2.297567e-19, 2.297519e-19, 2.297647e-19, 2.297092e-19, 
    2.297458e-19, 2.296853e-19, 2.297018e-19, 2.295666e-19, 2.295189e-19, 
    2.294962e-19, 2.294785e-19, 2.294334e-19, 2.294644e-19, 2.294521e-19, 
    2.29482e-19, 2.295006e-19, 2.294915e-19, 2.295486e-19, 2.295263e-19, 
    2.296427e-19, 2.295925e-19, 2.297251e-19, 2.296935e-19, 2.297328e-19, 
    2.297129e-19, 2.297469e-19, 2.297163e-19, 2.297697e-19, 2.297811e-19, 
    2.297732e-19, 2.298042e-19, 2.297145e-19, 2.297486e-19, 2.294911e-19, 
    2.294926e-19, 2.294997e-19, 2.294682e-19, 2.294665e-19, 2.294385e-19, 
    2.294637e-19, 2.294741e-19, 2.295019e-19, 2.295178e-19, 2.295331e-19, 
    2.295668e-19, 2.29604e-19, 2.296569e-19, 2.296955e-19, 2.297212e-19, 
    2.297056e-19, 2.297194e-19, 2.297039e-19, 2.296968e-19, 2.297766e-19, 
    2.297315e-19, 2.297997e-19, 2.297961e-19, 2.297649e-19, 2.297965e-19, 
    2.294936e-19, 2.294851e-19, 2.294547e-19, 2.294785e-19, 2.294355e-19, 
    2.294592e-19, 2.294726e-19, 2.295261e-19, 2.295386e-19, 2.295492e-19, 
    2.29571e-19, 2.295985e-19, 2.296467e-19, 2.296892e-19, 2.297284e-19, 
    2.297256e-19, 2.297266e-19, 2.29735e-19, 2.297137e-19, 2.297386e-19, 
    2.297425e-19, 2.297318e-19, 2.297956e-19, 2.297774e-19, 2.29796e-19, 
    2.297842e-19, 2.29488e-19, 2.295024e-19, 2.294946e-19, 2.295092e-19, 
    2.294987e-19, 2.295447e-19, 2.295585e-19, 2.29624e-19, 2.295978e-19, 
    2.296403e-19, 2.296023e-19, 2.296089e-19, 2.296404e-19, 2.296046e-19, 
    2.296863e-19, 2.296298e-19, 2.297354e-19, 2.296777e-19, 2.297389e-19, 
    2.297282e-19, 2.297462e-19, 2.29762e-19, 2.297825e-19, 2.298193e-19, 
    2.298109e-19, 2.298422e-19, 2.295243e-19, 2.295428e-19, 2.295417e-19, 
    2.295614e-19, 2.295759e-19, 2.296081e-19, 2.29659e-19, 2.2964e-19, 
    2.296755e-19, 2.296825e-19, 2.296289e-19, 2.296613e-19, 2.295556e-19, 
    2.295721e-19, 2.295627e-19, 2.295254e-19, 2.296437e-19, 2.295826e-19, 
    2.29696e-19, 2.29663e-19, 2.297597e-19, 2.29711e-19, 2.298061e-19, 
    2.298455e-19, 2.298852e-19, 2.299286e-19, 2.295535e-19, 2.295408e-19, 
    2.295639e-19, 2.29595e-19, 2.296253e-19, 2.296649e-19, 2.296692e-19, 
    2.296765e-19, 2.29696e-19, 2.297121e-19, 2.296783e-19, 2.297162e-19, 
    2.295748e-19, 2.296492e-19, 2.295355e-19, 2.29569e-19, 2.295934e-19, 
    2.295832e-19, 2.29638e-19, 2.296507e-19, 2.297024e-19, 2.29676e-19, 
    2.298353e-19, 2.297646e-19, 2.299636e-19, 2.299074e-19, 2.295363e-19, 
    2.295537e-19, 2.296135e-19, 2.295851e-19, 2.296678e-19, 2.296879e-19, 
    2.297048e-19, 2.297255e-19, 2.297281e-19, 2.297405e-19, 2.297202e-19, 
    2.297399e-19, 2.29665e-19, 2.296985e-19, 2.296073e-19, 2.296292e-19, 
    2.296193e-19, 2.296081e-19, 2.296427e-19, 2.296786e-19, 2.296803e-19, 
    2.296917e-19, 2.297223e-19, 2.296682e-19, 2.298428e-19, 2.297333e-19, 
    2.295726e-19, 2.29605e-19, 2.296107e-19, 2.295979e-19, 2.296859e-19, 
    2.296539e-19, 2.297403e-19, 2.297171e-19, 2.297554e-19, 2.297363e-19, 
    2.297334e-19, 2.297091e-19, 2.296938e-19, 2.296552e-19, 2.296241e-19, 
    2.295999e-19, 2.296056e-19, 2.296322e-19, 2.29681e-19, 2.29728e-19, 
    2.297176e-19, 2.297525e-19, 2.296618e-19, 2.296993e-19, 2.296845e-19, 
    2.297233e-19, 2.296393e-19, 2.297081e-19, 2.296215e-19, 2.296292e-19, 
    2.296533e-19, 2.297013e-19, 2.297132e-19, 2.297244e-19, 2.297177e-19, 
    2.296825e-19, 2.296771e-19, 2.296529e-19, 2.296458e-19, 2.296276e-19, 
    2.296122e-19, 2.296261e-19, 2.296405e-19, 2.296828e-19, 2.297206e-19, 
    2.297621e-19, 2.297726e-19, 2.298191e-19, 2.2978e-19, 2.298432e-19, 
    2.297877e-19, 2.298849e-19, 2.297134e-19, 2.297878e-19, 2.296547e-19, 
    2.296692e-19, 2.296945e-19, 2.297547e-19, 2.297231e-19, 2.297605e-19, 
    2.296769e-19, 2.296327e-19, 2.296223e-19, 2.296012e-19, 2.296228e-19, 
    2.296211e-19, 2.296417e-19, 2.296351e-19, 2.296842e-19, 2.296579e-19, 
    2.297331e-19, 2.297604e-19, 2.298386e-19, 2.298862e-19, 2.299361e-19, 
    2.299577e-19, 2.299644e-19, 2.299671e-19 ;

 MEG_methanol =
  5.797964e-17, 5.798532e-17, 5.798424e-17, 5.798877e-17, 5.79863e-17, 
    5.798923e-17, 5.798084e-17, 5.798551e-17, 5.798256e-17, 5.798023e-17, 
    5.799742e-17, 5.798898e-17, 5.800666e-17, 5.800119e-17, 5.801509e-17, 
    5.800574e-17, 5.8017e-17, 5.801493e-17, 5.802143e-17, 5.801957e-17, 
    5.802765e-17, 5.802229e-17, 5.803203e-17, 5.802644e-17, 5.802726e-17, 
    5.802209e-17, 5.799079e-17, 5.799633e-17, 5.799043e-17, 5.799122e-17, 
    5.799089e-17, 5.798631e-17, 5.798393e-17, 5.797929e-17, 5.798015e-17, 
    5.79836e-17, 5.799159e-17, 5.798895e-17, 5.799582e-17, 5.799566e-17, 
    5.800325e-17, 5.799983e-17, 5.801268e-17, 5.800905e-17, 5.801965e-17, 
    5.801697e-17, 5.801951e-17, 5.801875e-17, 5.801951e-17, 5.801558e-17, 
    5.801726e-17, 5.801384e-17, 5.800045e-17, 5.800434e-17, 5.799267e-17, 
    5.798551e-17, 5.798103e-17, 5.797777e-17, 5.797823e-17, 5.797909e-17, 
    5.798362e-17, 5.798799e-17, 5.799128e-17, 5.799347e-17, 5.799564e-17, 
    5.800194e-17, 5.800552e-17, 5.801337e-17, 5.801204e-17, 5.801435e-17, 
    5.80167e-17, 5.802052e-17, 5.80199e-17, 5.802156e-17, 5.801437e-17, 
    5.801912e-17, 5.801126e-17, 5.80134e-17, 5.799586e-17, 5.798968e-17, 
    5.798673e-17, 5.798443e-17, 5.797858e-17, 5.79826e-17, 5.798101e-17, 
    5.798488e-17, 5.798729e-17, 5.798612e-17, 5.799353e-17, 5.799064e-17, 
    5.800573e-17, 5.799922e-17, 5.801643e-17, 5.801232e-17, 5.801743e-17, 
    5.801484e-17, 5.801925e-17, 5.801528e-17, 5.802221e-17, 5.802368e-17, 
    5.802267e-17, 5.802669e-17, 5.801505e-17, 5.801947e-17, 5.798607e-17, 
    5.798625e-17, 5.798719e-17, 5.79831e-17, 5.798287e-17, 5.797925e-17, 
    5.798251e-17, 5.798387e-17, 5.798747e-17, 5.798953e-17, 5.799152e-17, 
    5.799588e-17, 5.800071e-17, 5.800758e-17, 5.801258e-17, 5.801592e-17, 
    5.80139e-17, 5.801568e-17, 5.801367e-17, 5.801275e-17, 5.802311e-17, 
    5.801726e-17, 5.80261e-17, 5.802563e-17, 5.802159e-17, 5.802569e-17, 
    5.79864e-17, 5.798529e-17, 5.798134e-17, 5.798443e-17, 5.797886e-17, 
    5.798193e-17, 5.798367e-17, 5.799061e-17, 5.799223e-17, 5.799361e-17, 
    5.799643e-17, 5.8e-17, 5.800625e-17, 5.801176e-17, 5.801685e-17, 
    5.801649e-17, 5.801662e-17, 5.801771e-17, 5.801494e-17, 5.801817e-17, 
    5.801868e-17, 5.80173e-17, 5.802556e-17, 5.802321e-17, 5.802562e-17, 
    5.802409e-17, 5.798566e-17, 5.798754e-17, 5.798652e-17, 5.798841e-17, 
    5.798705e-17, 5.799302e-17, 5.799481e-17, 5.80033e-17, 5.799991e-17, 
    5.800542e-17, 5.80005e-17, 5.800135e-17, 5.800544e-17, 5.800079e-17, 
    5.801139e-17, 5.800406e-17, 5.801776e-17, 5.801027e-17, 5.801822e-17, 
    5.801683e-17, 5.801916e-17, 5.802121e-17, 5.802386e-17, 5.802865e-17, 
    5.802755e-17, 5.803162e-17, 5.799037e-17, 5.799277e-17, 5.799263e-17, 
    5.799519e-17, 5.799707e-17, 5.800124e-17, 5.800785e-17, 5.800539e-17, 
    5.801e-17, 5.80109e-17, 5.800394e-17, 5.800814e-17, 5.799443e-17, 
    5.799657e-17, 5.799535e-17, 5.799052e-17, 5.800586e-17, 5.799793e-17, 
    5.801265e-17, 5.800836e-17, 5.802091e-17, 5.801459e-17, 5.802693e-17, 
    5.803204e-17, 5.803718e-17, 5.804282e-17, 5.799416e-17, 5.799252e-17, 
    5.799552e-17, 5.799954e-17, 5.800348e-17, 5.800861e-17, 5.800918e-17, 
    5.801012e-17, 5.801264e-17, 5.801474e-17, 5.801034e-17, 5.801527e-17, 
    5.799692e-17, 5.800658e-17, 5.799183e-17, 5.799617e-17, 5.799934e-17, 
    5.799802e-17, 5.800513e-17, 5.800677e-17, 5.801347e-17, 5.801005e-17, 
    5.803072e-17, 5.802155e-17, 5.804736e-17, 5.804007e-17, 5.799193e-17, 
    5.799419e-17, 5.800195e-17, 5.799826e-17, 5.800899e-17, 5.801161e-17, 
    5.80138e-17, 5.801648e-17, 5.801682e-17, 5.801842e-17, 5.801579e-17, 
    5.801834e-17, 5.800862e-17, 5.801298e-17, 5.800114e-17, 5.800398e-17, 
    5.80027e-17, 5.800124e-17, 5.800573e-17, 5.801039e-17, 5.801061e-17, 
    5.801209e-17, 5.801605e-17, 5.800904e-17, 5.803169e-17, 5.801748e-17, 
    5.799664e-17, 5.800084e-17, 5.800158e-17, 5.799993e-17, 5.801134e-17, 
    5.800719e-17, 5.80184e-17, 5.801538e-17, 5.802035e-17, 5.801787e-17, 
    5.80175e-17, 5.801435e-17, 5.801236e-17, 5.800735e-17, 5.800332e-17, 
    5.800018e-17, 5.800092e-17, 5.800437e-17, 5.801071e-17, 5.80168e-17, 
    5.801544e-17, 5.801997e-17, 5.800821e-17, 5.801307e-17, 5.801116e-17, 
    5.801618e-17, 5.80053e-17, 5.801422e-17, 5.800298e-17, 5.800399e-17, 
    5.800711e-17, 5.801333e-17, 5.801488e-17, 5.801633e-17, 5.801546e-17, 
    5.801089e-17, 5.80102e-17, 5.800705e-17, 5.800613e-17, 5.800378e-17, 
    5.800178e-17, 5.800358e-17, 5.800544e-17, 5.801094e-17, 5.801583e-17, 
    5.802123e-17, 5.802259e-17, 5.802861e-17, 5.802355e-17, 5.803175e-17, 
    5.802454e-17, 5.803715e-17, 5.801491e-17, 5.802456e-17, 5.800728e-17, 
    5.800917e-17, 5.801245e-17, 5.802025e-17, 5.801617e-17, 5.802101e-17, 
    5.801018e-17, 5.800443e-17, 5.800309e-17, 5.800035e-17, 5.800315e-17, 
    5.800293e-17, 5.80056e-17, 5.800475e-17, 5.801112e-17, 5.80077e-17, 
    5.801746e-17, 5.8021e-17, 5.803115e-17, 5.803732e-17, 5.804379e-17, 
    5.80466e-17, 5.804746e-17, 5.804782e-17 ;

 MEG_pinene_a =
  4.795984e-17, 4.796504e-17, 4.796405e-17, 4.79682e-17, 4.796594e-17, 
    4.796863e-17, 4.796094e-17, 4.796521e-17, 4.796251e-17, 4.796037e-17, 
    4.797613e-17, 4.79684e-17, 4.798461e-17, 4.79796e-17, 4.799235e-17, 
    4.798377e-17, 4.79941e-17, 4.799221e-17, 4.799817e-17, 4.799647e-17, 
    4.800389e-17, 4.799895e-17, 4.800791e-17, 4.800276e-17, 4.800353e-17, 
    4.799878e-17, 4.797005e-17, 4.797514e-17, 4.796973e-17, 4.797046e-17, 
    4.797015e-17, 4.796595e-17, 4.796377e-17, 4.795951e-17, 4.79603e-17, 
    4.796347e-17, 4.797079e-17, 4.796837e-17, 4.797467e-17, 4.797453e-17, 
    4.798149e-17, 4.797835e-17, 4.799014e-17, 4.798681e-17, 4.799654e-17, 
    4.799407e-17, 4.799641e-17, 4.799571e-17, 4.799641e-17, 4.79928e-17, 
    4.799435e-17, 4.799121e-17, 4.797892e-17, 4.798249e-17, 4.797179e-17, 
    4.796521e-17, 4.796111e-17, 4.795812e-17, 4.795854e-17, 4.795933e-17, 
    4.796349e-17, 4.796749e-17, 4.797051e-17, 4.797251e-17, 4.797451e-17, 
    4.798028e-17, 4.798357e-17, 4.799077e-17, 4.798955e-17, 4.799168e-17, 
    4.799383e-17, 4.799734e-17, 4.799677e-17, 4.79983e-17, 4.799169e-17, 
    4.799605e-17, 4.798884e-17, 4.79908e-17, 4.79747e-17, 4.796904e-17, 
    4.796633e-17, 4.796423e-17, 4.795886e-17, 4.796255e-17, 4.796109e-17, 
    4.796464e-17, 4.796685e-17, 4.796578e-17, 4.797257e-17, 4.796991e-17, 
    4.798376e-17, 4.797779e-17, 4.799358e-17, 4.798981e-17, 4.79945e-17, 
    4.799212e-17, 4.799617e-17, 4.799253e-17, 4.799889e-17, 4.800024e-17, 
    4.799931e-17, 4.8003e-17, 4.799232e-17, 4.799637e-17, 4.796573e-17, 
    4.79659e-17, 4.796675e-17, 4.796301e-17, 4.79628e-17, 4.795947e-17, 
    4.796246e-17, 4.796371e-17, 4.796701e-17, 4.79689e-17, 4.797072e-17, 
    4.797473e-17, 4.797916e-17, 4.798546e-17, 4.799005e-17, 4.799312e-17, 
    4.799126e-17, 4.79929e-17, 4.799105e-17, 4.79902e-17, 4.799971e-17, 
    4.799434e-17, 4.800247e-17, 4.800203e-17, 4.799832e-17, 4.800208e-17, 
    4.796603e-17, 4.796502e-17, 4.796139e-17, 4.796423e-17, 4.795911e-17, 
    4.796193e-17, 4.796353e-17, 4.796989e-17, 4.797138e-17, 4.797264e-17, 
    4.797523e-17, 4.797851e-17, 4.798424e-17, 4.79893e-17, 4.799397e-17, 
    4.799364e-17, 4.799375e-17, 4.799476e-17, 4.799222e-17, 4.799518e-17, 
    4.799565e-17, 4.799438e-17, 4.800197e-17, 4.79998e-17, 4.800202e-17, 
    4.800062e-17, 4.796535e-17, 4.796708e-17, 4.796614e-17, 4.796788e-17, 
    4.796663e-17, 4.79721e-17, 4.797374e-17, 4.798154e-17, 4.797842e-17, 
    4.798348e-17, 4.797896e-17, 4.797974e-17, 4.798349e-17, 4.797923e-17, 
    4.798895e-17, 4.798223e-17, 4.79948e-17, 4.798793e-17, 4.799522e-17, 
    4.799395e-17, 4.799609e-17, 4.799797e-17, 4.80004e-17, 4.80048e-17, 
    4.800379e-17, 4.800753e-17, 4.796967e-17, 4.797187e-17, 4.797174e-17, 
    4.79741e-17, 4.797582e-17, 4.797965e-17, 4.798571e-17, 4.798345e-17, 
    4.798768e-17, 4.79885e-17, 4.798212e-17, 4.798597e-17, 4.79734e-17, 
    4.797536e-17, 4.797424e-17, 4.796981e-17, 4.798388e-17, 4.797661e-17, 
    4.799011e-17, 4.798618e-17, 4.799769e-17, 4.799189e-17, 4.800323e-17, 
    4.800792e-17, 4.801264e-17, 4.801782e-17, 4.797315e-17, 4.797164e-17, 
    4.797439e-17, 4.797808e-17, 4.79817e-17, 4.798641e-17, 4.798692e-17, 
    4.798779e-17, 4.799011e-17, 4.799203e-17, 4.7988e-17, 4.799251e-17, 
    4.797568e-17, 4.798455e-17, 4.797101e-17, 4.797499e-17, 4.797789e-17, 
    4.797669e-17, 4.798321e-17, 4.798472e-17, 4.799087e-17, 4.798773e-17, 
    4.80067e-17, 4.799828e-17, 4.802198e-17, 4.801529e-17, 4.79711e-17, 
    4.797317e-17, 4.798029e-17, 4.797692e-17, 4.798676e-17, 4.798915e-17, 
    4.799116e-17, 4.799362e-17, 4.799394e-17, 4.799541e-17, 4.799299e-17, 
    4.799534e-17, 4.798641e-17, 4.799041e-17, 4.797956e-17, 4.798216e-17, 
    4.798098e-17, 4.797965e-17, 4.798376e-17, 4.798804e-17, 4.798824e-17, 
    4.79896e-17, 4.799324e-17, 4.79868e-17, 4.800759e-17, 4.799454e-17, 
    4.797543e-17, 4.797927e-17, 4.797995e-17, 4.797844e-17, 4.798891e-17, 
    4.79851e-17, 4.799539e-17, 4.799263e-17, 4.799718e-17, 4.799491e-17, 
    4.799457e-17, 4.799167e-17, 4.798985e-17, 4.798525e-17, 4.798155e-17, 
    4.797867e-17, 4.797935e-17, 4.798251e-17, 4.798833e-17, 4.799392e-17, 
    4.799268e-17, 4.799683e-17, 4.798604e-17, 4.79905e-17, 4.798874e-17, 
    4.799336e-17, 4.798337e-17, 4.799155e-17, 4.798124e-17, 4.798217e-17, 
    4.798502e-17, 4.799074e-17, 4.799216e-17, 4.799349e-17, 4.799269e-17, 
    4.79885e-17, 4.798786e-17, 4.798498e-17, 4.798413e-17, 4.798197e-17, 
    4.798013e-17, 4.798179e-17, 4.79835e-17, 4.798854e-17, 4.799304e-17, 
    4.799798e-17, 4.799924e-17, 4.800477e-17, 4.800012e-17, 4.800764e-17, 
    4.800103e-17, 4.80126e-17, 4.799219e-17, 4.800104e-17, 4.798519e-17, 
    4.798692e-17, 4.798994e-17, 4.79971e-17, 4.799334e-17, 4.799778e-17, 
    4.798784e-17, 4.798257e-17, 4.798134e-17, 4.797883e-17, 4.79814e-17, 
    4.798119e-17, 4.798365e-17, 4.798286e-17, 4.798871e-17, 4.798557e-17, 
    4.799453e-17, 4.799778e-17, 4.80071e-17, 4.801276e-17, 4.801871e-17, 
    4.802129e-17, 4.802208e-17, 4.80224e-17 ;

 MEG_thujene_a =
  1.210136e-18, 1.210262e-18, 1.210238e-18, 1.210339e-18, 1.210284e-18, 
    1.210349e-18, 1.210163e-18, 1.210266e-18, 1.210201e-18, 1.210149e-18, 
    1.210531e-18, 1.210343e-18, 1.210736e-18, 1.210615e-18, 1.210924e-18, 
    1.210716e-18, 1.210966e-18, 1.21092e-18, 1.211065e-18, 1.211024e-18, 
    1.211203e-18, 1.211084e-18, 1.211301e-18, 1.211176e-18, 1.211195e-18, 
    1.211079e-18, 1.210384e-18, 1.210507e-18, 1.210376e-18, 1.210393e-18, 
    1.210386e-18, 1.210284e-18, 1.210231e-18, 1.210128e-18, 1.210147e-18, 
    1.210224e-18, 1.210401e-18, 1.210343e-18, 1.210495e-18, 1.210492e-18, 
    1.210661e-18, 1.210585e-18, 1.21087e-18, 1.21079e-18, 1.211025e-18, 
    1.210966e-18, 1.211022e-18, 1.211005e-18, 1.211022e-18, 1.210935e-18, 
    1.210972e-18, 1.210896e-18, 1.210598e-18, 1.210685e-18, 1.210425e-18, 
    1.210266e-18, 1.210167e-18, 1.210094e-18, 1.210105e-18, 1.210124e-18, 
    1.210224e-18, 1.210321e-18, 1.210395e-18, 1.210443e-18, 1.210491e-18, 
    1.210631e-18, 1.210711e-18, 1.210885e-18, 1.210856e-18, 1.210907e-18, 
    1.21096e-18, 1.211045e-18, 1.211031e-18, 1.211068e-18, 1.210908e-18, 
    1.211013e-18, 1.210839e-18, 1.210886e-18, 1.210496e-18, 1.210359e-18, 
    1.210293e-18, 1.210242e-18, 1.210112e-18, 1.210202e-18, 1.210166e-18, 
    1.210252e-18, 1.210306e-18, 1.21028e-18, 1.210445e-18, 1.21038e-18, 
    1.210716e-18, 1.210571e-18, 1.210954e-18, 1.210862e-18, 1.210976e-18, 
    1.210918e-18, 1.211016e-18, 1.210928e-18, 1.211082e-18, 1.211115e-18, 
    1.211092e-18, 1.211182e-18, 1.210923e-18, 1.211021e-18, 1.210279e-18, 
    1.210283e-18, 1.210304e-18, 1.210213e-18, 1.210208e-18, 1.210127e-18, 
    1.2102e-18, 1.21023e-18, 1.21031e-18, 1.210356e-18, 1.2104e-18, 
    1.210497e-18, 1.210604e-18, 1.210757e-18, 1.210868e-18, 1.210942e-18, 
    1.210897e-18, 1.210937e-18, 1.210892e-18, 1.210872e-18, 1.211102e-18, 
    1.210972e-18, 1.211169e-18, 1.211158e-18, 1.211068e-18, 1.21116e-18, 
    1.210286e-18, 1.210261e-18, 1.210174e-18, 1.210242e-18, 1.210119e-18, 
    1.210187e-18, 1.210226e-18, 1.21038e-18, 1.210416e-18, 1.210446e-18, 
    1.210509e-18, 1.210588e-18, 1.210727e-18, 1.21085e-18, 1.210963e-18, 
    1.210955e-18, 1.210958e-18, 1.210982e-18, 1.21092e-18, 1.210992e-18, 
    1.211004e-18, 1.210973e-18, 1.211157e-18, 1.211104e-18, 1.211158e-18, 
    1.211124e-18, 1.21027e-18, 1.210311e-18, 1.210289e-18, 1.210331e-18, 
    1.2103e-18, 1.210433e-18, 1.210473e-18, 1.210662e-18, 1.210586e-18, 
    1.210709e-18, 1.210599e-18, 1.210618e-18, 1.210709e-18, 1.210606e-18, 
    1.210841e-18, 1.210678e-18, 1.210983e-18, 1.210817e-18, 1.210993e-18, 
    1.210963e-18, 1.211014e-18, 1.21106e-18, 1.211119e-18, 1.211225e-18, 
    1.211201e-18, 1.211292e-18, 1.210374e-18, 1.210428e-18, 1.210424e-18, 
    1.210481e-18, 1.210523e-18, 1.210616e-18, 1.210763e-18, 1.210708e-18, 
    1.210811e-18, 1.21083e-18, 1.210676e-18, 1.210769e-18, 1.210465e-18, 
    1.210512e-18, 1.210485e-18, 1.210378e-18, 1.210719e-18, 1.210542e-18, 
    1.21087e-18, 1.210774e-18, 1.211053e-18, 1.210913e-18, 1.211187e-18, 
    1.211301e-18, 1.211415e-18, 1.211541e-18, 1.210458e-18, 1.210422e-18, 
    1.210489e-18, 1.210578e-18, 1.210666e-18, 1.21078e-18, 1.210792e-18, 
    1.210813e-18, 1.210869e-18, 1.210916e-18, 1.210818e-18, 1.210928e-18, 
    1.21052e-18, 1.210735e-18, 1.210407e-18, 1.210503e-18, 1.210574e-18, 
    1.210544e-18, 1.210702e-18, 1.210739e-18, 1.210888e-18, 1.210812e-18, 
    1.211271e-18, 1.211067e-18, 1.211642e-18, 1.21148e-18, 1.210409e-18, 
    1.210459e-18, 1.210632e-18, 1.21055e-18, 1.210788e-18, 1.210846e-18, 
    1.210895e-18, 1.210955e-18, 1.210962e-18, 1.210998e-18, 1.210939e-18, 
    1.210996e-18, 1.21078e-18, 1.210877e-18, 1.210614e-18, 1.210677e-18, 
    1.210648e-18, 1.210616e-18, 1.210716e-18, 1.210819e-18, 1.210824e-18, 
    1.210857e-18, 1.210945e-18, 1.210789e-18, 1.211293e-18, 1.210977e-18, 
    1.210514e-18, 1.210607e-18, 1.210623e-18, 1.210587e-18, 1.21084e-18, 
    1.210748e-18, 1.210997e-18, 1.21093e-18, 1.211041e-18, 1.210986e-18, 
    1.210977e-18, 1.210907e-18, 1.210863e-18, 1.210752e-18, 1.210662e-18, 
    1.210592e-18, 1.210609e-18, 1.210685e-18, 1.210826e-18, 1.210962e-18, 
    1.210932e-18, 1.211032e-18, 1.210771e-18, 1.210879e-18, 1.210836e-18, 
    1.210948e-18, 1.210706e-18, 1.210904e-18, 1.210655e-18, 1.210677e-18, 
    1.210746e-18, 1.210885e-18, 1.210919e-18, 1.210951e-18, 1.210932e-18, 
    1.21083e-18, 1.210815e-18, 1.210745e-18, 1.210725e-18, 1.210672e-18, 
    1.210628e-18, 1.210668e-18, 1.210709e-18, 1.210832e-18, 1.21094e-18, 
    1.21106e-18, 1.211091e-18, 1.211225e-18, 1.211112e-18, 1.211294e-18, 
    1.211134e-18, 1.211415e-18, 1.21092e-18, 1.211134e-18, 1.21075e-18, 
    1.210792e-18, 1.210865e-18, 1.211039e-18, 1.210948e-18, 1.211055e-18, 
    1.210815e-18, 1.210687e-18, 1.210657e-18, 1.210596e-18, 1.210658e-18, 
    1.210653e-18, 1.210713e-18, 1.210694e-18, 1.210836e-18, 1.21076e-18, 
    1.210977e-18, 1.211055e-18, 1.211281e-18, 1.211418e-18, 1.211563e-18, 
    1.211625e-18, 1.211644e-18, 1.211652e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -9.889281e-26, 1.840507e-25, 2.856907e-25, 1.565805e-25, 7.691677e-26, 
    -3.845826e-26, 8.241083e-26, 2.747033e-26, 8.257808e-32, 1.346043e-25, 
    4.560062e-25, 1.565805e-25, -1.703155e-25, -2.829435e-25, -2.472314e-26, 
    -2.747024e-25, 8.241157e-27, 1.703156e-25, -1.346041e-25, -4.724882e-25, 
    1.538335e-25, 4.834764e-25, -3.488721e-25, -1.950387e-25, -1.840506e-25, 
    -1.071339e-25, -2.747024e-25, -3.241488e-25, -1.895446e-25, 
    -1.620744e-25, -4.285358e-25, -2.087738e-25, -2.554732e-25, 
    -2.032798e-25, 2.692085e-25, 1.0164e-25, 1.373521e-26, -2.582203e-25, 
    -3.296421e-26, 2.747033e-26, 1.098818e-26, 4.889705e-25, -1.840506e-25, 
    9.614595e-26, 6.785152e-25, -4.450179e-25, 1.867978e-25, -3.571131e-25, 
    8.790487e-26, -4.669934e-26, -6.043446e-26, 2.582204e-25, -8.241066e-26, 
    1.263632e-25, 3.021728e-25, -1.840506e-25, -2.774494e-25, -3.268959e-25, 
    -4.010655e-25, 5.494132e-27, -5.988513e-25, -1.346041e-25, -2.225089e-25, 
    1.181221e-25, 2.966788e-25, 1.236162e-25, -2.28003e-25, -5.164406e-25, 
    -4.395231e-26, 2.801966e-25, -2.197612e-26, -2.774494e-25, -1.620744e-25, 
    2.362442e-25, -2.444851e-25, -9.889281e-26, -2.582203e-25, 1.126281e-25, 
    -1.538333e-25, 1.098811e-25, -1.098802e-26, -3.571131e-25, -1.593274e-25, 
    6.867563e-25, -1.318571e-25, -6.043446e-26, 5.76876e-26, 1.675686e-25, 
    -3.021727e-25, 2.774496e-25, -1.922916e-25, -2.25256e-25, -1.565803e-25, 
    -3.598602e-25, 1.977859e-25, 1.126281e-25, 4.944653e-26, 1.071341e-25, 
    -9.339876e-26, 2.197628e-26, 3.57114e-26, 5.274289e-25, -1.565803e-25, 
    -3.488721e-25, -1.867976e-25, -5.109465e-25, -1.840506e-25, 8.515785e-26, 
    2.334972e-25, 9.339892e-26, -1.758095e-25, 1.373513e-25, -1.510863e-25, 
    -3.790893e-25, 1.236162e-25, -2.664613e-25, 3.928246e-25, -2.746942e-27, 
    6.86757e-26, -2.664613e-25, -1.620744e-25, 9.06519e-26, -1.922909e-26, 
    1.840507e-25, -5.494041e-26, 4.202949e-25, 2.08774e-25, -2.499792e-25, 
    1.236162e-25, 1.510864e-25, -3.928245e-25, 3.351371e-25, 1.346043e-25, 
    1.675686e-25, -2.637143e-25, 3.983187e-25, 1.648223e-26, -2.389911e-25, 
    -2.417381e-25, 2.225091e-25, -3.900774e-25, 1.208692e-25, -1.510863e-25, 
    -3.214018e-25, -2.582203e-25, -4.395239e-25, 2.11521e-25, -2.472321e-25, 
    1.730626e-25, 7.691677e-26, -4.148007e-25, -1.950387e-25, -3.296429e-25, 
    3.488722e-25, -6.043454e-25, -7.691661e-26, -1.620744e-25, -9.614578e-26, 
    1.373513e-25, -2.939316e-25, -7.691661e-26, -9.614578e-26, -5.439108e-25, 
    2.032799e-25, 8.790487e-26, -6.043446e-26, -1.016398e-25, -2.774494e-25, 
    -2.032798e-25, -1.126279e-25, -9.889281e-26, -1.620744e-25, 1.373513e-25, 
    6.592867e-26, 3.900776e-25, -1.593274e-25, -1.016398e-25, -5.768744e-26, 
    -1.18122e-25, 3.378841e-25, -3.983185e-25, -2.060268e-25, -2.472314e-26, 
    -1.071339e-25, 2.032799e-25, -2.747024e-25, -7.966364e-26, -2.472321e-25, 
    -4.340298e-25, -5.493967e-27, -4.010655e-25, 2.554734e-25, 1.291103e-25, 
    -3.845834e-25, -1.675684e-25, -4.422709e-25, 1.510864e-25, 1.813037e-25, 
    -2.774494e-25, -6.043446e-26, 2.692085e-25, -2.939316e-25, 5.494058e-26, 
    2.719555e-25, -1.867976e-25, 2.499793e-25, -2.499792e-25, 1.208692e-25, 
    -1.565803e-25, -3.241488e-25, 4.944653e-26, -1.565803e-25, -1.428452e-25, 
    -1.730625e-25, -2.664613e-25, -4.944636e-26, -2.554732e-25, 1.373521e-26, 
    2.747033e-26, -3.214018e-25, -4.58753e-25, 4.120545e-26, -2.747016e-26, 
    -1.126279e-25, -3.681012e-25, -1.263631e-25, -5.493967e-27, 
    -1.813036e-25, 2.801966e-25, 2.939317e-25, -1.483393e-25, -3.296421e-26, 
    2.747033e-26, 5.494058e-26, 9.889298e-26, 3.653544e-25, 3.104139e-25, 
    -2.472321e-25, -1.483393e-25, -3.351369e-25, -3.571131e-25, 1.703156e-25, 
    -2.527262e-25, -2.28003e-25, 1.346043e-25, 2.472331e-26, 3.351371e-25, 
    5.246818e-25, -6.867554e-26, 1.483394e-25, -2.747016e-26, 4.66995e-26, 
    5.658872e-25, 5.494132e-27, -2.3075e-25, -4.944636e-26, 1.950388e-25, 
    8.241083e-26, -4.944636e-26, -3.790893e-25, -5.494041e-26, 4.450181e-25, 
    -8.790471e-26, -2.801964e-25, 8.790487e-26, 4.120538e-25, 6.345628e-25, 
    -1.785565e-25, -2.005327e-25, 1.922926e-26, 3.543663e-25, 1.593275e-25, 
    2.747033e-26, 2.856907e-25, 1.648216e-25, 1.126281e-25, -1.18122e-25, 
    -4.944636e-26, 3.076668e-25, 1.181221e-25, -6.043446e-26, 1.840507e-25, 
    -4.669934e-26, 1.373513e-25, -9.614578e-26, -6.318148e-26, 2.582204e-25, 
    -2.609673e-25, -3.900774e-25, 2.08774e-25, -3.46125e-25, -5.494041e-26, 
    -3.626072e-25, -1.785565e-25, 2.362442e-25, 4.120545e-26, -2.472314e-26, 
    2.389912e-25, -6.867554e-26, 4.120545e-26, -5.494041e-26, -3.735953e-25, 
    -1.20869e-25, -2.225089e-25, -1.373512e-25, 8.241157e-27, 2.747033e-26, 
    2.801966e-25, 5.494058e-26, -1.016398e-25, 1.236162e-25, -3.268959e-25, 
    7.96638e-26, -2.417381e-25, -4.50512e-25, -2.33497e-25, 4.66995e-26, 
    -4.202947e-25, -3.516191e-25, -3.681012e-25, -2.197612e-26, 1.181221e-25, 
    3.26896e-25, -1.867976e-25, -2.032798e-25, 3.296438e-26, -2.966786e-25, 
    -2.444851e-25, 1.428454e-25, -1.455922e-25, 1.950388e-25, -1.813036e-25, 
    -2.664613e-25, -2.170149e-25, 2.692085e-25, -1.538333e-25, -3.681012e-25, 
    1.895448e-25 ;

 M_LITR2C_TO_LEACHING =
  1.483394e-25, -1.758095e-25, 1.64822e-26, 1.758096e-25, -1.428452e-25, 
    -2.3075e-25, 1.593275e-25, -1.428452e-25, -1.895447e-25, -1.922912e-26, 
    -1.895447e-25, -1.043869e-25, -1.400982e-25, 1.04387e-25, 5.219352e-26, 
    1.04387e-25, -2.087738e-25, 5.494055e-26, -5.219342e-26, 2.280031e-25, 
    -4.944639e-26, -2.911846e-25, -1.043869e-25, -6.592854e-26, 
    -1.730625e-25, 1.648215e-25, -1.648209e-26, 2.582204e-25, -3.021722e-26, 
    -2.884375e-25, -1.785566e-25, -5.493996e-27, 1.675686e-25, -6.592854e-26, 
    -2.197619e-25, -2.472317e-26, 1.977858e-25, -2.197614e-26, 5.351482e-32, 
    -2.417381e-25, -6.043449e-26, -1.263631e-25, -1.373512e-25, 
    -1.867976e-25, 5.494055e-26, -9.065177e-26, 5.351459e-32, 1.758096e-25, 
    -5.493996e-27, -2.389911e-25, -6.043449e-26, -7.142259e-26, 
    -2.829435e-25, 5.768757e-26, -4.395234e-26, 6.04346e-26, 5.494055e-26, 
    -3.845829e-26, 1.867977e-25, -2.28003e-25, -2.142679e-25, -1.098805e-26, 
    2.856906e-25, -1.071339e-25, -2.334971e-25, 1.0164e-25, -1.455923e-25, 
    -6.318152e-26, -2.472317e-26, -1.648209e-26, -1.648214e-25, 
    -3.296424e-26, 2.856906e-25, -1.895447e-25, 2.362442e-25, 8.241128e-27, 
    -1.703155e-25, 7.966377e-26, -6.043449e-26, -3.845829e-26, 8.790485e-26, 
    -2.142679e-25, 1.675686e-25, -1.703155e-25, -1.346042e-25, -2.115208e-25, 
    -3.296424e-26, -2.719554e-25, -4.120532e-26, 8.790485e-26, -1.428452e-25, 
    9.889295e-26, -6.043449e-26, 3.571138e-26, 3.021728e-25, -1.291101e-25, 
    -2.637143e-25, 1.373513e-25, -1.895447e-25, 2.74703e-26, -8.241069e-26, 
    6.04346e-26, -1.098809e-25, 3.84584e-26, -9.339879e-26, 9.339889e-26, 
    -8.515771e-26, -1.593274e-25, -6.318152e-26, -1.758095e-25, 9.614592e-26, 
    -1.620744e-25, 8.790485e-26, -2.197614e-26, -1.263631e-25, -3.021727e-25, 
    1.126281e-25, -2.197619e-25, -2.747024e-25, -1.483393e-25, -4.669937e-26, 
    -3.790894e-25, -2.472317e-26, 1.593275e-25, -2.74702e-26, -1.785566e-25, 
    -2.746971e-27, -7.691664e-26, -1.18122e-25, -1.538333e-25, 1.0164e-25, 
    -3.021722e-26, 3.296435e-26, -2.197614e-26, 4.94465e-26, -1.703155e-25, 
    -7.691664e-26, -5.219342e-26, 2.225091e-25, -1.098805e-26, 2.11521e-25, 
    1.098815e-26, 2.19762e-25, 3.076668e-25, -1.098809e-25, 1.703156e-25, 
    2.14268e-25, 7.14227e-26, 1.455924e-25, -1.813036e-25, -8.515771e-26, 
    8.790485e-26, 1.126281e-25, -1.758095e-25, 1.263632e-25, -2.472322e-25, 
    -8.241069e-26, -1.648214e-25, 4.94465e-26, -3.021722e-26, -1.730625e-25, 
    -1.098809e-25, 6.04346e-26, -1.318571e-25, -2.582203e-25, -1.373512e-25, 
    -2.142679e-25, -2.032798e-25, -2.74702e-26, 6.867567e-26, -5.768747e-26, 
    1.648215e-25, 2.417382e-25, -1.043869e-25, 7.416973e-26, -2.939316e-25, 
    -3.543661e-25, 8.790485e-26, -2.389911e-25, -6.043449e-26, -2.774495e-25, 
    2.17015e-25, 4.148008e-25, -4.944639e-26, -2.609673e-25, -1.291101e-25, 
    5.494103e-27, -4.395234e-26, 8.790485e-26, 2.966787e-25, 2.362442e-25, 
    4.505121e-25, -6.592854e-26, -2.3075e-25, 1.098815e-26, -3.543661e-25, 
    -2.527262e-25, 1.950388e-25, -1.538333e-25, 2.197625e-26, 1.04387e-25, 
    6.592865e-26, -5.493996e-27, -2.115208e-25, -1.098805e-26, 4.120543e-26, 
    -7.691664e-26, -1.455923e-25, 8.515782e-26, -2.032798e-25, 1.400983e-25, 
    3.818365e-25, -6.592854e-26, -1.12628e-25, 4.94465e-26, -1.648209e-26, 
    -9.065177e-26, -1.538333e-25, -5.493996e-27, -1.593274e-25, 1.428453e-25, 
    -1.043869e-25, -7.142259e-26, -1.373512e-25, 1.758096e-25, -7.966367e-26, 
    -3.131608e-25, -7.691664e-26, 1.373518e-26, 5.494103e-27, 3.763424e-25, 
    -3.214019e-25, -1.12628e-25, -2.527262e-25, -1.648209e-26, 8.24108e-26, 
    -8.515771e-26, 1.098815e-26, -5.219342e-26, 4.395245e-26, 1.208691e-25, 
    6.318163e-26, 3.845835e-25, 2.664615e-25, 1.867977e-25, 3.84584e-26, 
    -4.944639e-26, -2.582203e-25, -1.373512e-25, -2.197614e-26, 
    -7.691664e-26, 8.24108e-26, -2.856905e-25, 8.24108e-26, 1.867977e-25, 
    1.593275e-25, -1.236161e-25, 6.318163e-26, 6.04346e-26, 1.922923e-26, 
    5.768757e-26, 1.703156e-25, 1.538334e-25, -7.691664e-26, -7.416961e-26, 
    1.620745e-25, -5.219342e-26, 1.593275e-25, -2.389911e-25, 4.94465e-26, 
    9.339889e-26, 1.895448e-25, 2.444853e-25, -3.021722e-26, -3.076667e-25, 
    1.813037e-25, -1.922912e-26, -1.813036e-25, -8.241069e-26, -1.840506e-25, 
    3.021733e-26, -9.889284e-26, -8.241069e-26, -7.691664e-26, -1.15375e-25, 
    -1.428452e-25, 1.703156e-25, 1.703156e-25, -7.966367e-26, 2.087739e-25, 
    1.483394e-25, 1.840507e-25, 9.889295e-26, 7.416973e-26, 8.24108e-26, 
    2.197625e-26, -2.527262e-25, 9.614592e-26, -8.241021e-27, -6.043449e-26, 
    2.664615e-25, 3.296435e-26, -4.395234e-26, -2.087738e-25, -2.142679e-25, 
    3.296435e-26, -3.296424e-26, 9.339889e-26, 1.758096e-25, 3.571138e-26, 
    -6.043449e-26, -1.20869e-25, 1.0164e-25, 3.021728e-25, 1.593275e-25, 
    6.318163e-26, -1.373507e-26, -2.28003e-25, 8.790485e-26, -2.197614e-26, 
    1.455924e-25, -8.241069e-26, -3.571132e-25, 1.538334e-25, -5.494044e-26, 
    9.339889e-26, -1.510863e-25, 2.747078e-27, 1.703156e-25, -7.691664e-26, 
    -3.571132e-25, 2.74703e-26, -9.889284e-26, 3.296435e-26, -1.538333e-25, 
    -1.703155e-25, 6.592865e-26, -1.565804e-25 ;

 M_LITR3C_TO_LEACHING =
  6.867565e-26, 9.339887e-26, -1.922915e-26, -3.296427e-26, 1.510866e-26, 
    3.433784e-26, 8.241101e-27, 1.236161e-25, 1.181221e-25, -4.532588e-26, 
    2.884379e-26, 1.428453e-25, -1.002664e-25, 8.241101e-27, -2.746998e-27, 
    -1.400982e-25, -1.098807e-26, 1.648217e-26, -4.257886e-26, -4.395237e-26, 
    -1.552069e-25, -3.296427e-26, 4.120564e-27, -6.043452e-26, 9.614614e-27, 
    8.241101e-27, 9.889292e-26, -5.494047e-26, 8.653131e-26, 2.675742e-32, 
    -6.867559e-26, -2.746998e-27, 1.236164e-26, 6.043457e-26, -1.387247e-25, 
    1.098813e-26, 3.159081e-26, 7.004916e-26, 8.515779e-26, 5.356701e-26, 
    -1.909182e-25, -4.120535e-26, -2.197617e-26, 4.669945e-26, -1.648212e-26, 
    -1.922915e-26, 5.768755e-26, -4.395237e-26, 3.845837e-26, 1.098813e-26, 
    -1.785566e-25, -2.747022e-26, 1.785569e-26, -5.356696e-26, 4.12054e-26, 
    8.241101e-27, 3.02173e-26, -2.747022e-26, 5.356701e-26, -1.373486e-27, 
    2.609676e-26, 4.120564e-27, -1.483393e-25, -9.065179e-26, 4.669945e-26, 
    -1.043869e-25, -7.416964e-26, 5.494052e-26, 3.845837e-26, 4.532594e-26, 
    -6.867535e-27, 1.92292e-26, -2.197617e-26, -1.634479e-25, -1.043869e-25, 
    6.592862e-26, 2.675733e-32, -5.768749e-26, -8.790477e-26, -6.455506e-26, 
    -1.09881e-25, -1.648212e-26, 4.944647e-26, 2.362442e-25, 5.906106e-26, 
    -1.236161e-25, 1.373515e-26, 6.867565e-26, -1.098807e-26, -9.61456e-27, 
    1.140016e-25, 9.202536e-26, 5.081998e-26, 1.648217e-26, 1.236164e-26, 
    -1.15375e-25, -9.20253e-26, -7.966369e-26, 1.648217e-26, 2.197622e-26, 
    -2.458587e-25, 4.395242e-26, -1.098807e-26, 2.060271e-26, -5.631398e-26, 
    5.768755e-26, -3.296427e-26, -1.346042e-25, 6.867565e-26, -5.219344e-26, 
    6.043457e-26, -3.57113e-26, 2.197622e-26, 1.648217e-26, 3.571135e-26, 
    -1.277366e-25, -8.241047e-27, -1.510861e-26, -2.47232e-26, 4.12054e-26, 
    2.675731e-32, -1.098807e-26, 2.334974e-26, -7.416964e-26, -6.043452e-26, 
    -7.416964e-26, 1.92292e-26, 5.494076e-27, -1.593274e-25, 6.867589e-27, 
    -6.592857e-26, 1.771831e-25, 6.455511e-26, 7.691672e-26, -4.257886e-26, 
    6.31816e-26, -8.927828e-26, -9.889287e-26, 1.785569e-26, 1.09881e-25, 
    -2.609671e-26, -2.609671e-26, -9.61456e-27, 1.016399e-25, 1.785569e-26, 
    -6.318154e-26, -8.241071e-26, 1.703156e-25, -6.455506e-26, 1.098813e-26, 
    1.510866e-26, -6.043452e-26, 2.747052e-27, -1.37351e-26, -1.194956e-25, 
    -1.208691e-25, 3.02173e-26, 1.07134e-25, -3.845832e-26, 9.75194e-26, 
    3.433784e-26, 6.867589e-27, 4.807296e-26, -3.296427e-26, -1.758096e-25, 
    -1.71689e-25, 1.04387e-25, 2.197622e-26, -7.142262e-26, 3.571135e-26, 
    -6.043452e-26, -2.142679e-25, -1.249896e-25, 1.04387e-25, -1.263631e-25, 
    -1.950387e-25, -1.510863e-25, -1.277366e-25, 1.318572e-25, -3.296427e-26, 
    8.241077e-26, -8.515774e-26, -8.378423e-26, -9.889287e-26, -1.936652e-25, 
    1.92292e-26, -1.455923e-25, 9.889292e-26, -8.515774e-26, -1.112545e-25, 
    -4.669939e-26, -3.983183e-26, 4.395242e-26, -2.417381e-25, 3.845837e-26, 
    1.92292e-26, -7.279613e-26, -1.15375e-25, -4.120535e-26, 1.92292e-26, 
    -3.021725e-26, -1.387247e-25, 5.494076e-27, 8.790482e-26, -2.747022e-26, 
    -5.356696e-26, -2.060266e-26, 6.31816e-26, -7.279613e-26, -8.515774e-26, 
    4.669945e-26, 9.065185e-26, 6.592862e-26, 6.867565e-26, 8.515779e-26, 
    1.63448e-25, 1.373513e-25, -8.241071e-26, -1.648212e-26, -3.57113e-26, 
    2.197622e-26, 3.845837e-26, -1.249896e-25, -8.515774e-26, -6.730208e-26, 
    -2.609671e-26, 1.977858e-25, -2.19762e-25, -4.395237e-26, -4.120511e-27, 
    -7.279613e-26, 2.472325e-26, 2.609676e-26, -6.318154e-26, 5.631404e-26, 
    -6.318154e-26, -1.016399e-25, -5.494047e-26, -4.532588e-26, 
    -1.620744e-25, 9.065185e-26, -2.747022e-26, 7.416969e-26, 5.356701e-26, 
    -6.318154e-26, -6.867559e-26, -7.691667e-26, 3.708486e-26, 1.236161e-25, 
    3.296432e-26, 5.21935e-26, -2.197617e-26, -8.241047e-27, 1.291102e-25, 
    1.936653e-25, 2.060271e-26, 2.334974e-26, -4.395237e-26, -1.071339e-25, 
    2.266296e-25, -6.867559e-26, -1.236161e-25, 1.098813e-26, -3.845832e-26, 
    2.747028e-26, -4.257886e-26, 6.043457e-26, -1.785563e-26, 7.142267e-26, 
    -4.257886e-26, -3.845832e-26, 6.455511e-26, 5.494052e-26, 4.12054e-26, 
    -3.021725e-26, 3.433784e-26, -9.065179e-26, -1.12628e-25, -3.296427e-26, 
    6.043457e-26, -2.747022e-26, -1.236161e-25, -1.318572e-25, 7.691672e-26, 
    -1.785563e-26, -6.592857e-26, -1.09881e-25, 6.043457e-26, 1.098813e-26, 
    -7.00491e-26, 2.197622e-26, -1.922915e-26, -1.09881e-25, -1.167485e-25, 
    -1.922915e-26, 6.867565e-26, -3.296427e-26, -3.296427e-26, 1.181221e-25, 
    1.510866e-26, 5.494052e-26, 3.708486e-26, -2.47232e-26, 2.675733e-32, 
    -6.592857e-26, -7.142262e-26, 3.708486e-26, 1.181221e-25, -2.060266e-26, 
    1.098813e-26, 1.112545e-25, -4.395237e-26, -2.746998e-27, -1.085074e-25, 
    9.889292e-26, -9.61456e-27, -1.277366e-25, -2.47232e-26, -1.249896e-25, 
    2.17015e-25, -2.060266e-26, 2.747052e-27, 8.515779e-26, -1.37351e-26, 
    4.944647e-26, -3.021725e-26, 1.648217e-26, -4.395237e-26, -8.241047e-27, 
    7.416969e-26, -1.867977e-25, -6.318154e-26, -6.043452e-26, 1.208691e-25, 
    4.395242e-26, 5.768755e-26, -6.318154e-26, -5.494023e-27 ;

 M_SOIL1C_TO_LEACHING =
  1.809874e-20, -1.497994e-20, 2.602791e-20, 8.224344e-21, 2.435427e-21, 
    -1.520921e-20, -3.919158e-20, 9.897008e-21, -1.050034e-20, -2.709467e-20, 
    2.168064e-20, -3.037802e-20, -2.522382e-20, 1.112773e-20, 1.710422e-22, 
    -2.867825e-20, -2.152515e-20, 4.958533e-21, 1.373732e-20, 4.3173e-21, 
    -2.002838e-20, -1.146105e-20, -5.451902e-21, 3.007125e-21, 6.669744e-22, 
    -1.54111e-20, 2.761447e-21, 2.504853e-20, -2.492724e-20, -6.268707e-21, 
    1.713546e-20, 1.292308e-20, -1.905492e-20, 1.666048e-20, 8.142375e-21, 
    1.877417e-20, -2.65851e-21, 4.112328e-21, -2.346126e-20, 6.302648e-21, 
    -2.582181e-20, 2.011148e-20, 6.134119e-21, 3.869456e-21, 1.068976e-20, 
    -5.243807e-20, 8.758437e-21, -6.604881e-21, 2.323849e-20, -2.347713e-20, 
    2.069561e-20, 1.341443e-20, 1.312663e-20, 2.066483e-21, -9.093467e-21, 
    -5.06964e-21, 5.624079e-21, 3.823368e-21, -4.213818e-21, 1.397962e-20, 
    1.050656e-20, 3.181564e-21, 1.806424e-20, -1.149047e-20, -2.950352e-20, 
    -4.619762e-20, 1.455016e-20, 1.116135e-20, 3.349991e-20, -3.878417e-20, 
    -1.915472e-20, -1.167765e-20, -1.253637e-21, 7.165802e-21, 3.527633e-21, 
    -1.282297e-20, 8.645623e-21, 3.922494e-20, -3.327453e-21, -2.285596e-20, 
    -3.118664e-20, 1.464772e-20, 1.386624e-20, 3.785748e-21, 2.269311e-20, 
    6.008309e-21, 2.578845e-20, 1.025041e-20, 4.564517e-20, -1.115316e-20, 
    5.155595e-21, 3.180168e-21, 1.937669e-20, -1.679562e-20, 1.846545e-20, 
    -1.332396e-20, 7.437502e-21, -1.611566e-20, -3.681726e-21, 3.015919e-20, 
    -1.61637e-20, -3.253412e-20, -2.257407e-20, -1.189619e-20, 2.083215e-20, 
    -5.609098e-21, 3.679372e-20, -1.685838e-20, 2.000715e-20, -1.256117e-20, 
    2.926575e-20, -1.992318e-20, -2.056725e-20, -2.945517e-20, 1.200843e-20, 
    -7.85878e-21, -3.02392e-20, 8.406998e-21, -1.631358e-21, 1.616175e-20, 
    -2.47528e-20, 1.778884e-20, -2.275304e-20, -2.114403e-20, -1.12702e-20, 
    -8.65778e-21, -8.212759e-21, -2.315283e-20, -2.394753e-22, 6.32639e-21, 
    1.209549e-20, -2.227127e-20, 2.018387e-20, -3.636479e-21, -3.838322e-20, 
    5.527245e-20, 4.313358e-21, 5.843209e-21, -8.017093e-21, -1.541589e-20, 
    3.853646e-22, 8.664017e-21, -9.422849e-21, -4.524845e-21, 1.41032e-20, 
    6.791314e-22, -2.276492e-20, 1.058036e-20, -1.755986e-20, -1.980785e-20, 
    -1.884317e-20, 1.294794e-20, -9.542146e-21, -3.834903e-20, -2.329928e-20, 
    1.243959e-20, -5.023007e-21, 1.566554e-20, 4.670003e-20, -2.607117e-20, 
    -1.403137e-20, -9.112416e-21, -6.290742e-21, -1.292915e-21, 5.891558e-21, 
    6.446287e-22, 3.26817e-20, 1.181222e-20, 1.170222e-21, -8.128633e-22, 
    2.632366e-20, -3.304896e-20, 9.839326e-21, 1.082632e-20, -1.461946e-20, 
    8.034925e-21, -3.480812e-20, 3.716382e-20, 6.245227e-21, -1.997379e-20, 
    1.777803e-21, -2.091274e-20, 1.725223e-20, -6.987689e-21, -3.02847e-20, 
    -4.898314e-21, 1.627625e-20, -1.306555e-20, 2.656822e-20, -5.631705e-21, 
    4.832323e-20, -9.957487e-21, -1.674388e-20, 2.628576e-20, 2.194215e-20, 
    -1.249304e-20, 2.039281e-20, -7.917597e-21, 2.492384e-20, -2.243017e-20, 
    8.380166e-22, -2.620405e-20, -2.537509e-20, -7.635992e-21, -2.185341e-20, 
    4.668197e-20, -6.775351e-21, 3.114309e-20, -3.475921e-20, 3.902079e-20, 
    -1.426385e-21, 1.534097e-21, -7.990544e-21, -1.058034e-20, -2.076121e-20, 
    1.201549e-20, 1.93648e-20, -8.962609e-22, -2.721269e-21, 1.555331e-20, 
    -1.095637e-20, 1.54343e-21, 2.180415e-21, -3.456835e-20, 3.36314e-20, 
    3.421298e-20, -1.740406e-20, 4.72986e-20, -9.572134e-21, 2.196449e-20, 
    -1.33808e-20, 1.884486e-20, 1.882988e-20, -9.702476e-21, 1.952991e-20, 
    1.405963e-20, -2.390999e-20, 2.145332e-20, 2.027942e-20, 1.077204e-20, 
    1.816685e-20, -1.595761e-20, 5.372196e-20, -5.082369e-21, -1.824065e-20, 
    -1.707779e-20, 4.661215e-20, -2.344856e-20, -6.615921e-21, -8.804525e-21, 
    -2.51718e-20, -3.439988e-20, -1.769898e-21, 1.428072e-20, 2.035831e-20, 
    1.997832e-20, -2.14248e-20, -2.876732e-20, 2.680827e-20, 2.544775e-20, 
    -1.498163e-20, 9.526331e-21, 1.464432e-20, 5.412313e-21, 4.948751e-20, 
    3.535009e-20, 4.577017e-20, -7.515823e-21, -4.124484e-21, -3.215494e-21, 
    2.961942e-20, 4.821683e-21, -3.634645e-20, -5.577419e-21, -2.828834e-20, 
    -7.848591e-21, 4.811242e-21, 1.838203e-20, -4.165499e-20, 1.896108e-20, 
    -1.784023e-21, 3.300232e-20, -2.492271e-20, -2.055395e-20, 2.619329e-20, 
    4.071604e-21, -1.630422e-20, 5.462353e-21, -3.501563e-20, -2.012733e-20, 
    1.393289e-21, -1.27263e-20, 1.558921e-20, -3.061351e-20, 9.42738e-21, 
    3.415191e-20, -2.138065e-20, -7.176562e-21, -3.417029e-20, 7.116056e-21, 
    -1.866875e-21, -1.602716e-20, -8.703867e-21, 3.180327e-20, 4.592566e-20, 
    -7.99563e-21, 3.386976e-20, -2.016606e-20, 2.548337e-20, 1.593384e-20, 
    -1.293351e-20, 1.719935e-20, -9.85595e-22, -3.788337e-20, -2.424162e-20, 
    -2.368039e-20, -4.011159e-20, -2.065087e-21, -8.602359e-21, 
    -6.194585e-22, 1.024474e-20, -3.076252e-20, 1.878011e-20, 9.224375e-21, 
    3.890998e-20, -3.252422e-20, -1.704441e-20, -1.041578e-20, -3.257822e-20, 
    -8.10815e-21, 7.46918e-21, -9.500043e-21, 1.65044e-20, 1.568011e-21, 
    1.823528e-20, -1.2739e-20, -1.221424e-20, -5.562438e-21 ;

 M_SOIL2C_TO_LEACHING =
  -1.020176e-20, 6.864816e-20, 3.285445e-20, -8.911674e-21, -4.515437e-20, 
    -8.105593e-21, 2.167696e-20, -2.206629e-20, 3.776828e-20, 2.326845e-20, 
    -2.544407e-20, -2.949617e-20, -8.874909e-21, 7.675009e-21, 1.23409e-20, 
    -4.169437e-21, 1.767098e-20, -1.526209e-20, 6.004088e-21, -1.233895e-20, 
    -6.588756e-21, 6.655428e-20, -1.89568e-20, -4.057298e-20, -1.487646e-20, 
    1.160523e-20, -2.10623e-20, -8.121146e-21, -7.865572e-21, 6.436925e-21, 
    1.575489e-20, 1.585554e-20, -9.857418e-21, 8.995088e-21, 1.858278e-20, 
    -7.304342e-21, -5.21234e-20, -4.202796e-21, -2.292608e-20, -2.579807e-20, 
    -3.440579e-20, -1.240933e-20, -3.890744e-20, 8.661176e-21, 1.106836e-20, 
    -4.142713e-20, -2.36787e-20, 1.515835e-20, -1.121537e-20, -1.315716e-20, 
    -2.214572e-20, -8.761261e-21, 6.847443e-21, 1.208449e-20, -6.02698e-21, 
    -2.966128e-20, 1.35202e-20, 1.735459e-20, -2.998871e-23, -1.39895e-20, 
    -5.575167e-21, -1.827318e-20, -8.359766e-21, 2.850661e-20, 1.610829e-20, 
    -2.716647e-20, 4.207065e-22, -1.288233e-20, 2.269366e-20, 2.374964e-21, 
    -1.746399e-20, 2.020193e-20, -2.344035e-20, -4.250405e-20, -4.339976e-22, 
    3.075461e-20, -1.988585e-20, 1.476022e-20, -1.201946e-20, -1.233554e-20, 
    -3.723845e-21, -1.748066e-20, -2.630668e-20, -4.3495e-20, -5.866933e-21, 
    -4.536708e-21, 2.555885e-21, -2.327327e-20, 2.195573e-20, 1.634755e-21, 
    2.284532e-22, 1.113309e-20, 7.590494e-21, -1.339575e-21, 1.566048e-20, 
    -3.021372e-20, 3.719315e-21, 6.197176e-20, -7.978648e-21, -2.318987e-20, 
    2.952417e-20, 1.530989e-20, 1.253996e-20, 8.908295e-21, -2.840002e-20, 
    1.363187e-20, 1.269291e-20, 4.787764e-20, -7.08949e-21, -9.862211e-21, 
    3.602783e-20, -2.973194e-21, -1.059309e-20, 2.808591e-20, 1.544869e-20, 
    9.079621e-21, 1.018017e-22, -2.499793e-20, 8.619881e-21, -1.628219e-20, 
    -2.636634e-20, -1.351565e-20, -7.572383e-21, 1.02586e-20, -1.082121e-20, 
    -7.501404e-21, 2.012486e-21, -2.283532e-20, 1.957089e-20, -1.638057e-20, 
    -4.444533e-21, -9.844117e-21, 1.806821e-20, 2.168574e-20, 3.365683e-20, 
    -3.101301e-20, -3.096213e-20, -9.137303e-21, 1.241725e-20, 2.098484e-20, 
    2.907896e-21, 5.598647e-21, -3.668658e-20, 2.792363e-20, 1.551907e-20, 
    5.457e-23, -2.271798e-20, -2.796264e-20, 5.456694e-21, -4.731786e-21, 
    1.38295e-20, 1.386258e-20, -8.68295e-21, -4.238784e-20, -2.573529e-20, 
    1.398642e-20, -5.906801e-21, 2.270978e-20, -1.794183e-20, 3.928796e-20, 
    6.538155e-21, -7.15082e-21, -6.137515e-21, -3.535435e-20, 3.482108e-21, 
    -2.015763e-22, -4.808092e-20, -1.278226e-20, 9.985508e-21, 1.681969e-21, 
    -8.996572e-22, -1.681937e-20, -4.232768e-21, 2.701379e-20, -2.821497e-22, 
    7.47963e-21, 2.197383e-20, -6.581963e-21, -3.293163e-20, -3.605158e-20, 
    1.055348e-20, 2.183814e-20, 2.85476e-20, -9.633496e-21, -2.083783e-20, 
    1.591377e-20, 9.762982e-21, -1.962971e-20, -3.211961e-20, 1.161034e-20, 
    1.164456e-20, 1.837044e-20, 3.89028e-22, 3.341566e-20, -8.090612e-21, 
    -1.543144e-20, -7.594991e-21, -1.443483e-20, -2.6308e-21, -5.219481e-21, 
    -1.162306e-20, -3.308882e-20, -3.12785e-20, -2.087542e-20, -1.15159e-20, 
    -2.959313e-20, -2.285314e-20, 1.555308e-21, -3.767782e-20, 2.243072e-20, 
    -1.705459e-20, 1.689516e-20, -2.689477e-20, 2.071059e-20, 3.549317e-20, 
    1.565057e-20, 6.031494e-21, 1.322904e-21, -1.462143e-20, 3.212954e-20, 
    -4.842911e-21, -2.580909e-20, 2.75805e-21, 3.782662e-21, -1.538637e-21, 
    8.285423e-21, -1.256174e-20, 2.033824e-20, -4.522845e-21, 6.850294e-21, 
    7.95832e-21, -1.749228e-20, 5.906801e-21, -2.199503e-20, -2.934603e-20, 
    1.004713e-20, -4.740547e-21, 4.07246e-21, 1.139321e-20, -5.784737e-22, 
    1.085092e-20, -5.448506e-21, 1.958022e-20, 4.611191e-22, -1.017801e-20, 
    -4.129819e-20, 1.702944e-20, -4.401949e-20, 2.24084e-20, -1.171947e-20, 
    1.590357e-21, -1.079042e-20, -1.811373e-20, -2.099673e-20, -1.80309e-20, 
    -2.202191e-20, 1.338277e-20, 4.027223e-21, 3.343998e-20, 2.7726e-20, 
    -3.4278e-20, -9.754062e-22, 1.142486e-20, 1.724235e-20, 2.058759e-20, 
    -2.358823e-20, 3.565263e-20, -2.671855e-22, -4.213246e-21, 1.226928e-22, 
    5.884193e-21, -1.698166e-20, -2.092745e-20, 4.23502e-21, -1.366354e-20, 
    -2.44036e-20, -5.122912e-20, -5.218872e-20, 1.184274e-20, 1.450137e-21, 
    -1.847194e-20, 1.011637e-20, -2.955556e-20, 4.132393e-20, 1.955025e-20, 
    2.381895e-20, -4.55745e-20, -4.333584e-20, 2.492724e-20, 2.880406e-20, 
    -9.85514e-21, -1.612245e-20, -1.541392e-20, -1.558157e-20, -1.603395e-20, 
    1.39929e-20, 2.739784e-22, -1.43565e-20, -1.012855e-20, 5.520025e-21, 
    2.15011e-20, 2.32676e-20, 1.29601e-20, -3.487596e-20, 2.824962e-20, 
    -1.617134e-20, -3.39721e-20, 3.500575e-20, -4.207175e-20, 2.730752e-20, 
    -4.496777e-20, -1.921382e-20, -3.029769e-20, -2.534172e-20, 1.040535e-20, 
    3.144759e-20, 1.092303e-20, -4.019858e-21, 3.747991e-20, 1.666727e-20, 
    -2.216298e-20, -1.282579e-20, 4.002873e-20, -2.180559e-20, 1.555338e-23, 
    -3.695828e-20, -3.933633e-20, -3.073369e-20, 2.611895e-20, 3.619219e-21, 
    2.119181e-20, -1.130413e-20, -2.875231e-20, 3.267812e-21, -6.002094e-21, 
    -3.246314e-20, -5.802485e-21, 1.248534e-21 ;

 M_SOIL3C_TO_LEACHING =
  1.111669e-20, 2.599314e-20, -2.170723e-20, 4.078397e-21, -1.698166e-20, 
    -4.472237e-20, 1.115316e-20, 6.433877e-20, -2.399339e-20, -5.329485e-22, 
    -3.427322e-20, -2.209769e-20, 5.136367e-21, 1.557338e-20, 4.8708e-20, 
    -2.834434e-20, -5.376676e-21, -1.074264e-20, 4.775906e-21, 9.066329e-21, 
    -5.195184e-21, 2.021487e-22, -1.882365e-20, 1.204311e-22, -9.605214e-21, 
    -4.907931e-21, -3.809967e-20, -1.556547e-20, 7.18449e-21, 3.853903e-21, 
    -7.546096e-21, -1.135701e-20, 1.304126e-20, -8.937122e-21, 3.434314e-21, 
    6.061576e-22, -1.904644e-20, -1.512693e-20, 1.963624e-20, 4.312508e-21, 
    1.624883e-20, 1.673822e-20, 4.867754e-21, -1.764522e-20, -1.975497e-20, 
    -1.719341e-20, -4.170534e-20, -6.808208e-22, -4.300067e-21, 8.864181e-21, 
    -2.984779e-21, -3.151374e-20, -1.103695e-20, 1.905058e-21, -3.257051e-21, 
    -2.425547e-20, -4.20435e-20, 1.873668e-21, 2.936669e-20, 4.460348e-21, 
    2.978908e-20, -2.061107e-20, 9.689201e-21, 2.130771e-20, 1.128858e-20, 
    1.641676e-20, 1.695282e-20, -3.274221e-20, 2.078129e-20, -5.67722e-21, 
    6.99645e-21, 7.626097e-21, -1.470143e-20, 4.793641e-20, -1.358126e-20, 
    2.075158e-20, 1.650074e-20, 2.217174e-20, 6.789509e-21, -1.171496e-20, 
    -2.795754e-20, 7.04563e-22, 1.263495e-20, -3.76483e-21, 3.70233e-20, 
    -3.327063e-20, 6.231381e-21, -1.82254e-20, 2.693776e-20, -6.615456e-23, 
    -8.247417e-22, -1.194537e-20, -2.156096e-21, -3.107748e-20, 
    -2.122574e-20, 3.255934e-21, -4.612768e-21, 2.673815e-20, 1.421316e-20, 
    -5.407211e-21, 9.499471e-21, 1.341898e-20, -3.429639e-20, 1.941935e-20, 
    -2.463376e-20, 2.552975e-20, -1.37246e-20, 2.598863e-20, 6.294737e-21, 
    8.736538e-22, 1.555338e-23, 7.811003e-21, 2.873645e-20, 1.287273e-20, 
    5.108935e-21, -1.316735e-20, -1.590332e-20, -1.787651e-20, 6.177955e-21, 
    -1.785784e-20, 1.30107e-20, -6.093134e-21, -1.134882e-20, -1.895258e-20, 
    1.011356e-20, 1.37178e-20, -3.213125e-20, -4.628043e-21, -5.705224e-21, 
    -2.702041e-21, -2.791178e-20, -1.548488e-20, -7.08749e-21, -7.451658e-21, 
    -3.521696e-21, 1.864335e-21, 6.763767e-21, 1.330163e-20, -2.213585e-20, 
    -1.476164e-20, 3.490735e-20, 3.422737e-20, 1.610547e-20, -1.710096e-20, 
    -7.526312e-21, 1.182947e-20, -4.716092e-20, -1.402092e-20, 6.405819e-21, 
    -4.664804e-20, -2.487578e-20, 9.620195e-21, 7.5048e-21, -9.224669e-21, 
    3.490538e-20, 1.280064e-20, 3.177873e-22, 5.516939e-21, -1.508648e-21, 
    -1.05925e-20, -5.214885e-20, -2.626881e-20, -1.717296e-21, -2.782552e-20, 
    -2.118784e-20, -2.420544e-20, 1.342689e-20, 9.162735e-21, -3.508379e-20, 
    8.515876e-21, -1.14448e-21, 2.530453e-21, 3.221169e-21, -4.329457e-21, 
    -1.978211e-20, 1.779029e-20, -3.085356e-20, 6.750492e-21, 4.086586e-21, 
    7.7471e-21, -1.441759e-20, 1.077318e-20, -1.605402e-20, 2.311465e-20, 
    -1.728106e-20, 2.216525e-20, -6.329786e-21, -1.060748e-20, 2.517094e-20, 
    -3.693511e-20, -4.990179e-22, -3.563341e-20, 6.510445e-21, -1.77702e-20, 
    -1.025607e-20, 1.697938e-20, 8.973582e-21, 1.278566e-20, 2.728061e-21, 
    -3.101586e-20, 3.324999e-20, 3.876465e-20, -3.18355e-20, 1.572492e-20, 
    -7.284274e-21, -2.126157e-22, 4.253767e-20, 2.816823e-21, 1.466524e-20, 
    2.076374e-20, -1.419025e-20, -3.112414e-20, 2.931775e-20, -2.803813e-20, 
    1.684565e-20, -1.512102e-20, -2.017256e-20, -2.126672e-20, -1.852456e-21, 
    -7.878864e-21, 5.233655e-21, 1.533618e-20, 2.535331e-20, 2.113723e-20, 
    3.050213e-20, 1.075197e-20, -7.072509e-21, 7.626097e-21, 6.672695e-23, 
    -5.992477e-21, 4.500508e-20, 2.103941e-20, 7.5427e-21, -1.660055e-20, 
    -1.043022e-20, 2.044766e-20, 2.806554e-20, -7.991923e-21, 1.229567e-20, 
    4.564402e-21, -6.279576e-22, 9.971351e-21, -9.901088e-22, -1.168922e-20, 
    1.527736e-20, 7.44769e-21, -2.084005e-21, 1.957289e-20, -1.163947e-20, 
    -1.264659e-21, -1.679054e-20, -9.345672e-21, 2.100352e-20, 1.741339e-20, 
    -9.952973e-21, 1.235619e-20, -9.341598e-22, -7.506503e-22, 1.043841e-20, 
    -7.436384e-20, -9.466968e-21, 1.556207e-20, 1.195555e-20, 1.700173e-20, 
    1.050656e-20, -5.224011e-21, -1.229483e-20, 9.105624e-21, -1.430532e-20, 
    -1.204123e-20, 2.172502e-20, 1.918217e-20, -5.639632e-21, -3.594272e-20, 
    -1.341925e-20, 2.389929e-21, -1.616709e-20, 1.443992e-20, -2.41175e-20, 
    1.843717e-20, -3.117389e-20, -1.816094e-20, -1.091314e-20, 1.013251e-20, 
    2.760273e-20, 3.101812e-20, -2.008124e-20, 2.066111e-20, -1.187667e-20, 
    -2.475789e-20, -2.03196e-20, 5.239565e-21, 2.501315e-21, -7.637136e-21, 
    4.415133e-21, -7.710083e-21, 2.548222e-20, -1.274379e-20, 8.250348e-21, 
    -1.742073e-20, 3.855118e-20, 7.183355e-21, -8.643916e-21, -2.003543e-20, 
    -8.063752e-21, 1.371799e-21, 3.093218e-20, 1.640916e-20, -2.661685e-20, 
    -2.804493e-20, -2.246497e-20, -4.354139e-20, 2.872009e-20, 1.72723e-20, 
    -1.392309e-20, -1.194399e-20, 3.018432e-20, 8.773418e-21, -4.610489e-21, 
    6.597517e-21, 7.378104e-23, 1.255326e-20, 9.947037e-21, 8.780766e-21, 
    1.181337e-20, -1.69039e-20, -2.534343e-20, -1.041101e-20, 2.085281e-20, 
    -2.569231e-20, -2.052935e-20, 2.668131e-20, 7.628638e-21, 1.774249e-20, 
    -3.208145e-20, -3.945515e-21, -1.665877e-20, -2.58023e-20 ;

 NBP =
  -6.191079e-08, -6.218382e-08, -6.213074e-08, -6.235096e-08, -6.22288e-08, 
    -6.2373e-08, -6.196615e-08, -6.219464e-08, -6.204878e-08, -6.193537e-08, 
    -6.277832e-08, -6.236078e-08, -6.321213e-08, -6.294581e-08, 
    -6.361488e-08, -6.317068e-08, -6.370446e-08, -6.360209e-08, 
    -6.391026e-08, -6.382197e-08, -6.421612e-08, -6.395101e-08, 
    -6.442048e-08, -6.415281e-08, -6.419468e-08, -6.394226e-08, 
    -6.244482e-08, -6.272633e-08, -6.242814e-08, -6.246828e-08, 
    -6.245027e-08, -6.223132e-08, -6.212098e-08, -6.188993e-08, 
    -6.193188e-08, -6.210158e-08, -6.248633e-08, -6.235573e-08, 
    -6.268491e-08, -6.267748e-08, -6.304396e-08, -6.287872e-08, 
    -6.349475e-08, -6.331966e-08, -6.382565e-08, -6.369839e-08, 
    -6.381968e-08, -6.378291e-08, -6.382015e-08, -6.363351e-08, 
    -6.371348e-08, -6.354926e-08, -6.290966e-08, -6.309762e-08, 
    -6.253705e-08, -6.219999e-08, -6.197617e-08, -6.181733e-08, 
    -6.183978e-08, -6.188259e-08, -6.210257e-08, -6.230942e-08, 
    -6.246706e-08, -6.25725e-08, -6.267641e-08, -6.299089e-08, -6.315737e-08, 
    -6.353015e-08, -6.346289e-08, -6.357685e-08, -6.368574e-08, 
    -6.386854e-08, -6.383846e-08, -6.391899e-08, -6.357385e-08, 
    -6.380323e-08, -6.342457e-08, -6.352813e-08, -6.270461e-08, 
    -6.239097e-08, -6.225762e-08, -6.214094e-08, -6.185705e-08, -6.20531e-08, 
    -6.197581e-08, -6.215969e-08, -6.227652e-08, -6.221874e-08, 
    -6.257539e-08, -6.243673e-08, -6.316724e-08, -6.285257e-08, 
    -6.367303e-08, -6.34767e-08, -6.37201e-08, -6.35959e-08, -6.380871e-08, 
    -6.361718e-08, -6.394897e-08, -6.402121e-08, -6.397185e-08, 
    -6.416151e-08, -6.360656e-08, -6.381967e-08, -6.221712e-08, 
    -6.222654e-08, -6.227045e-08, -6.207744e-08, -6.206563e-08, 
    -6.188878e-08, -6.204615e-08, -6.211316e-08, -6.22833e-08, -6.238393e-08, 
    -6.247959e-08, -6.268994e-08, -6.292485e-08, -6.325337e-08, 
    -6.348942e-08, -6.364765e-08, -6.355063e-08, -6.363629e-08, 
    -6.354053e-08, -6.349565e-08, -6.399414e-08, -6.371423e-08, 
    -6.413423e-08, -6.411099e-08, -6.392091e-08, -6.411361e-08, 
    -6.223316e-08, -6.217893e-08, -6.199063e-08, -6.213799e-08, 
    -6.186952e-08, -6.201979e-08, -6.210619e-08, -6.243962e-08, 
    -6.251289e-08, -6.258082e-08, -6.271499e-08, -6.288717e-08, 
    -6.318925e-08, -6.34521e-08, -6.369208e-08, -6.367449e-08, -6.368068e-08, 
    -6.373428e-08, -6.36015e-08, -6.375608e-08, -6.378202e-08, -6.37142e-08, 
    -6.410788e-08, -6.39954e-08, -6.411049e-08, -6.403727e-08, -6.219656e-08, 
    -6.228781e-08, -6.22385e-08, -6.233122e-08, -6.22659e-08, -6.255637e-08, 
    -6.264347e-08, -6.305104e-08, -6.288379e-08, -6.315e-08, -6.291083e-08, 
    -6.295321e-08, -6.315866e-08, -6.292376e-08, -6.34376e-08, -6.30892e-08, 
    -6.373637e-08, -6.338842e-08, -6.375817e-08, -6.369104e-08, -6.38022e-08, 
    -6.390175e-08, -6.402701e-08, -6.425812e-08, -6.420461e-08, -6.43979e-08, 
    -6.242386e-08, -6.254222e-08, -6.253181e-08, -6.265568e-08, -6.27473e-08, 
    -6.294588e-08, -6.326439e-08, -6.314462e-08, -6.336451e-08, 
    -6.340865e-08, -6.307459e-08, -6.327969e-08, -6.262145e-08, 
    -6.272778e-08, -6.266447e-08, -6.243319e-08, -6.31722e-08, -6.279292e-08, 
    -6.349332e-08, -6.328784e-08, -6.388755e-08, -6.358929e-08, 
    -6.417515e-08, -6.442559e-08, -6.466136e-08, -6.493683e-08, 
    -6.260683e-08, -6.25264e-08, -6.267042e-08, -6.286966e-08, -6.305456e-08, 
    -6.330037e-08, -6.332552e-08, -6.337157e-08, -6.349087e-08, 
    -6.359117e-08, -6.338612e-08, -6.361631e-08, -6.275242e-08, 
    -6.320513e-08, -6.249599e-08, -6.27095e-08, -6.285792e-08, -6.279282e-08, 
    -6.313093e-08, -6.321061e-08, -6.353445e-08, -6.336705e-08, 
    -6.436377e-08, -6.392277e-08, -6.514664e-08, -6.480458e-08, -6.24983e-08, 
    -6.260656e-08, -6.298333e-08, -6.280406e-08, -6.331678e-08, -6.3443e-08, 
    -6.354561e-08, -6.367676e-08, -6.369093e-08, -6.376864e-08, 
    -6.364129e-08, -6.376361e-08, -6.33009e-08, -6.350767e-08, -6.294027e-08, 
    -6.307836e-08, -6.301484e-08, -6.294515e-08, -6.316022e-08, 
    -6.338935e-08, -6.339426e-08, -6.346773e-08, -6.367474e-08, 
    -6.331886e-08, -6.442066e-08, -6.374017e-08, -6.272461e-08, 
    -6.293312e-08, -6.296292e-08, -6.288214e-08, -6.343034e-08, -6.32317e-08, 
    -6.376674e-08, -6.362214e-08, -6.385908e-08, -6.374134e-08, 
    -6.372401e-08, -6.35728e-08, -6.347865e-08, -6.32408e-08, -6.30473e-08, 
    -6.289386e-08, -6.292954e-08, -6.309808e-08, -6.340337e-08, -6.36922e-08, 
    -6.362893e-08, -6.384107e-08, -6.327961e-08, -6.351502e-08, 
    -6.342403e-08, -6.36613e-08, -6.314143e-08, -6.358408e-08, -6.302828e-08, 
    -6.307702e-08, -6.322776e-08, -6.353098e-08, -6.359809e-08, 
    -6.366972e-08, -6.362552e-08, -6.341112e-08, -6.337601e-08, 
    -6.322409e-08, -6.318215e-08, -6.306641e-08, -6.297058e-08, 
    -6.305813e-08, -6.315008e-08, -6.341122e-08, -6.364657e-08, 
    -6.390317e-08, -6.396598e-08, -6.426577e-08, -6.402171e-08, 
    -6.442445e-08, -6.408201e-08, -6.467483e-08, -6.360975e-08, 
    -6.407196e-08, -6.323462e-08, -6.332483e-08, -6.348797e-08, 
    -6.386221e-08, -6.366019e-08, -6.389647e-08, -6.337463e-08, 
    -6.310389e-08, -6.303387e-08, -6.290318e-08, -6.303685e-08, 
    -6.302598e-08, -6.315389e-08, -6.311279e-08, -6.341989e-08, 
    -6.325493e-08, -6.372358e-08, -6.38946e-08, -6.437764e-08, -6.467376e-08, 
    -6.497525e-08, -6.510835e-08, -6.514885e-08, -6.516579e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.191079e-08, 6.218382e-08, 6.213074e-08, 6.235096e-08, 6.22288e-08, 
    6.2373e-08, 6.196615e-08, 6.219464e-08, 6.204878e-08, 6.193537e-08, 
    6.277832e-08, 6.236078e-08, 6.321213e-08, 6.294581e-08, 6.361488e-08, 
    6.317068e-08, 6.370446e-08, 6.360209e-08, 6.391026e-08, 6.382197e-08, 
    6.421612e-08, 6.395101e-08, 6.442048e-08, 6.415281e-08, 6.419468e-08, 
    6.394226e-08, 6.244482e-08, 6.272633e-08, 6.242814e-08, 6.246828e-08, 
    6.245027e-08, 6.223132e-08, 6.212098e-08, 6.188993e-08, 6.193188e-08, 
    6.210158e-08, 6.248633e-08, 6.235573e-08, 6.268491e-08, 6.267748e-08, 
    6.304396e-08, 6.287872e-08, 6.349475e-08, 6.331966e-08, 6.382565e-08, 
    6.369839e-08, 6.381968e-08, 6.378291e-08, 6.382015e-08, 6.363351e-08, 
    6.371348e-08, 6.354926e-08, 6.290966e-08, 6.309762e-08, 6.253705e-08, 
    6.219999e-08, 6.197617e-08, 6.181733e-08, 6.183978e-08, 6.188259e-08, 
    6.210257e-08, 6.230942e-08, 6.246706e-08, 6.25725e-08, 6.267641e-08, 
    6.299089e-08, 6.315737e-08, 6.353015e-08, 6.346289e-08, 6.357685e-08, 
    6.368574e-08, 6.386854e-08, 6.383846e-08, 6.391899e-08, 6.357385e-08, 
    6.380323e-08, 6.342457e-08, 6.352813e-08, 6.270461e-08, 6.239097e-08, 
    6.225762e-08, 6.214094e-08, 6.185705e-08, 6.20531e-08, 6.197581e-08, 
    6.215969e-08, 6.227652e-08, 6.221874e-08, 6.257539e-08, 6.243673e-08, 
    6.316724e-08, 6.285257e-08, 6.367303e-08, 6.34767e-08, 6.37201e-08, 
    6.35959e-08, 6.380871e-08, 6.361718e-08, 6.394897e-08, 6.402121e-08, 
    6.397185e-08, 6.416151e-08, 6.360656e-08, 6.381967e-08, 6.221712e-08, 
    6.222654e-08, 6.227045e-08, 6.207744e-08, 6.206563e-08, 6.188878e-08, 
    6.204615e-08, 6.211316e-08, 6.22833e-08, 6.238393e-08, 6.247959e-08, 
    6.268994e-08, 6.292485e-08, 6.325337e-08, 6.348942e-08, 6.364765e-08, 
    6.355063e-08, 6.363629e-08, 6.354053e-08, 6.349565e-08, 6.399414e-08, 
    6.371423e-08, 6.413423e-08, 6.411099e-08, 6.392091e-08, 6.411361e-08, 
    6.223316e-08, 6.217893e-08, 6.199063e-08, 6.213799e-08, 6.186952e-08, 
    6.201979e-08, 6.210619e-08, 6.243962e-08, 6.251289e-08, 6.258082e-08, 
    6.271499e-08, 6.288717e-08, 6.318925e-08, 6.34521e-08, 6.369208e-08, 
    6.367449e-08, 6.368068e-08, 6.373428e-08, 6.36015e-08, 6.375608e-08, 
    6.378202e-08, 6.37142e-08, 6.410788e-08, 6.39954e-08, 6.411049e-08, 
    6.403727e-08, 6.219656e-08, 6.228781e-08, 6.22385e-08, 6.233122e-08, 
    6.22659e-08, 6.255637e-08, 6.264347e-08, 6.305104e-08, 6.288379e-08, 
    6.315e-08, 6.291083e-08, 6.295321e-08, 6.315866e-08, 6.292376e-08, 
    6.34376e-08, 6.30892e-08, 6.373637e-08, 6.338842e-08, 6.375817e-08, 
    6.369104e-08, 6.38022e-08, 6.390175e-08, 6.402701e-08, 6.425812e-08, 
    6.420461e-08, 6.43979e-08, 6.242386e-08, 6.254222e-08, 6.253181e-08, 
    6.265568e-08, 6.27473e-08, 6.294588e-08, 6.326439e-08, 6.314462e-08, 
    6.336451e-08, 6.340865e-08, 6.307459e-08, 6.327969e-08, 6.262145e-08, 
    6.272778e-08, 6.266447e-08, 6.243319e-08, 6.31722e-08, 6.279292e-08, 
    6.349332e-08, 6.328784e-08, 6.388755e-08, 6.358929e-08, 6.417515e-08, 
    6.442559e-08, 6.466136e-08, 6.493683e-08, 6.260683e-08, 6.25264e-08, 
    6.267042e-08, 6.286966e-08, 6.305456e-08, 6.330037e-08, 6.332552e-08, 
    6.337157e-08, 6.349087e-08, 6.359117e-08, 6.338612e-08, 6.361631e-08, 
    6.275242e-08, 6.320513e-08, 6.249599e-08, 6.27095e-08, 6.285792e-08, 
    6.279282e-08, 6.313093e-08, 6.321061e-08, 6.353445e-08, 6.336705e-08, 
    6.436377e-08, 6.392277e-08, 6.514664e-08, 6.480458e-08, 6.24983e-08, 
    6.260656e-08, 6.298333e-08, 6.280406e-08, 6.331678e-08, 6.3443e-08, 
    6.354561e-08, 6.367676e-08, 6.369093e-08, 6.376864e-08, 6.364129e-08, 
    6.376361e-08, 6.33009e-08, 6.350767e-08, 6.294027e-08, 6.307836e-08, 
    6.301484e-08, 6.294515e-08, 6.316022e-08, 6.338935e-08, 6.339426e-08, 
    6.346773e-08, 6.367474e-08, 6.331886e-08, 6.442066e-08, 6.374017e-08, 
    6.272461e-08, 6.293312e-08, 6.296292e-08, 6.288214e-08, 6.343034e-08, 
    6.32317e-08, 6.376674e-08, 6.362214e-08, 6.385908e-08, 6.374134e-08, 
    6.372401e-08, 6.35728e-08, 6.347865e-08, 6.32408e-08, 6.30473e-08, 
    6.289386e-08, 6.292954e-08, 6.309808e-08, 6.340337e-08, 6.36922e-08, 
    6.362893e-08, 6.384107e-08, 6.327961e-08, 6.351502e-08, 6.342403e-08, 
    6.36613e-08, 6.314143e-08, 6.358408e-08, 6.302828e-08, 6.307702e-08, 
    6.322776e-08, 6.353098e-08, 6.359809e-08, 6.366972e-08, 6.362552e-08, 
    6.341112e-08, 6.337601e-08, 6.322409e-08, 6.318215e-08, 6.306641e-08, 
    6.297058e-08, 6.305813e-08, 6.315008e-08, 6.341122e-08, 6.364657e-08, 
    6.390317e-08, 6.396598e-08, 6.426577e-08, 6.402171e-08, 6.442445e-08, 
    6.408201e-08, 6.467483e-08, 6.360975e-08, 6.407196e-08, 6.323462e-08, 
    6.332483e-08, 6.348797e-08, 6.386221e-08, 6.366019e-08, 6.389647e-08, 
    6.337463e-08, 6.310389e-08, 6.303387e-08, 6.290318e-08, 6.303685e-08, 
    6.302598e-08, 6.315389e-08, 6.311279e-08, 6.341989e-08, 6.325493e-08, 
    6.372358e-08, 6.38946e-08, 6.437764e-08, 6.467376e-08, 6.497525e-08, 
    6.510835e-08, 6.514885e-08, 6.516579e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.191079e-08, -6.218382e-08, -6.213074e-08, -6.235096e-08, -6.22288e-08, 
    -6.2373e-08, -6.196615e-08, -6.219464e-08, -6.204878e-08, -6.193537e-08, 
    -6.277832e-08, -6.236078e-08, -6.321213e-08, -6.294581e-08, 
    -6.361488e-08, -6.317068e-08, -6.370446e-08, -6.360209e-08, 
    -6.391026e-08, -6.382197e-08, -6.421612e-08, -6.395101e-08, 
    -6.442048e-08, -6.415281e-08, -6.419468e-08, -6.394226e-08, 
    -6.244482e-08, -6.272633e-08, -6.242814e-08, -6.246828e-08, 
    -6.245027e-08, -6.223132e-08, -6.212098e-08, -6.188993e-08, 
    -6.193188e-08, -6.210158e-08, -6.248633e-08, -6.235573e-08, 
    -6.268491e-08, -6.267748e-08, -6.304396e-08, -6.287872e-08, 
    -6.349475e-08, -6.331966e-08, -6.382565e-08, -6.369839e-08, 
    -6.381968e-08, -6.378291e-08, -6.382015e-08, -6.363351e-08, 
    -6.371348e-08, -6.354926e-08, -6.290966e-08, -6.309762e-08, 
    -6.253705e-08, -6.219999e-08, -6.197617e-08, -6.181733e-08, 
    -6.183978e-08, -6.188259e-08, -6.210257e-08, -6.230942e-08, 
    -6.246706e-08, -6.25725e-08, -6.267641e-08, -6.299089e-08, -6.315737e-08, 
    -6.353015e-08, -6.346289e-08, -6.357685e-08, -6.368574e-08, 
    -6.386854e-08, -6.383846e-08, -6.391899e-08, -6.357385e-08, 
    -6.380323e-08, -6.342457e-08, -6.352813e-08, -6.270461e-08, 
    -6.239097e-08, -6.225762e-08, -6.214094e-08, -6.185705e-08, -6.20531e-08, 
    -6.197581e-08, -6.215969e-08, -6.227652e-08, -6.221874e-08, 
    -6.257539e-08, -6.243673e-08, -6.316724e-08, -6.285257e-08, 
    -6.367303e-08, -6.34767e-08, -6.37201e-08, -6.35959e-08, -6.380871e-08, 
    -6.361718e-08, -6.394897e-08, -6.402121e-08, -6.397185e-08, 
    -6.416151e-08, -6.360656e-08, -6.381967e-08, -6.221712e-08, 
    -6.222654e-08, -6.227045e-08, -6.207744e-08, -6.206563e-08, 
    -6.188878e-08, -6.204615e-08, -6.211316e-08, -6.22833e-08, -6.238393e-08, 
    -6.247959e-08, -6.268994e-08, -6.292485e-08, -6.325337e-08, 
    -6.348942e-08, -6.364765e-08, -6.355063e-08, -6.363629e-08, 
    -6.354053e-08, -6.349565e-08, -6.399414e-08, -6.371423e-08, 
    -6.413423e-08, -6.411099e-08, -6.392091e-08, -6.411361e-08, 
    -6.223316e-08, -6.217893e-08, -6.199063e-08, -6.213799e-08, 
    -6.186952e-08, -6.201979e-08, -6.210619e-08, -6.243962e-08, 
    -6.251289e-08, -6.258082e-08, -6.271499e-08, -6.288717e-08, 
    -6.318925e-08, -6.34521e-08, -6.369208e-08, -6.367449e-08, -6.368068e-08, 
    -6.373428e-08, -6.36015e-08, -6.375608e-08, -6.378202e-08, -6.37142e-08, 
    -6.410788e-08, -6.39954e-08, -6.411049e-08, -6.403727e-08, -6.219656e-08, 
    -6.228781e-08, -6.22385e-08, -6.233122e-08, -6.22659e-08, -6.255637e-08, 
    -6.264347e-08, -6.305104e-08, -6.288379e-08, -6.315e-08, -6.291083e-08, 
    -6.295321e-08, -6.315866e-08, -6.292376e-08, -6.34376e-08, -6.30892e-08, 
    -6.373637e-08, -6.338842e-08, -6.375817e-08, -6.369104e-08, -6.38022e-08, 
    -6.390175e-08, -6.402701e-08, -6.425812e-08, -6.420461e-08, -6.43979e-08, 
    -6.242386e-08, -6.254222e-08, -6.253181e-08, -6.265568e-08, -6.27473e-08, 
    -6.294588e-08, -6.326439e-08, -6.314462e-08, -6.336451e-08, 
    -6.340865e-08, -6.307459e-08, -6.327969e-08, -6.262145e-08, 
    -6.272778e-08, -6.266447e-08, -6.243319e-08, -6.31722e-08, -6.279292e-08, 
    -6.349332e-08, -6.328784e-08, -6.388755e-08, -6.358929e-08, 
    -6.417515e-08, -6.442559e-08, -6.466136e-08, -6.493683e-08, 
    -6.260683e-08, -6.25264e-08, -6.267042e-08, -6.286966e-08, -6.305456e-08, 
    -6.330037e-08, -6.332552e-08, -6.337157e-08, -6.349087e-08, 
    -6.359117e-08, -6.338612e-08, -6.361631e-08, -6.275242e-08, 
    -6.320513e-08, -6.249599e-08, -6.27095e-08, -6.285792e-08, -6.279282e-08, 
    -6.313093e-08, -6.321061e-08, -6.353445e-08, -6.336705e-08, 
    -6.436377e-08, -6.392277e-08, -6.514664e-08, -6.480458e-08, -6.24983e-08, 
    -6.260656e-08, -6.298333e-08, -6.280406e-08, -6.331678e-08, -6.3443e-08, 
    -6.354561e-08, -6.367676e-08, -6.369093e-08, -6.376864e-08, 
    -6.364129e-08, -6.376361e-08, -6.33009e-08, -6.350767e-08, -6.294027e-08, 
    -6.307836e-08, -6.301484e-08, -6.294515e-08, -6.316022e-08, 
    -6.338935e-08, -6.339426e-08, -6.346773e-08, -6.367474e-08, 
    -6.331886e-08, -6.442066e-08, -6.374017e-08, -6.272461e-08, 
    -6.293312e-08, -6.296292e-08, -6.288214e-08, -6.343034e-08, -6.32317e-08, 
    -6.376674e-08, -6.362214e-08, -6.385908e-08, -6.374134e-08, 
    -6.372401e-08, -6.35728e-08, -6.347865e-08, -6.32408e-08, -6.30473e-08, 
    -6.289386e-08, -6.292954e-08, -6.309808e-08, -6.340337e-08, -6.36922e-08, 
    -6.362893e-08, -6.384107e-08, -6.327961e-08, -6.351502e-08, 
    -6.342403e-08, -6.36613e-08, -6.314143e-08, -6.358408e-08, -6.302828e-08, 
    -6.307702e-08, -6.322776e-08, -6.353098e-08, -6.359809e-08, 
    -6.366972e-08, -6.362552e-08, -6.341112e-08, -6.337601e-08, 
    -6.322409e-08, -6.318215e-08, -6.306641e-08, -6.297058e-08, 
    -6.305813e-08, -6.315008e-08, -6.341122e-08, -6.364657e-08, 
    -6.390317e-08, -6.396598e-08, -6.426577e-08, -6.402171e-08, 
    -6.442445e-08, -6.408201e-08, -6.467483e-08, -6.360975e-08, 
    -6.407196e-08, -6.323462e-08, -6.332483e-08, -6.348797e-08, 
    -6.386221e-08, -6.366019e-08, -6.389647e-08, -6.337463e-08, 
    -6.310389e-08, -6.303387e-08, -6.290318e-08, -6.303685e-08, 
    -6.302598e-08, -6.315389e-08, -6.311279e-08, -6.341989e-08, 
    -6.325493e-08, -6.372358e-08, -6.38946e-08, -6.437764e-08, -6.467376e-08, 
    -6.497525e-08, -6.510835e-08, -6.514885e-08, -6.516579e-08 ;

 NET_NMIN =
  8.721729e-09, 8.760189e-09, 8.752712e-09, 8.783733e-09, 8.766526e-09, 
    8.786838e-09, 8.729527e-09, 8.761715e-09, 8.741167e-09, 8.725192e-09, 
    8.843934e-09, 8.785118e-09, 8.905044e-09, 8.867527e-09, 8.961777e-09, 
    8.899205e-09, 8.974395e-09, 8.959975e-09, 9.003385e-09, 8.990948e-09, 
    9.04647e-09, 9.009125e-09, 9.075257e-09, 9.037553e-09, 9.04345e-09, 
    9.007892e-09, 8.796956e-09, 8.836611e-09, 8.794606e-09, 8.80026e-09, 
    8.797723e-09, 8.766881e-09, 8.751337e-09, 8.718791e-09, 8.724699e-09, 
    8.748605e-09, 8.802803e-09, 8.784406e-09, 8.830776e-09, 8.829729e-09, 
    8.881354e-09, 8.858077e-09, 8.944855e-09, 8.920191e-09, 8.991467e-09, 
    8.973541e-09, 8.990625e-09, 8.985445e-09, 8.990693e-09, 8.964402e-09, 
    8.975666e-09, 8.952533e-09, 8.862436e-09, 8.888913e-09, 8.809947e-09, 
    8.762468e-09, 8.730938e-09, 8.708564e-09, 8.711726e-09, 8.717756e-09, 
    8.748745e-09, 8.777882e-09, 8.800089e-09, 8.814943e-09, 8.829579e-09, 
    8.873878e-09, 8.89733e-09, 8.949841e-09, 8.940367e-09, 8.956419e-09, 
    8.971758e-09, 8.997509e-09, 8.99327e-09, 9.004615e-09, 8.955997e-09, 
    8.988308e-09, 8.934969e-09, 8.949557e-09, 8.833551e-09, 8.78937e-09, 
    8.770585e-09, 8.754149e-09, 8.714158e-09, 8.741774e-09, 8.730888e-09, 
    8.75679e-09, 8.773248e-09, 8.765109e-09, 8.815348e-09, 8.795816e-09, 
    8.89872e-09, 8.854394e-09, 8.969969e-09, 8.942311e-09, 8.976598e-09, 
    8.959103e-09, 8.989081e-09, 8.9621e-09, 9.008838e-09, 9.019015e-09, 
    9.01206e-09, 9.038778e-09, 8.960605e-09, 8.990624e-09, 8.76488e-09, 
    8.766207e-09, 8.772393e-09, 8.745205e-09, 8.743541e-09, 8.718628e-09, 
    8.740797e-09, 8.750236e-09, 8.774203e-09, 8.788378e-09, 8.801854e-09, 
    8.831484e-09, 8.864576e-09, 8.910853e-09, 8.944104e-09, 8.966393e-09, 
    8.952726e-09, 8.964792e-09, 8.951304e-09, 8.944982e-09, 9.015201e-09, 
    8.97577e-09, 9.034935e-09, 9.031661e-09, 9.004885e-09, 9.03203e-09, 
    8.76714e-09, 8.759501e-09, 8.732976e-09, 8.753734e-09, 8.715915e-09, 
    8.737083e-09, 8.749255e-09, 8.796222e-09, 8.806544e-09, 8.816112e-09, 
    8.835013e-09, 8.859269e-09, 8.901821e-09, 8.938847e-09, 8.97265e-09, 
    8.970174e-09, 8.971046e-09, 8.978597e-09, 8.959891e-09, 8.981668e-09, 
    8.985322e-09, 8.975767e-09, 9.031223e-09, 9.015379e-09, 9.031591e-09, 
    9.021276e-09, 8.761984e-09, 8.774839e-09, 8.767892e-09, 8.780954e-09, 
    8.771751e-09, 8.812671e-09, 8.824939e-09, 8.882352e-09, 8.858791e-09, 
    8.896291e-09, 8.8626e-09, 8.86857e-09, 8.897511e-09, 8.864421e-09, 
    8.936804e-09, 8.887728e-09, 8.97889e-09, 8.929876e-09, 8.981962e-09, 
    8.972505e-09, 8.988163e-09, 9.002187e-09, 9.019831e-09, 9.052387e-09, 
    9.044848e-09, 9.072076e-09, 8.794003e-09, 8.810676e-09, 8.809209e-09, 
    8.826659e-09, 8.839565e-09, 8.867538e-09, 8.912404e-09, 8.895532e-09, 
    8.926508e-09, 8.932727e-09, 8.885668e-09, 8.914559e-09, 8.821836e-09, 
    8.836815e-09, 8.827898e-09, 8.795317e-09, 8.899419e-09, 8.845991e-09, 
    8.944653e-09, 8.915708e-09, 9.000187e-09, 8.958172e-09, 9.040698e-09, 
    9.075977e-09, 9.109188e-09, 9.147993e-09, 8.819777e-09, 8.808448e-09, 
    8.828735e-09, 8.856801e-09, 8.882847e-09, 8.917473e-09, 8.921017e-09, 
    8.927503e-09, 8.944308e-09, 8.958436e-09, 8.929553e-09, 8.961978e-09, 
    8.840286e-09, 8.904057e-09, 8.804164e-09, 8.83424e-09, 8.855147e-09, 
    8.845977e-09, 8.893605e-09, 8.90483e-09, 8.950447e-09, 8.926865e-09, 
    9.067269e-09, 9.005148e-09, 9.177545e-09, 9.129363e-09, 8.80449e-09, 
    8.819739e-09, 8.872814e-09, 8.84756e-09, 8.919785e-09, 8.937564e-09, 
    8.952018e-09, 8.970493e-09, 8.972489e-09, 8.983435e-09, 8.965497e-09, 
    8.982727e-09, 8.917547e-09, 8.946674e-09, 8.866748e-09, 8.8862e-09, 
    8.877252e-09, 8.867436e-09, 8.897731e-09, 8.930007e-09, 8.930699e-09, 
    8.941049e-09, 8.970209e-09, 8.920078e-09, 9.075283e-09, 8.979425e-09, 
    8.836368e-09, 8.865739e-09, 8.869938e-09, 8.858559e-09, 8.935781e-09, 
    8.9078e-09, 8.983169e-09, 8.962799e-09, 8.996175e-09, 8.97959e-09, 
    8.97715e-09, 8.955849e-09, 8.942586e-09, 8.909082e-09, 8.881823e-09, 
    8.860209e-09, 8.865236e-09, 8.888978e-09, 8.931982e-09, 8.972668e-09, 
    8.963756e-09, 8.993639e-09, 8.914548e-09, 8.94771e-09, 8.934892e-09, 
    8.968316e-09, 8.895084e-09, 8.957437e-09, 8.879145e-09, 8.88601e-09, 
    8.907245e-09, 8.949958e-09, 8.959412e-09, 8.969502e-09, 8.963276e-09, 
    8.933075e-09, 8.928128e-09, 8.906729e-09, 8.90082e-09, 8.884516e-09, 
    8.871017e-09, 8.88335e-09, 8.896301e-09, 8.933088e-09, 8.96624e-09, 
    9.002386e-09, 9.011234e-09, 9.053464e-09, 9.019083e-09, 9.075817e-09, 
    9.027579e-09, 9.111085e-09, 8.961055e-09, 9.026164e-09, 8.908211e-09, 
    8.920918e-09, 8.9439e-09, 8.996617e-09, 8.968159e-09, 9.001441e-09, 
    8.927934e-09, 8.889796e-09, 8.879931e-09, 8.861523e-09, 8.880352e-09, 
    8.878821e-09, 8.896839e-09, 8.891049e-09, 8.934309e-09, 8.911072e-09, 
    8.977088e-09, 9.001179e-09, 9.069222e-09, 9.110935e-09, 9.153403e-09, 
    9.172152e-09, 9.177858e-09, 9.180244e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.006537e-14, 5.020265e-14, 5.017598e-14, 5.028662e-14, 5.022528e-14, 
    5.029769e-14, 5.009324e-14, 5.020808e-14, 5.013479e-14, 5.007777e-14, 
    5.050107e-14, 5.029156e-14, 5.071864e-14, 5.058518e-14, 5.092029e-14, 
    5.069785e-14, 5.096511e-14, 5.091392e-14, 5.106806e-14, 5.102392e-14, 
    5.122079e-14, 5.108843e-14, 5.132283e-14, 5.118922e-14, 5.121011e-14, 
    5.108405e-14, 5.033379e-14, 5.047498e-14, 5.032541e-14, 5.034555e-14, 
    5.033653e-14, 5.022653e-14, 5.017103e-14, 5.005491e-14, 5.007601e-14, 
    5.016131e-14, 5.035461e-14, 5.028905e-14, 5.045433e-14, 5.04506e-14, 
    5.06344e-14, 5.055155e-14, 5.086021e-14, 5.077255e-14, 5.102576e-14, 
    5.096211e-14, 5.102276e-14, 5.100438e-14, 5.1023e-14, 5.092965e-14, 
    5.096965e-14, 5.088749e-14, 5.056706e-14, 5.066128e-14, 5.038009e-14, 
    5.021072e-14, 5.009827e-14, 5.001838e-14, 5.002968e-14, 5.00512e-14, 
    5.016181e-14, 5.026579e-14, 5.034497e-14, 5.039791e-14, 5.045006e-14, 
    5.060771e-14, 5.06912e-14, 5.08779e-14, 5.084426e-14, 5.090128e-14, 
    5.095578e-14, 5.104719e-14, 5.103216e-14, 5.107241e-14, 5.08998e-14, 
    5.101452e-14, 5.082509e-14, 5.087692e-14, 5.046407e-14, 5.030675e-14, 
    5.023969e-14, 5.01811e-14, 5.003836e-14, 5.013694e-14, 5.009808e-14, 
    5.019055e-14, 5.024925e-14, 5.022023e-14, 5.039936e-14, 5.032973e-14, 
    5.069615e-14, 5.053841e-14, 5.094942e-14, 5.085117e-14, 5.097297e-14, 
    5.091084e-14, 5.101727e-14, 5.092149e-14, 5.10874e-14, 5.112348e-14, 
    5.109882e-14, 5.119359e-14, 5.091617e-14, 5.102275e-14, 5.021941e-14, 
    5.022414e-14, 5.024621e-14, 5.014918e-14, 5.014325e-14, 5.005432e-14, 
    5.013346e-14, 5.016714e-14, 5.025267e-14, 5.030321e-14, 5.035125e-14, 
    5.045684e-14, 5.057466e-14, 5.073932e-14, 5.085754e-14, 5.093673e-14, 
    5.088819e-14, 5.093105e-14, 5.088313e-14, 5.086068e-14, 5.110995e-14, 
    5.097001e-14, 5.117996e-14, 5.116836e-14, 5.107336e-14, 5.116967e-14, 
    5.022747e-14, 5.020022e-14, 5.010555e-14, 5.017964e-14, 5.004464e-14, 
    5.01202e-14, 5.016362e-14, 5.033115e-14, 5.036798e-14, 5.040207e-14, 
    5.046942e-14, 5.055579e-14, 5.07072e-14, 5.083885e-14, 5.095896e-14, 
    5.095017e-14, 5.095326e-14, 5.098006e-14, 5.091364e-14, 5.099097e-14, 
    5.100393e-14, 5.097002e-14, 5.11668e-14, 5.111061e-14, 5.116811e-14, 
    5.113153e-14, 5.020908e-14, 5.025493e-14, 5.023015e-14, 5.027673e-14, 
    5.024391e-14, 5.038977e-14, 5.043348e-14, 5.063791e-14, 5.055408e-14, 
    5.068752e-14, 5.056766e-14, 5.058889e-14, 5.06918e-14, 5.057415e-14, 
    5.083156e-14, 5.065702e-14, 5.09811e-14, 5.08069e-14, 5.099201e-14, 
    5.095844e-14, 5.101404e-14, 5.106379e-14, 5.11264e-14, 5.124181e-14, 
    5.12151e-14, 5.131159e-14, 5.032327e-14, 5.038268e-14, 5.037748e-14, 
    5.043966e-14, 5.048562e-14, 5.058524e-14, 5.074485e-14, 5.068486e-14, 
    5.079501e-14, 5.081711e-14, 5.064976e-14, 5.07525e-14, 5.042246e-14, 
    5.047579e-14, 5.044406e-14, 5.032794e-14, 5.069864e-14, 5.050848e-14, 
    5.085949e-14, 5.07566e-14, 5.10567e-14, 5.090749e-14, 5.120039e-14, 
    5.132534e-14, 5.1443e-14, 5.158021e-14, 5.041513e-14, 5.037477e-14, 
    5.044706e-14, 5.054697e-14, 5.063971e-14, 5.076287e-14, 5.077549e-14, 
    5.079854e-14, 5.085828e-14, 5.090847e-14, 5.08058e-14, 5.092105e-14, 
    5.048809e-14, 5.071515e-14, 5.035948e-14, 5.046661e-14, 5.05411e-14, 
    5.050846e-14, 5.0678e-14, 5.071793e-14, 5.088006e-14, 5.079629e-14, 
    5.129449e-14, 5.107426e-14, 5.16847e-14, 5.151434e-14, 5.036066e-14, 
    5.041501e-14, 5.060398e-14, 5.05141e-14, 5.077111e-14, 5.08343e-14, 
    5.088568e-14, 5.095127e-14, 5.095838e-14, 5.099724e-14, 5.093355e-14, 
    5.099473e-14, 5.076314e-14, 5.086668e-14, 5.058243e-14, 5.065164e-14, 
    5.061982e-14, 5.058488e-14, 5.069268e-14, 5.080741e-14, 5.080991e-14, 
    5.084667e-14, 5.095012e-14, 5.077215e-14, 5.132279e-14, 5.098287e-14, 
    5.047425e-14, 5.057878e-14, 5.059377e-14, 5.055328e-14, 5.082796e-14, 
    5.072848e-14, 5.09963e-14, 5.092397e-14, 5.104247e-14, 5.098359e-14, 
    5.097493e-14, 5.089928e-14, 5.085215e-14, 5.073303e-14, 5.063607e-14, 
    5.055916e-14, 5.057705e-14, 5.066152e-14, 5.081443e-14, 5.0959e-14, 
    5.092734e-14, 5.103347e-14, 5.075249e-14, 5.087034e-14, 5.082478e-14, 
    5.094356e-14, 5.068325e-14, 5.090479e-14, 5.062656e-14, 5.065098e-14, 
    5.072651e-14, 5.08783e-14, 5.091194e-14, 5.094775e-14, 5.092566e-14, 
    5.081832e-14, 5.080075e-14, 5.072468e-14, 5.070365e-14, 5.064567e-14, 
    5.059763e-14, 5.064151e-14, 5.068757e-14, 5.081839e-14, 5.093617e-14, 
    5.10645e-14, 5.10959e-14, 5.124555e-14, 5.112367e-14, 5.132467e-14, 
    5.11537e-14, 5.144959e-14, 5.091769e-14, 5.114877e-14, 5.072996e-14, 
    5.077514e-14, 5.085678e-14, 5.104398e-14, 5.0943e-14, 5.106111e-14, 
    5.080007e-14, 5.066441e-14, 5.062935e-14, 5.056382e-14, 5.063085e-14, 
    5.06254e-14, 5.068951e-14, 5.066891e-14, 5.082273e-14, 5.074013e-14, 
    5.09747e-14, 5.106019e-14, 5.130146e-14, 5.144914e-14, 5.15994e-14, 
    5.166566e-14, 5.168583e-14, 5.169425e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.484155e-43, 0, 1.912772e-42, 
    3.629363e-43, 4.945042e-41, 1.242251e-41, 5.060599e-39, 9.290469e-41, 
    9.736725e-38, 1.98011e-39, 3.686572e-39, 8.117582e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.165713e-44, 2.802597e-45, 1.31652e-41, 
    1.734807e-42, 1.19825e-41, 6.695404e-42, 1.207219e-41, 6.067622e-43, 
    2.209848e-42, 1.527415e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.107026e-43, 3.643376e-44, 2.39622e-43, 1.41391e-42, 2.581612e-41, 
    1.610512e-41, 5.664469e-41, 2.284116e-43, 9.242965e-42, 1.961818e-44, 
    1.079e-43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.151867e-42, 
    4.624285e-44, 2.457878e-42, 3.279038e-43, 1.007954e-41, 4.652311e-43, 
    9.005024e-41, 2.726717e-40, 1.280843e-40, 2.25279e-39, 3.909623e-43, 
    1.19839e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    5.605194e-44, 7.637077e-43, 1.555441e-43, 6.347882e-43, 1.317221e-43, 
    6.305843e-44, 1.803401e-40, 2.237874e-42, 1.5001e-39, 1.059208e-39, 
    5.835567e-41, 1.101639e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.082857e-44, 1.566652e-42, 1.178492e-42, 1.303208e-42, 3.085659e-42, 
    3.601337e-43, 4.37065e-42, 6.605721e-42, 2.235071e-42, 1.01087e-39, 
    1.837845e-40, 1.051384e-39, 3.479578e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.382207e-44, 0, 3.190757e-42, 9.809089e-45, 4.519188e-42, 
    1.540027e-42, 9.090223e-42, 4.333936e-41, 2.977451e-40, 9.368527e-39, 
    4.266976e-39, 7.056501e-38, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 
    7.006492e-45, 1.401298e-44, 0, 1.401298e-45, 0, 0, 0, 0, 0, 0, 
    6.025583e-44, 1.401298e-45, 3.474379e-41, 2.942727e-43, 2.759103e-39, 
    1.047586e-37, 2.781373e-36, 1.085173e-34, 0, 0, 0, 0, 0, 2.802597e-45, 
    4.203895e-45, 8.407791e-45, 5.745324e-44, 3.040818e-43, 9.809089e-45, 
    4.582246e-43, 0, 0, 0, 0, 0, 0, 0, 0, 1.191104e-43, 7.006492e-45, 
    4.333622e-38, 6.009609e-41, 1.567935e-33, 1.911503e-35, 0, 0, 0, 0, 
    2.802597e-45, 2.662467e-44, 1.429324e-43, 1.223334e-42, 1.537224e-42, 
    5.338947e-42, 6.880375e-43, 4.926965e-42, 2.802597e-45, 7.707142e-44, 0, 
    0, 0, 0, 0, 9.809089e-45, 1.121039e-44, 3.923636e-44, 1.1869e-42, 
    2.802597e-45, 9.780159e-38, 3.396747e-42, 0, 0, 0, 0, 2.101948e-44, 0, 
    5.179199e-42, 5.044674e-43, 2.225822e-41, 3.454201e-42, 2.617626e-42, 
    2.242078e-43, 4.764415e-44, 1.401298e-45, 0, 0, 0, 0, 1.261169e-44, 
    1.569454e-42, 5.63322e-43, 1.677915e-41, 1.401298e-45, 8.68805e-44, 
    1.821688e-44, 9.52883e-43, 0, 2.704506e-43, 0, 0, 0, 1.121039e-43, 
    3.405155e-43, 1.091612e-42, 5.324934e-43, 1.541428e-44, 8.407791e-45, 0, 
    0, 0, 0, 0, 0, 1.541428e-44, 7.496947e-43, 4.430766e-41, 1.170028e-40, 
    1.048755e-38, 2.749264e-40, 1.032221e-37, 6.868086e-40, 3.346619e-36, 
    4.119817e-43, 5.894758e-40, 1.401298e-45, 2.802597e-45, 5.465064e-44, 
    2.339888e-41, 9.360674e-43, 3.99356e-41, 8.407791e-45, 0, 0, 0, 0, 0, 0, 
    0, 1.821688e-44, 1.401298e-45, 2.599409e-42, 3.878654e-41, 5.282891e-38, 
    3.295288e-36, 1.781647e-34, 9.699692e-34, 1.611632e-33, 1.990581e-33 ;

 POT_F_NIT =
  3.83111e-11, 3.86413e-11, 3.857699e-11, 3.884415e-11, 3.869583e-11, 
    3.887093e-11, 3.837791e-11, 3.86544e-11, 3.847777e-11, 3.834074e-11, 
    3.936533e-11, 3.885606e-11, 3.98981e-11, 3.957057e-11, 4.039603e-11, 
    3.984702e-11, 4.050721e-11, 4.038015e-11, 4.076324e-11, 4.065329e-11, 
    4.114531e-11, 4.081402e-11, 4.140161e-11, 4.106607e-11, 4.111845e-11, 
    4.080309e-11, 3.895832e-11, 3.930177e-11, 3.893801e-11, 3.898688e-11, 
    3.896494e-11, 3.869887e-11, 3.856513e-11, 3.828589e-11, 3.83365e-11, 
    3.854164e-11, 3.900883e-11, 3.884991e-11, 3.925108e-11, 3.9242e-11, 
    3.96911e-11, 3.948828e-11, 4.024715e-11, 4.003069e-11, 4.065787e-11, 
    4.049965e-11, 4.065042e-11, 4.060466e-11, 4.0651e-11, 4.04191e-11, 
    4.051836e-11, 4.031462e-11, 3.952627e-11, 3.975713e-11, 3.907066e-11, 
    3.866087e-11, 3.838999e-11, 3.819836e-11, 3.822542e-11, 3.827702e-11, 
    3.854283e-11, 3.879364e-11, 3.898534e-11, 3.911384e-11, 3.924068e-11, 
    3.962589e-11, 3.983061e-11, 4.029098e-11, 4.02077e-11, 4.034883e-11, 
    4.048392e-11, 4.071124e-11, 4.067378e-11, 4.077408e-11, 4.034509e-11, 
    4.062992e-11, 4.016026e-11, 4.028843e-11, 3.927519e-11, 3.889277e-11, 
    3.873077e-11, 3.85893e-11, 3.824622e-11, 3.848297e-11, 3.838954e-11, 
    3.861199e-11, 3.875368e-11, 3.868356e-11, 3.911736e-11, 3.89484e-11, 
    3.984275e-11, 3.945622e-11, 4.046816e-11, 4.022477e-11, 4.052659e-11, 
    4.037244e-11, 4.063675e-11, 4.039882e-11, 4.081144e-11, 4.090158e-11, 
    4.083996e-11, 4.107691e-11, 4.038562e-11, 4.065036e-11, 3.868163e-11, 
    3.869306e-11, 3.874633e-11, 3.851241e-11, 3.849812e-11, 3.828447e-11, 
    3.847454e-11, 3.855563e-11, 3.87619e-11, 3.888416e-11, 3.900058e-11, 
    3.925719e-11, 3.954482e-11, 3.994888e-11, 4.024052e-11, 4.043663e-11, 
    4.031632e-11, 4.042251e-11, 4.03038e-11, 4.024821e-11, 4.086778e-11, 
    4.051927e-11, 4.104277e-11, 4.101371e-11, 4.077643e-11, 4.101697e-11, 
    3.870107e-11, 3.863531e-11, 3.840744e-11, 3.85857e-11, 3.826124e-11, 
    3.844267e-11, 3.854719e-11, 3.89519e-11, 3.904113e-11, 3.912395e-11, 
    3.928781e-11, 3.949861e-11, 3.986984e-11, 4.019433e-11, 4.049177e-11, 
    4.046993e-11, 4.047761e-11, 4.054419e-11, 4.037935e-11, 4.057128e-11, 
    4.060353e-11, 4.051922e-11, 4.100981e-11, 4.086933e-11, 4.101307e-11, 
    4.092158e-11, 3.865668e-11, 3.876738e-11, 3.870753e-11, 3.88201e-11, 
    3.874076e-11, 3.909415e-11, 3.920043e-11, 3.969977e-11, 3.949445e-11, 
    3.98215e-11, 3.95276e-11, 3.957959e-11, 3.983215e-11, 3.954344e-11, 
    4.017638e-11, 3.974666e-11, 4.054677e-11, 4.011556e-11, 4.057387e-11, 
    4.049044e-11, 4.06286e-11, 4.075255e-11, 4.090877e-11, 4.119784e-11, 
    4.11308e-11, 4.137317e-11, 3.893274e-11, 3.90769e-11, 3.90642e-11, 
    3.921535e-11, 3.932732e-11, 3.957062e-11, 3.996246e-11, 3.981487e-11, 
    4.008604e-11, 4.014059e-11, 3.972869e-11, 3.998131e-11, 3.91735e-11, 
    3.93034e-11, 3.922603e-11, 3.894403e-11, 3.984879e-11, 3.938309e-11, 
    4.024529e-11, 3.999133e-11, 4.073485e-11, 4.036417e-11, 4.109392e-11, 
    4.140795e-11, 4.170469e-11, 4.205282e-11, 3.91557e-11, 3.90576e-11, 
    3.923334e-11, 3.947714e-11, 3.970408e-11, 4.000685e-11, 4.003789e-11, 
    4.009476e-11, 4.024229e-11, 4.036654e-11, 4.011273e-11, 4.039771e-11, 
    3.933354e-11, 3.988936e-11, 3.902048e-11, 3.928104e-11, 3.946269e-11, 
    3.938296e-11, 3.979796e-11, 3.989609e-11, 4.02962e-11, 4.008911e-11, 
    4.13303e-11, 4.077871e-11, 4.231895e-11, 4.188549e-11, 3.902335e-11, 
    3.915535e-11, 3.961657e-11, 3.939677e-11, 4.00271e-11, 4.018305e-11, 
    4.031007e-11, 4.047274e-11, 4.049032e-11, 4.058688e-11, 4.04287e-11, 
    4.058062e-11, 4.000745e-11, 4.026305e-11, 3.956367e-11, 3.973329e-11, 
    3.965521e-11, 3.956964e-11, 3.983401e-11, 4.011666e-11, 4.012272e-11, 
    4.021358e-11, 4.047016e-11, 4.002958e-11, 4.140172e-11, 4.055142e-11, 
    3.929955e-11, 3.955493e-11, 3.95915e-11, 3.949241e-11, 4.016739e-11, 
    3.992212e-11, 4.058453e-11, 4.040494e-11, 4.06994e-11, 4.055293e-11, 
    4.053139e-11, 4.034374e-11, 4.022712e-11, 3.993331e-11, 3.969508e-11, 
    3.950672e-11, 3.955047e-11, 3.975753e-11, 4.013398e-11, 4.049184e-11, 
    4.04133e-11, 4.067692e-11, 3.998112e-11, 4.027211e-11, 4.015949e-11, 
    4.045345e-11, 3.981093e-11, 4.035776e-11, 3.967177e-11, 3.973166e-11, 
    3.991725e-11, 4.029194e-11, 4.03751e-11, 4.046398e-11, 4.040912e-11, 
    4.01436e-11, 4.010018e-11, 3.991271e-11, 3.986101e-11, 3.971858e-11, 
    3.960084e-11, 3.970839e-11, 3.982149e-11, 4.014368e-11, 4.043518e-11, 
    4.075426e-11, 4.083255e-11, 4.120736e-11, 4.090208e-11, 4.140646e-11, 
    4.09774e-11, 4.172163e-11, 4.038958e-11, 4.096494e-11, 3.992571e-11, 
    4.003699e-11, 4.023868e-11, 4.070329e-11, 4.045212e-11, 4.074595e-11, 
    4.009848e-11, 3.976468e-11, 3.967857e-11, 3.951815e-11, 3.968223e-11, 
    3.966888e-11, 3.982619e-11, 3.97756e-11, 4.015439e-11, 3.995068e-11, 
    4.053079e-11, 4.074358e-11, 4.134767e-11, 4.172029e-11, 4.210143e-11, 
    4.227026e-11, 4.232172e-11, 4.234324e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005857516, 0.0005857558, 0.000585755, 0.0005857584, 0.0005857565, 
    0.0005857587, 0.0005857525, 0.0005857559, 0.0005857538, 0.000585752, 
    0.0005857648, 0.0005857585, 0.0005857716, 0.0005857676, 0.0005857779, 
    0.0005857709, 0.0005857793, 0.0005857777, 0.0005857825, 0.0005857812, 
    0.0005857872, 0.0005857832, 0.0005857904, 0.0005857862, 0.0005857869, 
    0.000585783, 0.0005857598, 0.0005857639, 0.0005857596, 0.0005857602, 
    0.0005857599, 0.0005857565, 0.0005857548, 0.0005857513, 0.000585752, 
    0.0005857545, 0.0005857604, 0.0005857585, 0.0005857635, 0.0005857634, 
    0.0005857691, 0.0005857665, 0.0005857761, 0.0005857734, 0.0005857812, 
    0.0005857793, 0.0005857811, 0.0005857805, 0.0005857811, 0.0005857782, 
    0.0005857794, 0.0005857769, 0.000585767, 0.0005857699, 0.0005857612, 
    0.0005857559, 0.0005857526, 0.0005857502, 0.0005857506, 0.0005857512, 
    0.0005857545, 0.0005857578, 0.0005857602, 0.0005857618, 0.0005857634, 
    0.0005857681, 0.0005857708, 0.0005857766, 0.0005857756, 0.0005857773, 
    0.000585779, 0.0005857819, 0.0005857814, 0.0005857826, 0.0005857773, 
    0.0005857808, 0.000585775, 0.0005857766, 0.0005857636, 0.000585759, 
    0.0005857568, 0.0005857552, 0.0005857508, 0.0005857538, 0.0005857526, 
    0.0005857554, 0.0005857573, 0.0005857564, 0.0005857619, 0.0005857597, 
    0.0005857709, 0.0005857661, 0.0005857788, 0.0005857758, 0.0005857795, 
    0.0005857776, 0.0005857809, 0.000585778, 0.0005857832, 0.0005857842, 
    0.0005857834, 0.0005857865, 0.0005857778, 0.0005857811, 0.0005857563, 
    0.0005857565, 0.0005857571, 0.0005857542, 0.000585754, 0.0005857513, 
    0.0005857537, 0.0005857547, 0.0005857574, 0.0005857589, 0.0005857604, 
    0.0005857636, 0.0005857671, 0.0005857723, 0.000585776, 0.0005857784, 
    0.0005857769, 0.0005857783, 0.0005857768, 0.0005857761, 0.0005857838, 
    0.0005857794, 0.000585786, 0.0005857857, 0.0005857827, 0.0005857857, 
    0.0005857566, 0.0005857557, 0.0005857528, 0.0005857551, 0.000585751, 
    0.0005857533, 0.0005857546, 0.0005857597, 0.0005857609, 0.0005857619, 
    0.000585764, 0.0005857666, 0.0005857713, 0.0005857754, 0.0005857791, 
    0.0005857788, 0.000585779, 0.0005857798, 0.0005857777, 0.0005857801, 
    0.0005857805, 0.0005857795, 0.0005857856, 0.0005857839, 0.0005857857, 
    0.0005857846, 0.000585756, 0.0005857574, 0.0005857567, 0.0005857581, 
    0.0005857571, 0.0005857615, 0.0005857628, 0.0005857691, 0.0005857666, 
    0.0005857706, 0.000585767, 0.0005857677, 0.0005857707, 0.0005857672, 
    0.0005857751, 0.0005857697, 0.0005857798, 0.0005857743, 0.0005857801, 
    0.0005857791, 0.0005857809, 0.0005857824, 0.0005857844, 0.0005857879, 
    0.0005857871, 0.0005857901, 0.0005857595, 0.0005857613, 0.0005857612, 
    0.0005857631, 0.0005857645, 0.0005857676, 0.0005857724, 0.0005857706, 
    0.0005857741, 0.0005857747, 0.0005857696, 0.0005857727, 0.0005857626, 
    0.0005857641, 0.0005857632, 0.0005857596, 0.000585771, 0.0005857651, 
    0.000585776, 0.0005857729, 0.0005857822, 0.0005857775, 0.0005857866, 
    0.0005857904, 0.0005857943, 0.0005857985, 0.0005857623, 0.0005857611, 
    0.0005857633, 0.0005857663, 0.0005857692, 0.000585773, 0.0005857734, 
    0.0005857741, 0.000585776, 0.0005857776, 0.0005857743, 0.000585778, 
    0.0005857644, 0.0005857715, 0.0005857606, 0.0005857638, 0.0005857662, 
    0.0005857652, 0.0005857705, 0.0005857717, 0.0005857766, 0.0005857741, 
    0.0005857894, 0.0005857826, 0.0005858019, 0.0005857964, 0.0005857607, 
    0.0005857624, 0.0005857681, 0.0005857653, 0.0005857733, 0.0005857752, 
    0.0005857769, 0.0005857788, 0.0005857791, 0.0005857803, 0.0005857783, 
    0.0005857802, 0.000585773, 0.0005857763, 0.0005857675, 0.0005857696, 
    0.0005857687, 0.0005857676, 0.0005857709, 0.0005857744, 0.0005857745, 
    0.0005857756, 0.0005857786, 0.0005857733, 0.0005857902, 0.0005857796, 
    0.0005857642, 0.0005857673, 0.0005857678, 0.0005857666, 0.0005857751, 
    0.000585772, 0.0005857803, 0.000585778, 0.0005857818, 0.0005857799, 
    0.0005857796, 0.0005857773, 0.0005857758, 0.0005857721, 0.0005857691, 
    0.0005857668, 0.0005857673, 0.0005857699, 0.0005857746, 0.0005857791, 
    0.0005857781, 0.0005857815, 0.0005857727, 0.0005857763, 0.0005857749, 
    0.0005857787, 0.0005857706, 0.0005857772, 0.0005857688, 0.0005857696, 
    0.0005857719, 0.0005857765, 0.0005857777, 0.0005857787, 0.0005857781, 
    0.0005857747, 0.0005857742, 0.0005857719, 0.0005857712, 0.0005857694, 
    0.000585768, 0.0005857693, 0.0005857707, 0.0005857748, 0.0005857784, 
    0.0005857824, 0.0005857834, 0.0005857879, 0.0005857841, 0.0005857903, 
    0.0005857848, 0.0005857943, 0.0005857777, 0.0005857849, 0.000585772, 
    0.0005857734, 0.0005857759, 0.0005857817, 0.0005857786, 0.0005857822, 
    0.0005857742, 0.0005857699, 0.000585769, 0.0005857669, 0.000585769, 
    0.0005857688, 0.0005857708, 0.0005857702, 0.0005857749, 0.0005857723, 
    0.0005857796, 0.0005857822, 0.0005857898, 0.0005857944, 0.0005857992, 
    0.0005858013, 0.000585802, 0.0005858022 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  -2.839813e-07, -2.84087e-07, -2.840669e-07, -2.841511e-07, -2.84105e-07, 
    -2.841597e-07, -2.840035e-07, -2.840906e-07, -2.840354e-07, 
    -2.839918e-07, -2.843121e-07, -2.84155e-07, -2.844815e-07, -2.843805e-07, 
    -2.846356e-07, -2.844648e-07, -2.846702e-07, -2.846323e-07, 
    -2.847502e-07, -2.847165e-07, -2.848637e-07, -2.847657e-07, 
    -2.849423e-07, -2.848412e-07, -2.848564e-07, -2.847623e-07, 
    -2.841882e-07, -2.842921e-07, -2.841817e-07, -2.841966e-07, 
    -2.841902e-07, -2.841054e-07, -2.840616e-07, -2.839743e-07, 
    -2.839904e-07, -2.840551e-07, -2.842033e-07, -2.841541e-07, -2.84281e-07, 
    -2.842782e-07, -2.844184e-07, -2.843552e-07, -2.845912e-07, 
    -2.845246e-07, -2.84718e-07, -2.846692e-07, -2.847154e-07, -2.847016e-07, 
    -2.847156e-07, -2.846441e-07, -2.846747e-07, -2.846122e-07, 
    -2.843667e-07, -2.844386e-07, -2.842233e-07, -2.840912e-07, -2.84007e-07, 
    -2.83946e-07, -2.839546e-07, -2.839708e-07, -2.840555e-07, -2.841362e-07, 
    -2.841972e-07, -2.842377e-07, -2.842777e-07, -2.843951e-07, 
    -2.844605e-07, -2.846039e-07, -2.845794e-07, -2.846219e-07, 
    -2.846644e-07, -2.847339e-07, -2.847226e-07, -2.847529e-07, 
    -2.846218e-07, -2.847085e-07, -2.845651e-07, -2.846042e-07, 
    -2.842834e-07, -2.841676e-07, -2.841138e-07, -2.840706e-07, 
    -2.839612e-07, -2.840365e-07, -2.840067e-07, -2.840786e-07, 
    -2.841235e-07, -2.841015e-07, -2.842388e-07, -2.841853e-07, 
    -2.844643e-07, -2.843443e-07, -2.846595e-07, -2.845845e-07, 
    -2.846776e-07, -2.846304e-07, -2.847108e-07, -2.846384e-07, 
    -2.847646e-07, -2.847914e-07, -2.847729e-07, -2.848455e-07, 
    -2.846343e-07, -2.847149e-07, -2.841007e-07, -2.841042e-07, 
    -2.841214e-07, -2.840458e-07, -2.840414e-07, -2.839736e-07, 
    -2.840344e-07, -2.840599e-07, -2.841265e-07, -2.841649e-07, 
    -2.842016e-07, -2.842824e-07, -2.843719e-07, -2.844981e-07, 
    -2.845893e-07, -2.846501e-07, -2.846132e-07, -2.846458e-07, 
    -2.846091e-07, -2.845922e-07, -2.84781e-07, -2.846747e-07, -2.84835e-07, 
    -2.848264e-07, -2.847534e-07, -2.848274e-07, -2.841068e-07, 
    -2.840862e-07, -2.840128e-07, -2.840702e-07, -2.839663e-07, 
    -2.840238e-07, -2.840565e-07, -2.841853e-07, -2.842147e-07, 
    -2.842404e-07, -2.842924e-07, -2.843584e-07, -2.844737e-07, 
    -2.845745e-07, -2.846671e-07, -2.846604e-07, -2.846627e-07, 
    -2.846828e-07, -2.846323e-07, -2.846912e-07, -2.847006e-07, 
    -2.846753e-07, -2.848252e-07, -2.847825e-07, -2.848262e-07, 
    -2.847985e-07, -2.84093e-07, -2.841279e-07, -2.84109e-07, -2.841443e-07, 
    -2.84119e-07, -2.842299e-07, -2.84263e-07, -2.844198e-07, -2.843568e-07, 
    -2.844584e-07, -2.843676e-07, -2.843834e-07, -2.844595e-07, 
    -2.843728e-07, -2.84568e-07, -2.844338e-07, -2.846836e-07, -2.845479e-07, 
    -2.84692e-07, -2.846667e-07, -2.847091e-07, -2.847465e-07, -2.847944e-07, 
    -2.848811e-07, -2.848613e-07, -2.849346e-07, -2.841804e-07, 
    -2.842251e-07, -2.842221e-07, -2.842696e-07, -2.843044e-07, 
    -2.843812e-07, -2.845029e-07, -2.844575e-07, -2.845419e-07, 
    -2.845585e-07, -2.844308e-07, -2.845083e-07, -2.842557e-07, 
    -2.842955e-07, -2.842725e-07, -2.841833e-07, -2.844666e-07, 
    -2.843207e-07, -2.845906e-07, -2.845121e-07, -2.84741e-07, -2.846263e-07, 
    -2.848501e-07, -2.849428e-07, -2.850344e-07, -2.851359e-07, 
    -2.842505e-07, -2.842201e-07, -2.842755e-07, -2.843504e-07, 
    -2.844225e-07, -2.845167e-07, -2.845269e-07, -2.845442e-07, 
    -2.845903e-07, -2.846285e-07, -2.845487e-07, -2.846382e-07, 
    -2.843028e-07, -2.844797e-07, -2.842076e-07, -2.842883e-07, 
    -2.843464e-07, -2.843219e-07, -2.844526e-07, -2.84483e-07, -2.846058e-07, 
    -2.845429e-07, -2.849191e-07, -2.84753e-07, -2.852163e-07, -2.850867e-07, 
    -2.842092e-07, -2.842509e-07, -2.843946e-07, -2.843264e-07, 
    -2.845235e-07, -2.845715e-07, -2.846113e-07, -2.846604e-07, 
    -2.846665e-07, -2.846957e-07, -2.846477e-07, -2.846942e-07, 
    -2.845169e-07, -2.845964e-07, -2.843793e-07, -2.844317e-07, -2.84408e-07, 
    -2.843812e-07, -2.844637e-07, -2.845498e-07, -2.845532e-07, 
    -2.845805e-07, -2.846544e-07, -2.845244e-07, -2.849376e-07, 
    -2.846801e-07, -2.842962e-07, -2.843744e-07, -2.843875e-07, 
    -2.843569e-07, -2.845666e-07, -2.844906e-07, -2.846952e-07, 
    -2.846404e-07, -2.847306e-07, -2.846857e-07, -2.84679e-07, -2.846215e-07, 
    -2.845852e-07, -2.844938e-07, -2.844196e-07, -2.843615e-07, 
    -2.843752e-07, -2.84439e-07, -2.845554e-07, -2.846663e-07, -2.846418e-07, 
    -2.847238e-07, -2.845092e-07, -2.845985e-07, -2.845635e-07, -2.84655e-07, 
    -2.84456e-07, -2.846207e-07, -2.844131e-07, -2.844317e-07, -2.844891e-07, 
    -2.846035e-07, -2.846311e-07, -2.846578e-07, -2.846417e-07, 
    -2.845586e-07, -2.845457e-07, -2.844881e-07, -2.844713e-07, 
    -2.844278e-07, -2.84391e-07, -2.844242e-07, -2.844588e-07, -2.845593e-07, 
    -2.846488e-07, -2.847468e-07, -2.847713e-07, -2.848813e-07, 
    -2.847896e-07, -2.849387e-07, -2.848087e-07, -2.850351e-07, 
    -2.846326e-07, -2.848081e-07, -2.844922e-07, -2.845267e-07, 
    -2.845874e-07, -2.847297e-07, -2.846546e-07, -2.847432e-07, 
    -2.845454e-07, -2.844404e-07, -2.844152e-07, -2.843648e-07, 
    -2.844163e-07, -2.844122e-07, -2.844614e-07, -2.844456e-07, 
    -2.845627e-07, -2.844999e-07, -2.846784e-07, -2.847428e-07, 
    -2.849263e-07, -2.850373e-07, -2.851526e-07, -2.852025e-07, 
    -2.852179e-07, -2.852242e-07 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  9.441314e-06, 9.466045e-06, 9.461244e-06, 9.481187e-06, 9.470137e-06, 
    9.483187e-06, 9.446343e-06, 9.467012e-06, 9.453825e-06, 9.443563e-06, 
    9.519893e-06, 9.482081e-06, 9.559419e-06, 9.535218e-06, 9.596115e-06, 
    9.555627e-06, 9.604296e-06, 9.594987e-06, 9.623115e-06, 9.615056e-06, 
    9.650985e-06, 9.626836e-06, 9.669698e-06, 9.645238e-06, 9.649047e-06, 
    9.626033e-06, 9.489723e-06, 9.515168e-06, 9.488207e-06, 9.491836e-06, 
    9.490216e-06, 9.470352e-06, 9.460321e-06, 9.439452e-06, 9.443246e-06, 
    9.45859e-06, 9.493468e-06, 9.481648e-06, 9.511528e-06, 9.510853e-06, 
    9.54415e-06, 9.52913e-06, 9.585201e-06, 9.569259e-06, 9.615393e-06, 
    9.603776e-06, 9.61484e-06, 9.61149e-06, 9.614883e-06, 9.59785e-06, 
    9.605144e-06, 9.590175e-06, 9.531935e-06, 9.549022e-06, 9.498082e-06, 
    9.46746e-06, 9.447242e-06, 9.432877e-06, 9.434907e-06, 9.43877e-06, 
    9.458679e-06, 9.477449e-06, 9.491752e-06, 9.501319e-06, 9.510756e-06, 
    9.53925e-06, 9.554435e-06, 9.588407e-06, 9.582306e-06, 9.592668e-06, 
    9.602622e-06, 9.619296e-06, 9.616556e-06, 9.623896e-06, 9.59242e-06, 
    9.613322e-06, 9.578824e-06, 9.58825e-06, 9.513186e-06, 9.484843e-06, 
    9.472691e-06, 9.462162e-06, 9.436466e-06, 9.4542e-06, 9.447204e-06, 
    9.463881e-06, 9.474465e-06, 9.469235e-06, 9.501581e-06, 9.488995e-06, 
    9.555334e-06, 9.526732e-06, 9.601461e-06, 9.583561e-06, 9.605758e-06, 
    9.594435e-06, 9.613829e-06, 9.596375e-06, 9.62664e-06, 9.633221e-06, 
    9.62872e-06, 9.646056e-06, 9.595404e-06, 9.614827e-06, 9.469082e-06, 
    9.469934e-06, 9.47392e-06, 9.456403e-06, 9.45534e-06, 9.439341e-06, 
    9.453588e-06, 9.459647e-06, 9.475089e-06, 9.484203e-06, 9.492879e-06, 
    9.511971e-06, 9.533297e-06, 9.563194e-06, 9.584719e-06, 9.599154e-06, 
    9.590311e-06, 9.598117e-06, 9.589386e-06, 9.5853e-06, 9.630746e-06, 
    9.605204e-06, 9.643562e-06, 9.641443e-06, 9.624066e-06, 9.641682e-06, 
    9.470535e-06, 9.465628e-06, 9.448556e-06, 9.461915e-06, 9.437601e-06, 
    9.451191e-06, 9.458999e-06, 9.489228e-06, 9.495909e-06, 9.502062e-06, 
    9.514254e-06, 9.529898e-06, 9.55736e-06, 9.581305e-06, 9.603207e-06, 
    9.601604e-06, 9.602167e-06, 9.607048e-06, 9.59494e-06, 9.609038e-06, 
    9.611392e-06, 9.605217e-06, 9.641159e-06, 9.630887e-06, 9.641398e-06, 
    9.634712e-06, 9.467226e-06, 9.475491e-06, 9.471022e-06, 9.479417e-06, 
    9.473492e-06, 9.499815e-06, 9.507714e-06, 9.54476e-06, 9.529582e-06, 
    9.553782e-06, 9.53205e-06, 9.535891e-06, 9.554514e-06, 9.533233e-06, 
    9.579958e-06, 9.548217e-06, 9.607238e-06, 9.575447e-06, 9.609229e-06, 
    9.603112e-06, 9.613254e-06, 9.622327e-06, 9.633771e-06, 9.654861e-06, 
    9.649982e-06, 9.667653e-06, 9.487829e-06, 9.498547e-06, 9.497628e-06, 
    9.508868e-06, 9.51718e-06, 9.535242e-06, 9.564212e-06, 9.553321e-06, 
    9.573348e-06, 9.57736e-06, 9.546954e-06, 9.565593e-06, 9.505742e-06, 
    9.515373e-06, 9.509657e-06, 9.488659e-06, 9.555795e-06, 9.521295e-06, 
    9.58507e-06, 9.566354e-06, 9.621029e-06, 9.593794e-06, 9.64729e-06, 
    9.670129e-06, 9.691766e-06, 9.716935e-06, 9.504426e-06, 9.497138e-06, 
    9.510212e-06, 9.528272e-06, 9.545117e-06, 9.56749e-06, 9.569794e-06, 
    9.573982e-06, 9.584862e-06, 9.594002e-06, 9.57528e-06, 9.596296e-06, 
    9.517556e-06, 9.558805e-06, 9.49436e-06, 9.513707e-06, 9.527219e-06, 
    9.521316e-06, 9.552084e-06, 9.559332e-06, 9.588805e-06, 9.57358e-06, 
    9.664466e-06, 9.624207e-06, 9.736204e-06, 9.704834e-06, 9.494586e-06, 
    9.504413e-06, 9.538621e-06, 9.522341e-06, 9.568998e-06, 9.580486e-06, 
    9.589853e-06, 9.601789e-06, 9.603097e-06, 9.610177e-06, 9.598574e-06, 
    9.609728e-06, 9.567538e-06, 9.586385e-06, 9.534739e-06, 9.547282e-06, 
    9.54152e-06, 9.535182e-06, 9.554747e-06, 9.575569e-06, 9.576055e-06, 
    9.582729e-06, 9.601472e-06, 9.569188e-06, 9.66959e-06, 9.607459e-06, 
    9.515133e-06, 9.534033e-06, 9.536784e-06, 9.529451e-06, 9.579333e-06, 
    9.56124e-06, 9.61001e-06, 9.596827e-06, 9.618442e-06, 9.607695e-06, 
    9.606112e-06, 9.592328e-06, 9.583739e-06, 9.562062e-06, 9.544452e-06, 
    9.530519e-06, 9.533762e-06, 9.54907e-06, 9.576853e-06, 9.603197e-06, 
    9.597418e-06, 9.616799e-06, 9.565611e-06, 9.587038e-06, 9.57874e-06, 
    9.600391e-06, 9.553023e-06, 9.593228e-06, 9.542744e-06, 9.547174e-06, 
    9.560882e-06, 9.588464e-06, 9.594633e-06, 9.601147e-06, 9.597136e-06, 
    9.577566e-06, 9.57438e-06, 9.560558e-06, 9.556724e-06, 9.546213e-06, 
    9.537494e-06, 9.54545e-06, 9.553798e-06, 9.577591e-06, 9.599034e-06, 
    9.622449e-06, 9.628199e-06, 9.655491e-06, 9.633215e-06, 9.669929e-06, 
    9.638625e-06, 9.692884e-06, 9.595621e-06, 9.637789e-06, 9.56152e-06, 
    9.569733e-06, 9.584553e-06, 9.618673e-06, 9.60029e-06, 9.62181e-06, 
    9.574258e-06, 9.549578e-06, 9.543248e-06, 9.531359e-06, 9.54352e-06, 
    9.542532e-06, 9.554173e-06, 9.550434e-06, 9.578383e-06, 9.563367e-06, 
    9.606061e-06, 9.621651e-06, 9.665785e-06, 9.692856e-06, 9.720512e-06, 
    9.732709e-06, 9.736427e-06, 9.737979e-06 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.68652, 81.68573, 81.68588, 81.68524, 81.68559, 81.68518, 81.68636, 
    81.6857, 81.68612, 81.68644, 81.68404, 81.68522, 81.68274, 81.68351, 
    81.68156, 81.68287, 81.6813, 81.68159, 81.68068, 81.68094, 81.67981, 
    81.68056, 81.6792, 81.67998, 81.67986, 81.68059, 81.68496, 81.68419, 
    81.68501, 81.6849, 81.68494, 81.68559, 81.68592, 81.68658, 81.68645, 
    81.68597, 81.68485, 81.68522, 81.68426, 81.68428, 81.68322, 81.6837, 
    81.6819, 81.68241, 81.68092, 81.6813, 81.68095, 81.68105, 81.68095, 
    81.6815, 81.68126, 81.68174, 81.68361, 81.68307, 81.6847, 81.6857, 
    81.68633, 81.68679, 81.68672, 81.6866, 81.68597, 81.68536, 81.68489, 
    81.68459, 81.68428, 81.6834, 81.6829, 81.68181, 81.68199, 81.68166, 
    81.68134, 81.68081, 81.68089, 81.68066, 81.68166, 81.681, 81.6821, 
    81.6818, 81.68425, 81.68512, 81.68553, 81.68585, 81.68668, 81.68611, 
    81.68633, 81.68579, 81.68545, 81.68562, 81.68458, 81.68498, 81.68287, 
    81.68378, 81.68137, 81.68195, 81.68124, 81.68159, 81.68098, 81.68153, 
    81.68057, 81.68037, 81.6805, 81.67995, 81.68157, 81.68095, 81.68562, 
    81.6856, 81.68547, 81.68604, 81.68607, 81.68658, 81.68612, 81.68594, 
    81.68542, 81.68514, 81.68486, 81.68425, 81.68357, 81.68261, 81.68192, 
    81.68145, 81.68173, 81.68148, 81.68176, 81.68189, 81.68044, 81.68126, 
    81.68002, 81.68009, 81.68066, 81.68008, 81.68558, 81.68573, 81.68629, 
    81.68585, 81.68664, 81.6862, 81.68596, 81.68499, 81.68476, 81.68457, 
    81.68417, 81.68367, 81.6828, 81.68203, 81.68132, 81.68137, 81.68135, 
    81.6812, 81.68159, 81.68113, 81.68106, 81.68125, 81.6801, 81.68043, 
    81.68009, 81.68031, 81.68568, 81.68542, 81.68556, 81.6853, 81.68549, 
    81.68465, 81.6844, 81.68321, 81.68369, 81.68291, 81.6836, 81.68349, 
    81.68291, 81.68356, 81.68208, 81.68311, 81.68119, 81.68224, 81.68113, 
    81.68132, 81.68099, 81.68071, 81.68034, 81.67967, 81.67982, 81.67926, 
    81.68502, 81.68468, 81.68471, 81.68435, 81.68408, 81.6835, 81.68257, 
    81.68292, 81.68227, 81.68215, 81.68312, 81.68253, 81.68446, 81.68415, 
    81.68433, 81.685, 81.68285, 81.68396, 81.68191, 81.6825, 81.68075, 
    81.68163, 81.67991, 81.6792, 81.67848, 81.6777, 81.68449, 81.68472, 
    81.6843, 81.68374, 81.68319, 81.68247, 81.68239, 81.68226, 81.68191, 
    81.68161, 81.68223, 81.68154, 81.6841, 81.68275, 81.68481, 81.68421, 
    81.68377, 81.68395, 81.68295, 81.68272, 81.68179, 81.68227, 81.67938, 
    81.68066, 81.67706, 81.67808, 81.6848, 81.68449, 81.6834, 81.68391, 
    81.68242, 81.68205, 81.68175, 81.68137, 81.68132, 81.6811, 81.68147, 
    81.68111, 81.68246, 81.68186, 81.68351, 81.68311, 81.6833, 81.6835, 
    81.68287, 81.68222, 81.68219, 81.68198, 81.68143, 81.68241, 81.67924, 
    81.68123, 81.68414, 81.68356, 81.68345, 81.68369, 81.68209, 81.68267, 
    81.6811, 81.68152, 81.68083, 81.68118, 81.68123, 81.68166, 81.68195, 
    81.68265, 81.68321, 81.68365, 81.68355, 81.68306, 81.68217, 81.68133, 
    81.68151, 81.68089, 81.68253, 81.68185, 81.68211, 81.68141, 81.68293, 
    81.68169, 81.68326, 81.68311, 81.68268, 81.68181, 81.68159, 81.68139, 
    81.68151, 81.68215, 81.68225, 81.68269, 81.68282, 81.68314, 81.68343, 
    81.68317, 81.68291, 81.68214, 81.68146, 81.68071, 81.68052, 81.67968, 
    81.68038, 81.67924, 81.68024, 81.67849, 81.68159, 81.68024, 81.68266, 
    81.68239, 81.68193, 81.68084, 81.68141, 81.68074, 81.68225, 81.68305, 
    81.68324, 81.68362, 81.68324, 81.68327, 81.68289, 81.68301, 81.68211, 
    81.68259, 81.68123, 81.68074, 81.67932, 81.67846, 81.67756, 81.67717, 
    81.67705, 81.677 ;

 RH2M_R =
  81.68652, 81.68573, 81.68588, 81.68524, 81.68559, 81.68518, 81.68636, 
    81.6857, 81.68612, 81.68644, 81.68404, 81.68522, 81.68274, 81.68351, 
    81.68156, 81.68287, 81.6813, 81.68159, 81.68068, 81.68094, 81.67981, 
    81.68056, 81.6792, 81.67998, 81.67986, 81.68059, 81.68496, 81.68419, 
    81.68501, 81.6849, 81.68494, 81.68559, 81.68592, 81.68658, 81.68645, 
    81.68597, 81.68485, 81.68522, 81.68426, 81.68428, 81.68322, 81.6837, 
    81.6819, 81.68241, 81.68092, 81.6813, 81.68095, 81.68105, 81.68095, 
    81.6815, 81.68126, 81.68174, 81.68361, 81.68307, 81.6847, 81.6857, 
    81.68633, 81.68679, 81.68672, 81.6866, 81.68597, 81.68536, 81.68489, 
    81.68459, 81.68428, 81.6834, 81.6829, 81.68181, 81.68199, 81.68166, 
    81.68134, 81.68081, 81.68089, 81.68066, 81.68166, 81.681, 81.6821, 
    81.6818, 81.68425, 81.68512, 81.68553, 81.68585, 81.68668, 81.68611, 
    81.68633, 81.68579, 81.68545, 81.68562, 81.68458, 81.68498, 81.68287, 
    81.68378, 81.68137, 81.68195, 81.68124, 81.68159, 81.68098, 81.68153, 
    81.68057, 81.68037, 81.6805, 81.67995, 81.68157, 81.68095, 81.68562, 
    81.6856, 81.68547, 81.68604, 81.68607, 81.68658, 81.68612, 81.68594, 
    81.68542, 81.68514, 81.68486, 81.68425, 81.68357, 81.68261, 81.68192, 
    81.68145, 81.68173, 81.68148, 81.68176, 81.68189, 81.68044, 81.68126, 
    81.68002, 81.68009, 81.68066, 81.68008, 81.68558, 81.68573, 81.68629, 
    81.68585, 81.68664, 81.6862, 81.68596, 81.68499, 81.68476, 81.68457, 
    81.68417, 81.68367, 81.6828, 81.68203, 81.68132, 81.68137, 81.68135, 
    81.6812, 81.68159, 81.68113, 81.68106, 81.68125, 81.6801, 81.68043, 
    81.68009, 81.68031, 81.68568, 81.68542, 81.68556, 81.6853, 81.68549, 
    81.68465, 81.6844, 81.68321, 81.68369, 81.68291, 81.6836, 81.68349, 
    81.68291, 81.68356, 81.68208, 81.68311, 81.68119, 81.68224, 81.68113, 
    81.68132, 81.68099, 81.68071, 81.68034, 81.67967, 81.67982, 81.67926, 
    81.68502, 81.68468, 81.68471, 81.68435, 81.68408, 81.6835, 81.68257, 
    81.68292, 81.68227, 81.68215, 81.68312, 81.68253, 81.68446, 81.68415, 
    81.68433, 81.685, 81.68285, 81.68396, 81.68191, 81.6825, 81.68075, 
    81.68163, 81.67991, 81.6792, 81.67848, 81.6777, 81.68449, 81.68472, 
    81.6843, 81.68374, 81.68319, 81.68247, 81.68239, 81.68226, 81.68191, 
    81.68161, 81.68223, 81.68154, 81.6841, 81.68275, 81.68481, 81.68421, 
    81.68377, 81.68395, 81.68295, 81.68272, 81.68179, 81.68227, 81.67938, 
    81.68066, 81.67706, 81.67808, 81.6848, 81.68449, 81.6834, 81.68391, 
    81.68242, 81.68205, 81.68175, 81.68137, 81.68132, 81.6811, 81.68147, 
    81.68111, 81.68246, 81.68186, 81.68351, 81.68311, 81.6833, 81.6835, 
    81.68287, 81.68222, 81.68219, 81.68198, 81.68143, 81.68241, 81.67924, 
    81.68123, 81.68414, 81.68356, 81.68345, 81.68369, 81.68209, 81.68267, 
    81.6811, 81.68152, 81.68083, 81.68118, 81.68123, 81.68166, 81.68195, 
    81.68265, 81.68321, 81.68365, 81.68355, 81.68306, 81.68217, 81.68133, 
    81.68151, 81.68089, 81.68253, 81.68185, 81.68211, 81.68141, 81.68293, 
    81.68169, 81.68326, 81.68311, 81.68268, 81.68181, 81.68159, 81.68139, 
    81.68151, 81.68215, 81.68225, 81.68269, 81.68282, 81.68314, 81.68343, 
    81.68317, 81.68291, 81.68214, 81.68146, 81.68071, 81.68052, 81.67968, 
    81.68038, 81.67924, 81.68024, 81.67849, 81.68159, 81.68024, 81.68266, 
    81.68239, 81.68193, 81.68084, 81.68141, 81.68074, 81.68225, 81.68305, 
    81.68324, 81.68362, 81.68324, 81.68327, 81.68289, 81.68301, 81.68211, 
    81.68259, 81.68123, 81.68074, 81.67932, 81.67846, 81.67756, 81.67717, 
    81.67705, 81.677 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004362544, 0.0004380977, 0.0004377393, 0.000439226, 0.0004384012, 
    0.0004393746, 0.0004366279, 0.0004381705, 0.0004371857, 0.00043642, 
    0.0004421107, 0.0004392919, 0.0004450391, 0.0004432412, 0.0004477576, 
    0.0004447591, 0.0004483621, 0.000447671, 0.0004497511, 0.0004491551, 
    0.0004518154, 0.000450026, 0.0004531946, 0.000451388, 0.0004516706, 
    0.0004499667, 0.0004398596, 0.0004417601, 0.0004397469, 0.0004400179, 
    0.0004398962, 0.000438418, 0.0004376731, 0.0004361131, 0.0004363963, 
    0.000437542, 0.0004401394, 0.0004392576, 0.0004414798, 0.0004414296, 
    0.0004439035, 0.0004427881, 0.0004469464, 0.0004457645, 0.0004491799, 
    0.0004483208, 0.0004491394, 0.0004488911, 0.0004491425, 0.0004478827, 
    0.0004484224, 0.0004473139, 0.0004429976, 0.0004442663, 0.0004404821, 
    0.0004382065, 0.0004366953, 0.000435623, 0.0004357744, 0.0004360634, 
    0.0004375486, 0.0004389449, 0.0004400091, 0.0004407209, 0.0004414222, 
    0.0004435452, 0.000444669, 0.0004471853, 0.0004467312, 0.0004475004, 
    0.0004482353, 0.0004494691, 0.0004492661, 0.0004498096, 0.0004474798, 
    0.0004490281, 0.0004464721, 0.0004471711, 0.0004416132, 0.0004394958, 
    0.0004385955, 0.0004378077, 0.000435891, 0.0004372145, 0.0004366927, 
    0.000437934, 0.0004387228, 0.0004383326, 0.0004407403, 0.0004398041, 
    0.0004447355, 0.0004426114, 0.0004481497, 0.0004468243, 0.0004484672, 
    0.0004476288, 0.0004490652, 0.0004477724, 0.0004500118, 0.0004504994, 
    0.0004501661, 0.0004514463, 0.0004477004, 0.0004491388, 0.000438322, 
    0.0004383856, 0.0004386819, 0.0004373788, 0.0004372991, 0.000436105, 
    0.0004371674, 0.0004376198, 0.0004387684, 0.0004394476, 0.0004400934, 
    0.0004415134, 0.0004430992, 0.0004453168, 0.0004469101, 0.0004479781, 
    0.0004473232, 0.0004479013, 0.0004472549, 0.0004469519, 0.0004503166, 
    0.0004484272, 0.000451262, 0.0004511052, 0.0004498221, 0.0004511227, 
    0.0004384301, 0.000438064, 0.0004367927, 0.0004377875, 0.0004359749, 
    0.0004369894, 0.0004375727, 0.0004398235, 0.0004403181, 0.0004407767, 
    0.0004416824, 0.0004428447, 0.0004448839, 0.0004466581, 0.0004482779, 
    0.0004481591, 0.0004482009, 0.0004485626, 0.0004476663, 0.0004487096, 
    0.0004488847, 0.0004484268, 0.000451084, 0.0004503248, 0.0004511016, 
    0.0004506072, 0.0004381829, 0.0004387989, 0.0004384659, 0.0004390919, 
    0.0004386507, 0.0004406118, 0.0004411997, 0.000443951, 0.0004428218, 
    0.0004446189, 0.0004430043, 0.0004432904, 0.0004446772, 0.0004430914, 
    0.00044656, 0.0004442082, 0.0004485766, 0.0004462279, 0.0004487237, 
    0.0004482704, 0.0004490207, 0.0004496927, 0.000450538, 0.0004520979, 
    0.0004517366, 0.0004530412, 0.0004397173, 0.0004405163, 0.0004404459, 
    0.0004412821, 0.0004419005, 0.0004432411, 0.0004453911, 0.0004445825, 
    0.0004460668, 0.0004463647, 0.0004441096, 0.0004454941, 0.0004410505, 
    0.0004417683, 0.0004413409, 0.0004397795, 0.0004447683, 0.0004422078, 
    0.0004469358, 0.0004455486, 0.0004495967, 0.0004475834, 0.0004515377, 
    0.0004532281, 0.0004548192, 0.0004566784, 0.0004409524, 0.0004404093, 
    0.0004413815, 0.0004427265, 0.0004439746, 0.0004456339, 0.0004458036, 
    0.0004461144, 0.0004469196, 0.0004475966, 0.0004462125, 0.0004477662, 
    0.0004419346, 0.0004449905, 0.0004402033, 0.0004416447, 0.0004426465, 
    0.0004422071, 0.0004444894, 0.0004450272, 0.0004472131, 0.0004460831, 
    0.0004528107, 0.0004498342, 0.0004580941, 0.0004557857, 0.0004402195, 
    0.0004409503, 0.0004434937, 0.0004422835, 0.0004457445, 0.0004465965, 
    0.000447289, 0.0004481743, 0.0004482698, 0.0004487944, 0.0004479347, 
    0.0004487603, 0.0004456368, 0.0004470326, 0.0004432024, 0.0004441345, 
    0.0004437057, 0.0004432352, 0.000444687, 0.0004462336, 0.0004462667, 
    0.0004467626, 0.0004481599, 0.0004457576, 0.0004531945, 0.0004486013, 
    0.0004417472, 0.0004431547, 0.0004433558, 0.0004428105, 0.0004465109, 
    0.0004451701, 0.0004487816, 0.0004478054, 0.0004494047, 0.00044861, 
    0.0004484929, 0.0004474722, 0.0004468366, 0.0004452311, 0.0004439247, 
    0.0004428889, 0.0004431297, 0.0004442675, 0.0004463281, 0.0004482777, 
    0.0004478506, 0.0004492824, 0.0004454924, 0.0004470816, 0.0004464673, 
    0.0004480689, 0.0004445608, 0.0004475488, 0.0004437969, 0.0004441258, 
    0.0004451433, 0.0004471901, 0.000447643, 0.0004481265, 0.0004478281, 
    0.0004463809, 0.0004461437, 0.0004451182, 0.000444835, 0.0004440537, 
    0.0004434067, 0.0004439977, 0.0004446182, 0.0004463811, 0.0004479696, 
    0.0004497016, 0.0004501255, 0.0004521489, 0.0004505015, 0.0004532198, 
    0.0004509085, 0.0004549095, 0.0004477219, 0.0004508418, 0.0004451896, 
    0.0004457985, 0.0004468997, 0.0004494257, 0.000448062, 0.0004496569, 
    0.0004461344, 0.0004443068, 0.000443834, 0.0004429518, 0.000443854, 
    0.0004437806, 0.000444644, 0.0004443665, 0.0004464394, 0.0004453259, 
    0.0004484892, 0.0004496436, 0.0004529038, 0.0004549024, 0.000456937, 
    0.0004578352, 0.0004581086, 0.0004582228 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.475499e-14, 3.485026e-14, 3.483175e-14, 3.490853e-14, 3.486596e-14, 
    3.491621e-14, 3.477432e-14, 3.485402e-14, 3.480316e-14, 3.476359e-14, 
    3.505735e-14, 3.491196e-14, 3.520834e-14, 3.511572e-14, 3.534828e-14, 
    3.519391e-14, 3.537938e-14, 3.534386e-14, 3.545083e-14, 3.54202e-14, 
    3.555682e-14, 3.546496e-14, 3.562763e-14, 3.553491e-14, 3.554941e-14, 
    3.546193e-14, 3.494126e-14, 3.503925e-14, 3.493545e-14, 3.494943e-14, 
    3.494316e-14, 3.486682e-14, 3.482831e-14, 3.474773e-14, 3.476237e-14, 
    3.482157e-14, 3.495571e-14, 3.491022e-14, 3.502492e-14, 3.502233e-14, 
    3.514988e-14, 3.509239e-14, 3.530658e-14, 3.524575e-14, 3.542147e-14, 
    3.53773e-14, 3.541939e-14, 3.540664e-14, 3.541956e-14, 3.535477e-14, 
    3.538253e-14, 3.532552e-14, 3.510315e-14, 3.516853e-14, 3.49734e-14, 
    3.485586e-14, 3.477781e-14, 3.472238e-14, 3.473022e-14, 3.474515e-14, 
    3.482191e-14, 3.489407e-14, 3.494902e-14, 3.498576e-14, 3.502196e-14, 
    3.513136e-14, 3.51893e-14, 3.531886e-14, 3.529552e-14, 3.533508e-14, 
    3.537291e-14, 3.543635e-14, 3.542591e-14, 3.545384e-14, 3.533406e-14, 
    3.541368e-14, 3.528222e-14, 3.531818e-14, 3.503168e-14, 3.49225e-14, 
    3.487596e-14, 3.48353e-14, 3.473624e-14, 3.480465e-14, 3.477769e-14, 
    3.484186e-14, 3.48826e-14, 3.486246e-14, 3.498677e-14, 3.493845e-14, 
    3.519273e-14, 3.508327e-14, 3.53685e-14, 3.530031e-14, 3.538484e-14, 
    3.534172e-14, 3.541558e-14, 3.534911e-14, 3.546425e-14, 3.548929e-14, 
    3.547217e-14, 3.553794e-14, 3.534542e-14, 3.541938e-14, 3.486189e-14, 
    3.486517e-14, 3.488048e-14, 3.481315e-14, 3.480903e-14, 3.474732e-14, 
    3.480224e-14, 3.482561e-14, 3.488497e-14, 3.492004e-14, 3.495338e-14, 
    3.502666e-14, 3.510842e-14, 3.522269e-14, 3.530473e-14, 3.535969e-14, 
    3.5326e-14, 3.535574e-14, 3.532249e-14, 3.530691e-14, 3.54799e-14, 
    3.538279e-14, 3.552849e-14, 3.552043e-14, 3.545451e-14, 3.552134e-14, 
    3.486748e-14, 3.484857e-14, 3.478287e-14, 3.483429e-14, 3.47406e-14, 
    3.479304e-14, 3.482317e-14, 3.493943e-14, 3.496499e-14, 3.498865e-14, 
    3.503539e-14, 3.509533e-14, 3.52004e-14, 3.529176e-14, 3.537511e-14, 
    3.536901e-14, 3.537116e-14, 3.538976e-14, 3.534366e-14, 3.539733e-14, 
    3.540632e-14, 3.538279e-14, 3.551935e-14, 3.548036e-14, 3.552026e-14, 
    3.549487e-14, 3.485472e-14, 3.488654e-14, 3.486934e-14, 3.490167e-14, 
    3.487889e-14, 3.498011e-14, 3.501045e-14, 3.515231e-14, 3.509414e-14, 
    3.518674e-14, 3.510356e-14, 3.51183e-14, 3.518971e-14, 3.510807e-14, 
    3.52867e-14, 3.516558e-14, 3.539048e-14, 3.526959e-14, 3.539805e-14, 
    3.537476e-14, 3.541334e-14, 3.544787e-14, 3.549132e-14, 3.55714e-14, 
    3.555287e-14, 3.561983e-14, 3.493396e-14, 3.497519e-14, 3.497158e-14, 
    3.501474e-14, 3.504663e-14, 3.511576e-14, 3.522653e-14, 3.518489e-14, 
    3.526134e-14, 3.527667e-14, 3.516054e-14, 3.523184e-14, 3.50028e-14, 
    3.503981e-14, 3.501779e-14, 3.493721e-14, 3.519446e-14, 3.506249e-14, 
    3.530608e-14, 3.523469e-14, 3.544294e-14, 3.53394e-14, 3.554266e-14, 
    3.562937e-14, 3.571103e-14, 3.580624e-14, 3.499771e-14, 3.49697e-14, 
    3.501987e-14, 3.508921e-14, 3.515356e-14, 3.523904e-14, 3.524779e-14, 
    3.526379e-14, 3.530524e-14, 3.534008e-14, 3.526883e-14, 3.534881e-14, 
    3.504835e-14, 3.520592e-14, 3.495909e-14, 3.503344e-14, 3.508513e-14, 
    3.506248e-14, 3.518014e-14, 3.520785e-14, 3.532036e-14, 3.526223e-14, 
    3.560796e-14, 3.545513e-14, 3.587875e-14, 3.576053e-14, 3.495991e-14, 
    3.499763e-14, 3.512877e-14, 3.506639e-14, 3.524475e-14, 3.528861e-14, 
    3.532426e-14, 3.536978e-14, 3.537471e-14, 3.540168e-14, 3.535748e-14, 
    3.539994e-14, 3.523922e-14, 3.531108e-14, 3.511382e-14, 3.516185e-14, 
    3.513976e-14, 3.511551e-14, 3.519033e-14, 3.526994e-14, 3.527168e-14, 
    3.529719e-14, 3.536898e-14, 3.524548e-14, 3.56276e-14, 3.539171e-14, 
    3.503874e-14, 3.511128e-14, 3.512169e-14, 3.509358e-14, 3.528421e-14, 
    3.521517e-14, 3.540103e-14, 3.535083e-14, 3.543307e-14, 3.539221e-14, 
    3.53862e-14, 3.53337e-14, 3.530099e-14, 3.521833e-14, 3.515103e-14, 
    3.509766e-14, 3.511008e-14, 3.51687e-14, 3.527482e-14, 3.537514e-14, 
    3.535317e-14, 3.542682e-14, 3.523183e-14, 3.531362e-14, 3.5282e-14, 
    3.536443e-14, 3.518378e-14, 3.533752e-14, 3.514444e-14, 3.516139e-14, 
    3.52138e-14, 3.531914e-14, 3.534248e-14, 3.536734e-14, 3.535201e-14, 
    3.527752e-14, 3.526533e-14, 3.521254e-14, 3.519794e-14, 3.51577e-14, 
    3.512436e-14, 3.515481e-14, 3.518678e-14, 3.527756e-14, 3.53593e-14, 
    3.544835e-14, 3.547015e-14, 3.5574e-14, 3.548942e-14, 3.562891e-14, 
    3.551026e-14, 3.57156e-14, 3.534647e-14, 3.550684e-14, 3.521619e-14, 
    3.524755e-14, 3.53042e-14, 3.543412e-14, 3.536404e-14, 3.544601e-14, 
    3.526485e-14, 3.517071e-14, 3.514638e-14, 3.51009e-14, 3.514742e-14, 
    3.514363e-14, 3.518813e-14, 3.517383e-14, 3.528058e-14, 3.522325e-14, 
    3.538603e-14, 3.544537e-14, 3.56128e-14, 3.571529e-14, 3.581956e-14, 
    3.586554e-14, 3.587954e-14, 3.588538e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.155628e-14, 1.158799e-14, 1.158183e-14, 1.160739e-14, 1.159322e-14, 
    1.160994e-14, 1.156272e-14, 1.158924e-14, 1.157231e-14, 1.155914e-14, 
    1.165692e-14, 1.160853e-14, 1.170718e-14, 1.167635e-14, 1.175376e-14, 
    1.170237e-14, 1.176411e-14, 1.175229e-14, 1.178789e-14, 1.177769e-14, 
    1.182317e-14, 1.179259e-14, 1.184674e-14, 1.181588e-14, 1.18207e-14, 
    1.179158e-14, 1.161828e-14, 1.165089e-14, 1.161635e-14, 1.1621e-14, 
    1.161891e-14, 1.15935e-14, 1.158069e-14, 1.155386e-14, 1.155874e-14, 
    1.157844e-14, 1.162309e-14, 1.160795e-14, 1.164612e-14, 1.164526e-14, 
    1.168772e-14, 1.166858e-14, 1.173988e-14, 1.171963e-14, 1.177812e-14, 
    1.176342e-14, 1.177743e-14, 1.177318e-14, 1.177748e-14, 1.175592e-14, 
    1.176516e-14, 1.174618e-14, 1.167216e-14, 1.169393e-14, 1.162898e-14, 
    1.158985e-14, 1.156388e-14, 1.154543e-14, 1.154804e-14, 1.155301e-14, 
    1.157856e-14, 1.160257e-14, 1.162086e-14, 1.163309e-14, 1.164514e-14, 
    1.168155e-14, 1.170084e-14, 1.174396e-14, 1.17362e-14, 1.174936e-14, 
    1.176195e-14, 1.178307e-14, 1.17796e-14, 1.178889e-14, 1.174902e-14, 
    1.177552e-14, 1.173177e-14, 1.174374e-14, 1.164838e-14, 1.161203e-14, 
    1.159655e-14, 1.158301e-14, 1.155004e-14, 1.157281e-14, 1.156384e-14, 
    1.158519e-14, 1.159876e-14, 1.159205e-14, 1.163343e-14, 1.161734e-14, 
    1.170198e-14, 1.166555e-14, 1.176049e-14, 1.173779e-14, 1.176593e-14, 
    1.175157e-14, 1.177616e-14, 1.175403e-14, 1.179236e-14, 1.180069e-14, 
    1.1795e-14, 1.181689e-14, 1.17528e-14, 1.177742e-14, 1.159186e-14, 
    1.159295e-14, 1.159805e-14, 1.157564e-14, 1.157427e-14, 1.155373e-14, 
    1.157201e-14, 1.157979e-14, 1.159954e-14, 1.161122e-14, 1.162232e-14, 
    1.16467e-14, 1.167392e-14, 1.171195e-14, 1.173926e-14, 1.175755e-14, 
    1.174634e-14, 1.175624e-14, 1.174517e-14, 1.173999e-14, 1.179757e-14, 
    1.176524e-14, 1.181374e-14, 1.181106e-14, 1.178911e-14, 1.181136e-14, 
    1.159372e-14, 1.158743e-14, 1.156556e-14, 1.158267e-14, 1.155149e-14, 
    1.156894e-14, 1.157897e-14, 1.161767e-14, 1.162618e-14, 1.163405e-14, 
    1.164961e-14, 1.166956e-14, 1.170453e-14, 1.173494e-14, 1.176269e-14, 
    1.176066e-14, 1.176137e-14, 1.176756e-14, 1.175222e-14, 1.177008e-14, 
    1.177308e-14, 1.176524e-14, 1.18107e-14, 1.179772e-14, 1.1811e-14, 
    1.180255e-14, 1.158948e-14, 1.160007e-14, 1.159434e-14, 1.16051e-14, 
    1.159752e-14, 1.163121e-14, 1.164131e-14, 1.168853e-14, 1.166917e-14, 
    1.169999e-14, 1.16723e-14, 1.167721e-14, 1.170098e-14, 1.16738e-14, 
    1.173326e-14, 1.169294e-14, 1.17678e-14, 1.172756e-14, 1.177032e-14, 
    1.176257e-14, 1.177541e-14, 1.17869e-14, 1.180137e-14, 1.182802e-14, 
    1.182185e-14, 1.184414e-14, 1.161585e-14, 1.162957e-14, 1.162837e-14, 
    1.164274e-14, 1.165335e-14, 1.167636e-14, 1.171323e-14, 1.169937e-14, 
    1.172482e-14, 1.172992e-14, 1.169127e-14, 1.1715e-14, 1.163876e-14, 
    1.165108e-14, 1.164375e-14, 1.161693e-14, 1.170256e-14, 1.165863e-14, 
    1.173971e-14, 1.171595e-14, 1.178526e-14, 1.17508e-14, 1.181846e-14, 
    1.184732e-14, 1.18745e-14, 1.190619e-14, 1.163707e-14, 1.162775e-14, 
    1.164444e-14, 1.166752e-14, 1.168895e-14, 1.171739e-14, 1.172031e-14, 
    1.172563e-14, 1.173943e-14, 1.175103e-14, 1.172731e-14, 1.175393e-14, 
    1.165392e-14, 1.170637e-14, 1.162422e-14, 1.164896e-14, 1.166617e-14, 
    1.165863e-14, 1.169779e-14, 1.170701e-14, 1.174446e-14, 1.172511e-14, 
    1.184019e-14, 1.178932e-14, 1.193033e-14, 1.189098e-14, 1.162449e-14, 
    1.163704e-14, 1.168069e-14, 1.165993e-14, 1.17193e-14, 1.173389e-14, 
    1.174576e-14, 1.176091e-14, 1.176255e-14, 1.177153e-14, 1.175682e-14, 
    1.177095e-14, 1.171745e-14, 1.174137e-14, 1.167571e-14, 1.16917e-14, 
    1.168435e-14, 1.167628e-14, 1.170118e-14, 1.172768e-14, 1.172826e-14, 
    1.173675e-14, 1.176065e-14, 1.171954e-14, 1.184673e-14, 1.176821e-14, 
    1.165073e-14, 1.167487e-14, 1.167833e-14, 1.166898e-14, 1.173243e-14, 
    1.170945e-14, 1.177131e-14, 1.175461e-14, 1.178198e-14, 1.176838e-14, 
    1.176638e-14, 1.17489e-14, 1.173802e-14, 1.17105e-14, 1.16881e-14, 
    1.167034e-14, 1.167447e-14, 1.169398e-14, 1.17293e-14, 1.17627e-14, 
    1.175538e-14, 1.17799e-14, 1.1715e-14, 1.174222e-14, 1.17317e-14, 
    1.175913e-14, 1.1699e-14, 1.175017e-14, 1.168591e-14, 1.169155e-14, 
    1.170899e-14, 1.174406e-14, 1.175183e-14, 1.17601e-14, 1.1755e-14, 
    1.17302e-14, 1.172614e-14, 1.170857e-14, 1.170371e-14, 1.169032e-14, 
    1.167922e-14, 1.168936e-14, 1.17e-14, 1.173022e-14, 1.175742e-14, 
    1.178707e-14, 1.179432e-14, 1.182889e-14, 1.180074e-14, 1.184716e-14, 
    1.180767e-14, 1.187602e-14, 1.175316e-14, 1.180653e-14, 1.170979e-14, 
    1.172023e-14, 1.173909e-14, 1.178233e-14, 1.1759e-14, 1.178628e-14, 
    1.172599e-14, 1.169465e-14, 1.168655e-14, 1.167142e-14, 1.16869e-14, 
    1.168564e-14, 1.170045e-14, 1.169569e-14, 1.173122e-14, 1.171214e-14, 
    1.176632e-14, 1.178607e-14, 1.18418e-14, 1.187592e-14, 1.191063e-14, 
    1.192593e-14, 1.193059e-14, 1.193254e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.145939e-11, -8.181889e-11, -8.1749e-11, -8.203896e-11, -8.187812e-11, 
    -8.206798e-11, -8.153229e-11, -8.183315e-11, -8.164109e-11, 
    -8.149177e-11, -8.260167e-11, -8.20519e-11, -8.317288e-11, -8.28222e-11, 
    -8.370318e-11, -8.31183e-11, -8.382113e-11, -8.368634e-11, -8.40921e-11, 
    -8.397585e-11, -8.449484e-11, -8.414575e-11, -8.476393e-11, 
    -8.441148e-11, -8.446661e-11, -8.413423e-11, -8.216255e-11, 
    -8.253322e-11, -8.214059e-11, -8.219344e-11, -8.216973e-11, 
    -8.188144e-11, -8.173615e-11, -8.143194e-11, -8.148716e-11, 
    -8.171061e-11, -8.221721e-11, -8.204525e-11, -8.247868e-11, 
    -8.246889e-11, -8.295144e-11, -8.273387e-11, -8.3545e-11, -8.331446e-11, 
    -8.39807e-11, -8.381314e-11, -8.397283e-11, -8.392442e-11, -8.397346e-11, 
    -8.372772e-11, -8.3833e-11, -8.361677e-11, -8.277461e-11, -8.30221e-11, 
    -8.228399e-11, -8.184019e-11, -8.154548e-11, -8.133634e-11, 
    -8.136591e-11, -8.142226e-11, -8.171192e-11, -8.198427e-11, 
    -8.219184e-11, -8.233068e-11, -8.246748e-11, -8.288156e-11, 
    -8.310078e-11, -8.359161e-11, -8.350304e-11, -8.36531e-11, -8.379648e-11, 
    -8.403717e-11, -8.399756e-11, -8.410361e-11, -8.364915e-11, 
    -8.395117e-11, -8.345259e-11, -8.358896e-11, -8.250461e-11, 
    -8.209165e-11, -8.191606e-11, -8.176244e-11, -8.138864e-11, 
    -8.164677e-11, -8.154501e-11, -8.178712e-11, -8.194095e-11, 
    -8.186488e-11, -8.233447e-11, -8.21519e-11, -8.311377e-11, -8.269944e-11, 
    -8.377975e-11, -8.352122e-11, -8.384172e-11, -8.367818e-11, -8.39584e-11, 
    -8.37062e-11, -8.414307e-11, -8.42382e-11, -8.41732e-11, -8.442293e-11, 
    -8.369223e-11, -8.397282e-11, -8.186274e-11, -8.187515e-11, 
    -8.193296e-11, -8.167882e-11, -8.166328e-11, -8.143042e-11, 
    -8.163763e-11, -8.172586e-11, -8.194988e-11, -8.208238e-11, 
    -8.220834e-11, -8.24853e-11, -8.279461e-11, -8.322718e-11, -8.353798e-11, 
    -8.374632e-11, -8.361858e-11, -8.373136e-11, -8.360528e-11, 
    -8.354619e-11, -8.420255e-11, -8.383398e-11, -8.438701e-11, 
    -8.435641e-11, -8.410612e-11, -8.435986e-11, -8.188386e-11, 
    -8.181245e-11, -8.156453e-11, -8.175855e-11, -8.140506e-11, 
    -8.160292e-11, -8.171668e-11, -8.21557e-11, -8.225218e-11, -8.234161e-11, 
    -8.251828e-11, -8.274501e-11, -8.314274e-11, -8.348884e-11, 
    -8.380482e-11, -8.378167e-11, -8.378982e-11, -8.38604e-11, -8.368556e-11, 
    -8.38891e-11, -8.392326e-11, -8.383395e-11, -8.435231e-11, -8.420422e-11, 
    -8.435576e-11, -8.425934e-11, -8.183567e-11, -8.195582e-11, 
    -8.189089e-11, -8.201298e-11, -8.192697e-11, -8.230944e-11, 
    -8.242412e-11, -8.296077e-11, -8.274054e-11, -8.309106e-11, 
    -8.277615e-11, -8.283194e-11, -8.310246e-11, -8.279317e-11, 
    -8.346975e-11, -8.301101e-11, -8.386314e-11, -8.3405e-11, -8.389185e-11, 
    -8.380345e-11, -8.394982e-11, -8.408091e-11, -8.424584e-11, 
    -8.455014e-11, -8.447968e-11, -8.473419e-11, -8.213495e-11, -8.22908e-11, 
    -8.227709e-11, -8.244019e-11, -8.256083e-11, -8.28223e-11, -8.324168e-11, 
    -8.308398e-11, -8.337351e-11, -8.343163e-11, -8.299177e-11, 
    -8.326182e-11, -8.239511e-11, -8.253512e-11, -8.245177e-11, 
    -8.214724e-11, -8.31203e-11, -8.26209e-11, -8.354312e-11, -8.327256e-11, 
    -8.406222e-11, -8.366948e-11, -8.444088e-11, -8.477065e-11, 
    -8.508109e-11, -8.544382e-11, -8.237587e-11, -8.226998e-11, 
    -8.245959e-11, -8.272194e-11, -8.29654e-11, -8.328906e-11, -8.332218e-11, 
    -8.338281e-11, -8.353988e-11, -8.367194e-11, -8.340197e-11, 
    -8.370506e-11, -8.256757e-11, -8.316365e-11, -8.222992e-11, 
    -8.251106e-11, -8.270648e-11, -8.262076e-11, -8.306595e-11, 
    -8.317088e-11, -8.359727e-11, -8.337685e-11, -8.468925e-11, 
    -8.410858e-11, -8.572006e-11, -8.526967e-11, -8.223297e-11, 
    -8.237551e-11, -8.287161e-11, -8.263557e-11, -8.331067e-11, 
    -8.347685e-11, -8.361196e-11, -8.378465e-11, -8.38033e-11, -8.390563e-11, 
    -8.373795e-11, -8.389901e-11, -8.328974e-11, -8.3562e-11, -8.281491e-11, 
    -8.299673e-11, -8.291309e-11, -8.282134e-11, -8.310453e-11, 
    -8.340622e-11, -8.341269e-11, -8.350942e-11, -8.3782e-11, -8.33134e-11, 
    -8.476416e-11, -8.386814e-11, -8.253095e-11, -8.280549e-11, 
    -8.284473e-11, -8.273837e-11, -8.346019e-11, -8.319864e-11, 
    -8.390313e-11, -8.371273e-11, -8.402471e-11, -8.386968e-11, 
    -8.384687e-11, -8.364776e-11, -8.35238e-11, -8.321063e-11, -8.295583e-11, 
    -8.27538e-11, -8.280078e-11, -8.302271e-11, -8.342468e-11, -8.380498e-11, 
    -8.372168e-11, -8.4001e-11, -8.326172e-11, -8.357169e-11, -8.345188e-11, 
    -8.37643e-11, -8.307978e-11, -8.366262e-11, -8.29308e-11, -8.299497e-11, 
    -8.319345e-11, -8.35927e-11, -8.368107e-11, -8.377538e-11, -8.371719e-11, 
    -8.343488e-11, -8.338864e-11, -8.318863e-11, -8.313339e-11, -8.2981e-11, 
    -8.285482e-11, -8.29701e-11, -8.309116e-11, -8.343501e-11, -8.374489e-11, 
    -8.408277e-11, -8.416547e-11, -8.456021e-11, -8.423885e-11, 
    -8.476915e-11, -8.431825e-11, -8.509882e-11, -8.369643e-11, 
    -8.430502e-11, -8.320249e-11, -8.332126e-11, -8.353608e-11, 
    -8.402884e-11, -8.376283e-11, -8.407394e-11, -8.338683e-11, 
    -8.303035e-11, -8.293815e-11, -8.276608e-11, -8.294208e-11, 
    -8.292777e-11, -8.309618e-11, -8.304207e-11, -8.344643e-11, 
    -8.322922e-11, -8.384629e-11, -8.407149e-11, -8.470751e-11, 
    -8.509743e-11, -8.54944e-11, -8.566964e-11, -8.572299e-11, -8.574529e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.963328e-12, -1.97199e-12, -1.970306e-12, -1.977293e-12, -1.973418e-12, 
    -1.977992e-12, -1.965084e-12, -1.972334e-12, -1.967706e-12, 
    -1.964108e-12, -1.990853e-12, -1.977605e-12, -2.004617e-12, 
    -1.996167e-12, -2.017395e-12, -2.003302e-12, -2.020237e-12, 
    -2.016989e-12, -2.026767e-12, -2.023966e-12, -2.036471e-12, -2.02806e-12, 
    -2.042955e-12, -2.034463e-12, -2.035791e-12, -2.027782e-12, 
    -1.980271e-12, -1.989203e-12, -1.979742e-12, -1.981016e-12, 
    -1.980444e-12, -1.973497e-12, -1.969996e-12, -1.962666e-12, 
    -1.963997e-12, -1.969381e-12, -1.981588e-12, -1.977445e-12, 
    -1.987889e-12, -1.987653e-12, -1.999281e-12, -1.994038e-12, 
    -2.013584e-12, -2.008028e-12, -2.024083e-12, -2.020045e-12, 
    -2.023893e-12, -2.022726e-12, -2.023908e-12, -2.017986e-12, 
    -2.020524e-12, -2.015313e-12, -1.99502e-12, -2.000983e-12, -1.983197e-12, 
    -1.972503e-12, -1.965402e-12, -1.960362e-12, -1.961075e-12, 
    -1.962433e-12, -1.969412e-12, -1.975975e-12, -1.980977e-12, 
    -1.984322e-12, -1.987619e-12, -1.997597e-12, -2.002879e-12, 
    -2.014707e-12, -2.012573e-12, -2.016188e-12, -2.019643e-12, 
    -2.025443e-12, -2.024489e-12, -2.027044e-12, -2.016093e-12, 
    -2.023371e-12, -2.011357e-12, -2.014643e-12, -1.988514e-12, 
    -1.978563e-12, -1.974332e-12, -1.97063e-12, -1.961622e-12, -1.967843e-12, 
    -1.965391e-12, -1.971225e-12, -1.974932e-12, -1.973098e-12, 
    -1.984414e-12, -1.980014e-12, -2.003192e-12, -1.993209e-12, -2.01924e-12, 
    -2.013011e-12, -2.020733e-12, -2.016793e-12, -2.023545e-12, 
    -2.017468e-12, -2.027995e-12, -2.030287e-12, -2.028721e-12, 
    -2.034739e-12, -2.017131e-12, -2.023893e-12, -1.973047e-12, 
    -1.973346e-12, -1.974739e-12, -1.968615e-12, -1.96824e-12, -1.962629e-12, 
    -1.967622e-12, -1.969748e-12, -1.975147e-12, -1.978339e-12, 
    -1.981374e-12, -1.988048e-12, -1.995502e-12, -2.005925e-12, 
    -2.013414e-12, -2.018435e-12, -2.015356e-12, -2.018074e-12, 
    -2.015036e-12, -2.013612e-12, -2.029428e-12, -2.020547e-12, 
    -2.033873e-12, -2.033136e-12, -2.027105e-12, -2.033219e-12, 
    -1.973556e-12, -1.971835e-12, -1.965861e-12, -1.970536e-12, 
    -1.962018e-12, -1.966786e-12, -1.969527e-12, -1.980106e-12, 
    -1.982431e-12, -1.984586e-12, -1.988843e-12, -1.994306e-12, 
    -2.003891e-12, -2.01223e-12, -2.019844e-12, -2.019286e-12, -2.019483e-12, 
    -2.021184e-12, -2.016971e-12, -2.021875e-12, -2.022698e-12, 
    -2.020546e-12, -2.033037e-12, -2.029468e-12, -2.03312e-12, -2.030797e-12, 
    -1.972394e-12, -1.97529e-12, -1.973725e-12, -1.976667e-12, -1.974594e-12, 
    -1.983811e-12, -1.986574e-12, -1.999506e-12, -1.994199e-12, 
    -2.002645e-12, -1.995057e-12, -1.996401e-12, -2.00292e-12, -1.995467e-12, 
    -2.01177e-12, -2.000716e-12, -2.02125e-12, -2.01021e-12, -2.021941e-12, 
    -2.019811e-12, -2.023338e-12, -2.026497e-12, -2.030471e-12, 
    -2.037804e-12, -2.036106e-12, -2.042239e-12, -1.979606e-12, 
    -1.983362e-12, -1.983031e-12, -1.986962e-12, -1.989868e-12, 
    -1.996169e-12, -2.006274e-12, -2.002474e-12, -2.009451e-12, 
    -2.010852e-12, -2.000252e-12, -2.00676e-12, -1.985875e-12, -1.989249e-12, 
    -1.98724e-12, -1.979902e-12, -2.00335e-12, -1.991316e-12, -2.013538e-12, 
    -2.007019e-12, -2.026047e-12, -2.016583e-12, -2.035171e-12, 
    -2.043117e-12, -2.050598e-12, -2.059338e-12, -1.985411e-12, -1.98286e-12, 
    -1.987429e-12, -1.993751e-12, -1.999617e-12, -2.007416e-12, 
    -2.008214e-12, -2.009675e-12, -2.01346e-12, -2.016642e-12, -2.010137e-12, 
    -2.01744e-12, -1.990031e-12, -2.004394e-12, -1.981895e-12, -1.988669e-12, 
    -1.993378e-12, -1.991313e-12, -2.00204e-12, -2.004569e-12, -2.014843e-12, 
    -2.009532e-12, -2.041156e-12, -2.027164e-12, -2.065995e-12, 
    -2.055142e-12, -1.981968e-12, -1.985403e-12, -1.997357e-12, 
    -1.991669e-12, -2.007937e-12, -2.011941e-12, -2.015197e-12, 
    -2.019358e-12, -2.019808e-12, -2.022273e-12, -2.018233e-12, 
    -2.022114e-12, -2.007433e-12, -2.013993e-12, -1.995991e-12, 
    -2.000372e-12, -1.998357e-12, -1.996146e-12, -2.00297e-12, -2.010239e-12, 
    -2.010395e-12, -2.012726e-12, -2.019294e-12, -2.008003e-12, 
    -2.042961e-12, -2.02137e-12, -1.989148e-12, -1.995764e-12, -1.996709e-12, 
    -1.994147e-12, -2.01154e-12, -2.005238e-12, -2.022213e-12, -2.017625e-12, 
    -2.025143e-12, -2.021407e-12, -2.020858e-12, -2.01606e-12, -2.013073e-12, 
    -2.005526e-12, -1.999387e-12, -1.994518e-12, -1.99565e-12, -2.000998e-12, 
    -2.010684e-12, -2.019848e-12, -2.017841e-12, -2.024572e-12, 
    -2.006757e-12, -2.014227e-12, -2.01134e-12, -2.018868e-12, -2.002373e-12, 
    -2.016418e-12, -1.998784e-12, -2.00033e-12, -2.005112e-12, -2.014733e-12, 
    -2.016862e-12, -2.019135e-12, -2.017733e-12, -2.01093e-12, -2.009816e-12, 
    -2.004996e-12, -2.003665e-12, -1.999993e-12, -1.996953e-12, -1.99973e-12, 
    -2.002648e-12, -2.010933e-12, -2.0184e-12, -2.026542e-12, -2.028535e-12, 
    -2.038047e-12, -2.030303e-12, -2.043081e-12, -2.032216e-12, 
    -2.051025e-12, -2.017233e-12, -2.031897e-12, -2.00533e-12, -2.008192e-12, 
    -2.013369e-12, -2.025242e-12, -2.018833e-12, -2.026329e-12, 
    -2.009772e-12, -2.001182e-12, -1.99896e-12, -1.994814e-12, -1.999055e-12, 
    -1.99871e-12, -2.002769e-12, -2.001465e-12, -2.011208e-12, -2.005974e-12, 
    -2.020844e-12, -2.02627e-12, -2.041596e-12, -2.050992e-12, -2.060557e-12, 
    -2.06478e-12, -2.066065e-12, -2.066603e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.754104e-15, 3.764405e-15, 3.762403e-15, 3.770706e-15, 3.766102e-15, 
    3.771536e-15, 3.756195e-15, 3.764812e-15, 3.759312e-15, 3.755034e-15, 
    3.786797e-15, 3.771076e-15, 3.803123e-15, 3.793109e-15, 3.818254e-15, 
    3.801563e-15, 3.821618e-15, 3.817777e-15, 3.829343e-15, 3.826031e-15, 
    3.840804e-15, 3.830871e-15, 3.848461e-15, 3.838435e-15, 3.840002e-15, 
    3.830543e-15, 3.774245e-15, 3.78484e-15, 3.773616e-15, 3.775128e-15, 
    3.77445e-15, 3.766196e-15, 3.762032e-15, 3.753319e-15, 3.754902e-15, 
    3.761303e-15, 3.775807e-15, 3.770888e-15, 3.78329e-15, 3.783011e-15, 
    3.796801e-15, 3.790585e-15, 3.813746e-15, 3.807168e-15, 3.826169e-15, 
    3.821393e-15, 3.825944e-15, 3.824565e-15, 3.825962e-15, 3.818957e-15, 
    3.821958e-15, 3.815794e-15, 3.791749e-15, 3.798819e-15, 3.777719e-15, 
    3.765011e-15, 3.756572e-15, 3.750578e-15, 3.751425e-15, 3.75304e-15, 
    3.76134e-15, 3.769142e-15, 3.775084e-15, 3.779057e-15, 3.78297e-15, 
    3.794799e-15, 3.801064e-15, 3.815074e-15, 3.81255e-15, 3.816828e-15, 
    3.820918e-15, 3.827777e-15, 3.826649e-15, 3.829669e-15, 3.816717e-15, 
    3.825326e-15, 3.811111e-15, 3.815e-15, 3.784021e-15, 3.772216e-15, 
    3.767184e-15, 3.762788e-15, 3.752077e-15, 3.759474e-15, 3.756558e-15, 
    3.763497e-15, 3.767902e-15, 3.765724e-15, 3.779165e-15, 3.77394e-15, 
    3.801435e-15, 3.7896e-15, 3.820441e-15, 3.813068e-15, 3.822208e-15, 
    3.817546e-15, 3.825532e-15, 3.818344e-15, 3.830794e-15, 3.833502e-15, 
    3.831651e-15, 3.838763e-15, 3.817946e-15, 3.825943e-15, 3.765662e-15, 
    3.766017e-15, 3.767673e-15, 3.760392e-15, 3.759947e-15, 3.753275e-15, 
    3.759213e-15, 3.76174e-15, 3.768158e-15, 3.77195e-15, 3.775555e-15, 
    3.783478e-15, 3.792319e-15, 3.804675e-15, 3.813546e-15, 3.819488e-15, 
    3.815846e-15, 3.819062e-15, 3.815466e-15, 3.813781e-15, 3.832487e-15, 
    3.821986e-15, 3.83774e-15, 3.83687e-15, 3.82974e-15, 3.836967e-15, 
    3.766267e-15, 3.764222e-15, 3.757118e-15, 3.762678e-15, 3.752548e-15, 
    3.758218e-15, 3.761476e-15, 3.774047e-15, 3.776811e-15, 3.779369e-15, 
    3.784422e-15, 3.790903e-15, 3.802264e-15, 3.812143e-15, 3.821156e-15, 
    3.820496e-15, 3.820728e-15, 3.82274e-15, 3.817755e-15, 3.823558e-15, 
    3.82453e-15, 3.821986e-15, 3.836753e-15, 3.832536e-15, 3.836851e-15, 
    3.834106e-15, 3.764887e-15, 3.768328e-15, 3.766468e-15, 3.769963e-15, 
    3.7675e-15, 3.778445e-15, 3.781726e-15, 3.797065e-15, 3.790775e-15, 
    3.800788e-15, 3.791793e-15, 3.793387e-15, 3.801109e-15, 3.79228e-15, 
    3.811596e-15, 3.798499e-15, 3.822818e-15, 3.809746e-15, 3.823636e-15, 
    3.821117e-15, 3.825289e-15, 3.829023e-15, 3.833721e-15, 3.842381e-15, 
    3.840377e-15, 3.847617e-15, 3.773456e-15, 3.777913e-15, 3.777523e-15, 
    3.782189e-15, 3.785638e-15, 3.793113e-15, 3.80509e-15, 3.800588e-15, 
    3.808854e-15, 3.810512e-15, 3.797955e-15, 3.805664e-15, 3.780898e-15, 
    3.7849e-15, 3.782519e-15, 3.773806e-15, 3.801622e-15, 3.787353e-15, 
    3.813692e-15, 3.805972e-15, 3.82849e-15, 3.817294e-15, 3.839273e-15, 
    3.848649e-15, 3.857478e-15, 3.867774e-15, 3.780349e-15, 3.77732e-15, 
    3.782745e-15, 3.790242e-15, 3.7972e-15, 3.806442e-15, 3.807389e-15, 
    3.809119e-15, 3.813601e-15, 3.817367e-15, 3.809663e-15, 3.818312e-15, 
    3.785823e-15, 3.802861e-15, 3.776172e-15, 3.784212e-15, 3.789801e-15, 
    3.787352e-15, 3.800074e-15, 3.80307e-15, 3.815235e-15, 3.80895e-15, 
    3.846333e-15, 3.829808e-15, 3.875615e-15, 3.862831e-15, 3.776261e-15, 
    3.780339e-15, 3.79452e-15, 3.787775e-15, 3.80706e-15, 3.811802e-15, 
    3.815657e-15, 3.82058e-15, 3.821113e-15, 3.824028e-15, 3.81925e-15, 
    3.823841e-15, 3.806462e-15, 3.814232e-15, 3.792903e-15, 3.798096e-15, 
    3.795708e-15, 3.793086e-15, 3.801176e-15, 3.809784e-15, 3.809972e-15, 
    3.81273e-15, 3.820493e-15, 3.807139e-15, 3.848458e-15, 3.82295e-15, 
    3.784785e-15, 3.792629e-15, 3.793753e-15, 3.790715e-15, 3.811326e-15, 
    3.803861e-15, 3.823958e-15, 3.818531e-15, 3.827423e-15, 3.823005e-15, 
    3.822354e-15, 3.816678e-15, 3.813142e-15, 3.804203e-15, 3.796927e-15, 
    3.791156e-15, 3.792499e-15, 3.798837e-15, 3.810311e-15, 3.821159e-15, 
    3.818783e-15, 3.826747e-15, 3.805663e-15, 3.814507e-15, 3.811088e-15, 
    3.82e-15, 3.800467e-15, 3.817091e-15, 3.796214e-15, 3.798046e-15, 
    3.803713e-15, 3.815103e-15, 3.817628e-15, 3.820316e-15, 3.818658e-15, 
    3.810603e-15, 3.809285e-15, 3.803576e-15, 3.801998e-15, 3.797648e-15, 
    3.794043e-15, 3.797336e-15, 3.800791e-15, 3.810608e-15, 3.819446e-15, 
    3.829076e-15, 3.831432e-15, 3.842662e-15, 3.833516e-15, 3.848599e-15, 
    3.835769e-15, 3.857973e-15, 3.818059e-15, 3.835399e-15, 3.803972e-15, 
    3.807363e-15, 3.813489e-15, 3.827536e-15, 3.819959e-15, 3.828822e-15, 
    3.809233e-15, 3.799054e-15, 3.796423e-15, 3.791506e-15, 3.796536e-15, 
    3.796127e-15, 3.800938e-15, 3.799392e-15, 3.810934e-15, 3.804736e-15, 
    3.822337e-15, 3.828753e-15, 3.846857e-15, 3.857939e-15, 3.869214e-15, 
    3.874186e-15, 3.8757e-15, 3.876332e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.528752e-09, -8.566361e-09, -8.55905e-09, -8.589383e-09, -8.572558e-09, 
    -8.59242e-09, -8.536378e-09, -8.567853e-09, -8.54776e-09, -8.532139e-09, 
    -8.648252e-09, -8.590738e-09, -8.708009e-09, -8.671323e-09, 
    -8.763486e-09, -8.702298e-09, -8.775825e-09, -8.761723e-09, 
    -8.804172e-09, -8.792011e-09, -8.846304e-09, -8.809785e-09, 
    -8.874453e-09, -8.837584e-09, -8.84335e-09, -8.80858e-09, -8.602314e-09, 
    -8.641091e-09, -8.600016e-09, -8.605545e-09, -8.603064e-09, 
    -8.572904e-09, -8.557705e-09, -8.52588e-09, -8.531657e-09, -8.555033e-09, 
    -8.608032e-09, -8.590042e-09, -8.635385e-09, -8.634362e-09, 
    -8.684844e-09, -8.662082e-09, -8.746938e-09, -8.72282e-09, -8.792519e-09, 
    -8.77499e-09, -8.791694e-09, -8.786629e-09, -8.791761e-09, -8.766053e-09, 
    -8.777067e-09, -8.754446e-09, -8.666344e-09, -8.692234e-09, 
    -8.615018e-09, -8.568589e-09, -8.537758e-09, -8.515879e-09, 
    -8.518971e-09, -8.524868e-09, -8.55517e-09, -8.583663e-09, -8.605377e-09, 
    -8.619902e-09, -8.634214e-09, -8.677532e-09, -8.700465e-09, 
    -8.751814e-09, -8.742549e-09, -8.758247e-09, -8.773245e-09, 
    -8.798426e-09, -8.794282e-09, -8.805375e-09, -8.757834e-09, 
    -8.789429e-09, -8.737271e-09, -8.751536e-09, -8.638098e-09, 
    -8.594895e-09, -8.576527e-09, -8.560455e-09, -8.52135e-09, -8.548354e-09, 
    -8.537708e-09, -8.563037e-09, -8.579131e-09, -8.571171e-09, 
    -8.620299e-09, -8.601199e-09, -8.701824e-09, -8.65848e-09, -8.771496e-09, 
    -8.74445e-09, -8.777978e-09, -8.76087e-09, -8.790185e-09, -8.763802e-09, 
    -8.809504e-09, -8.819456e-09, -8.812655e-09, -8.838781e-09, 
    -8.762339e-09, -8.791694e-09, -8.570948e-09, -8.572246e-09, 
    -8.578295e-09, -8.551708e-09, -8.550082e-09, -8.525721e-09, 
    -8.547397e-09, -8.556628e-09, -8.580065e-09, -8.593926e-09, 
    -8.607103e-09, -8.636078e-09, -8.668437e-09, -8.713689e-09, 
    -8.746204e-09, -8.767999e-09, -8.754635e-09, -8.766434e-09, 
    -8.753243e-09, -8.747062e-09, -8.815727e-09, -8.777169e-09, 
    -8.835023e-09, -8.831822e-09, -8.805639e-09, -8.832183e-09, 
    -8.573158e-09, -8.565688e-09, -8.53975e-09, -8.560049e-09, -8.523068e-09, 
    -8.543767e-09, -8.555668e-09, -8.601597e-09, -8.611689e-09, 
    -8.621046e-09, -8.639528e-09, -8.663247e-09, -8.704856e-09, 
    -8.741063e-09, -8.774118e-09, -8.771696e-09, -8.772549e-09, 
    -8.779933e-09, -8.761642e-09, -8.782935e-09, -8.786509e-09, 
    -8.777166e-09, -8.831393e-09, -8.815901e-09, -8.831754e-09, 
    -8.821667e-09, -8.568116e-09, -8.580686e-09, -8.573894e-09, 
    -8.586666e-09, -8.577667e-09, -8.61768e-09, -8.629677e-09, -8.685819e-09, 
    -8.66278e-09, -8.699449e-09, -8.666505e-09, -8.672342e-09, -8.700643e-09, 
    -8.668286e-09, -8.739065e-09, -8.691075e-09, -8.780219e-09, 
    -8.732291e-09, -8.783223e-09, -8.773975e-09, -8.789288e-09, 
    -8.803001e-09, -8.820255e-09, -8.852089e-09, -8.844718e-09, 
    -8.871343e-09, -8.599426e-09, -8.61573e-09, -8.614296e-09, -8.63136e-09, 
    -8.643979e-09, -8.671333e-09, -8.715206e-09, -8.698708e-09, 
    -8.728997e-09, -8.735078e-09, -8.689062e-09, -8.717313e-09, 
    -8.626643e-09, -8.641289e-09, -8.63257e-09, -8.600712e-09, -8.702508e-09, 
    -8.650264e-09, -8.746741e-09, -8.718437e-09, -8.801045e-09, -8.75996e-09, 
    -8.84066e-09, -8.875157e-09, -8.907632e-09, -8.945579e-09, -8.62463e-09, 
    -8.613552e-09, -8.633389e-09, -8.660834e-09, -8.686303e-09, 
    -8.720162e-09, -8.723628e-09, -8.729971e-09, -8.746403e-09, 
    -8.760218e-09, -8.731975e-09, -8.763681e-09, -8.644684e-09, 
    -8.707043e-09, -8.609362e-09, -8.638772e-09, -8.659216e-09, 
    -8.650249e-09, -8.696823e-09, -8.7078e-09, -8.752406e-09, -8.729347e-09, 
    -8.866642e-09, -8.805896e-09, -8.974476e-09, -8.927361e-09, -8.60968e-09, 
    -8.624593e-09, -8.676492e-09, -8.651798e-09, -8.722424e-09, 
    -8.739809e-09, -8.753942e-09, -8.772009e-09, -8.77396e-09, -8.784665e-09, 
    -8.767123e-09, -8.783972e-09, -8.720234e-09, -8.748717e-09, -8.67056e-09, 
    -8.689581e-09, -8.680832e-09, -8.671233e-09, -8.700858e-09, 
    -8.732419e-09, -8.733096e-09, -8.743216e-09, -8.771731e-09, -8.72271e-09, 
    -8.874478e-09, -8.780743e-09, -8.640853e-09, -8.669574e-09, -8.67368e-09, 
    -8.662553e-09, -8.738065e-09, -8.710703e-09, -8.784403e-09, 
    -8.764485e-09, -8.797122e-09, -8.780904e-09, -8.778517e-09, 
    -8.757689e-09, -8.74472e-09, -8.711957e-09, -8.685302e-09, -8.664167e-09, 
    -8.669081e-09, -8.692298e-09, -8.73435e-09, -8.774136e-09, -8.76542e-09, 
    -8.794641e-09, -8.717302e-09, -8.749731e-09, -8.737196e-09, 
    -8.769879e-09, -8.69827e-09, -8.759242e-09, -8.682684e-09, -8.689397e-09, 
    -8.710161e-09, -8.751928e-09, -8.761172e-09, -8.771039e-09, 
    -8.764951e-09, -8.735419e-09, -8.730581e-09, -8.709656e-09, 
    -8.703878e-09, -8.687935e-09, -8.674736e-09, -8.686795e-09, -8.69946e-09, 
    -8.735432e-09, -8.76785e-09, -8.803196e-09, -8.811847e-09, -8.853142e-09, 
    -8.819523e-09, -8.874999e-09, -8.82783e-09, -8.909488e-09, -8.76278e-09, 
    -8.826446e-09, -8.711106e-09, -8.723531e-09, -8.746005e-09, 
    -8.797554e-09, -8.769726e-09, -8.802272e-09, -8.730392e-09, 
    -8.693099e-09, -8.683452e-09, -8.665451e-09, -8.683864e-09, 
    -8.682367e-09, -8.699986e-09, -8.694323e-09, -8.736626e-09, 
    -8.713903e-09, -8.778457e-09, -8.802015e-09, -8.868551e-09, 
    -8.909342e-09, -8.950868e-09, -8.969202e-09, -8.974783e-09, -8.977115e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.0121e-10, -1.016564e-10, -1.015697e-10, -1.019298e-10, -1.0173e-10, 
    -1.019658e-10, -1.013005e-10, -1.016742e-10, -1.014356e-10, 
    -1.012502e-10, -1.026286e-10, -1.019458e-10, -1.03338e-10, -1.029025e-10, 
    -1.039967e-10, -1.032703e-10, -1.041432e-10, -1.039757e-10, 
    -1.044797e-10, -1.043353e-10, -1.049799e-10, -1.045463e-10, 
    -1.053141e-10, -1.048764e-10, -1.049448e-10, -1.04532e-10, -1.020833e-10, 
    -1.025436e-10, -1.02056e-10, -1.021216e-10, -1.020922e-10, -1.017341e-10, 
    -1.015537e-10, -1.011759e-10, -1.012445e-10, -1.01522e-10, -1.021511e-10, 
    -1.019376e-10, -1.024759e-10, -1.024637e-10, -1.03063e-10, -1.027928e-10, 
    -1.038002e-10, -1.035139e-10, -1.043413e-10, -1.041332e-10, 
    -1.043316e-10, -1.042714e-10, -1.043323e-10, -1.040271e-10, 
    -1.041579e-10, -1.038893e-10, -1.028434e-10, -1.031508e-10, 
    -1.022341e-10, -1.016829e-10, -1.013169e-10, -1.010571e-10, 
    -1.010939e-10, -1.011639e-10, -1.015236e-10, -1.018618e-10, 
    -1.021196e-10, -1.022921e-10, -1.02462e-10, -1.029762e-10, -1.032485e-10, 
    -1.038581e-10, -1.037481e-10, -1.039345e-10, -1.041125e-10, 
    -1.044115e-10, -1.043623e-10, -1.04494e-10, -1.039296e-10, -1.043047e-10, 
    -1.036854e-10, -1.038548e-10, -1.025081e-10, -1.019952e-10, 
    -1.017771e-10, -1.015863e-10, -1.011221e-10, -1.014427e-10, 
    -1.013163e-10, -1.01617e-10, -1.01808e-10, -1.017136e-10, -1.022968e-10, 
    -1.0207e-10, -1.032646e-10, -1.0275e-10, -1.040918e-10, -1.037707e-10, 
    -1.041687e-10, -1.039656e-10, -1.043136e-10, -1.040004e-10, -1.04543e-10, 
    -1.046612e-10, -1.045804e-10, -1.048906e-10, -1.039831e-10, 
    -1.043316e-10, -1.017109e-10, -1.017263e-10, -1.017981e-10, 
    -1.014825e-10, -1.014632e-10, -1.01174e-10, -1.014313e-10, -1.015409e-10, 
    -1.018191e-10, -1.019837e-10, -1.021401e-10, -1.024841e-10, 
    -1.028682e-10, -1.034055e-10, -1.037915e-10, -1.040502e-10, 
    -1.038916e-10, -1.040317e-10, -1.038751e-10, -1.038017e-10, 
    -1.046169e-10, -1.041591e-10, -1.04846e-10, -1.04808e-10, -1.044971e-10, 
    -1.048123e-10, -1.017371e-10, -1.016485e-10, -1.013405e-10, 
    -1.015815e-10, -1.011425e-10, -1.013882e-10, -1.015295e-10, 
    -1.020747e-10, -1.021946e-10, -1.023056e-10, -1.025251e-10, 
    -1.028066e-10, -1.033006e-10, -1.037305e-10, -1.041229e-10, 
    -1.040941e-10, -1.041043e-10, -1.041919e-10, -1.039748e-10, 
    -1.042276e-10, -1.0427e-10, -1.041591e-10, -1.048029e-10, -1.046189e-10, 
    -1.048072e-10, -1.046874e-10, -1.016773e-10, -1.018265e-10, 
    -1.017459e-10, -1.018975e-10, -1.017907e-10, -1.022657e-10, 
    -1.024081e-10, -1.030746e-10, -1.028011e-10, -1.032364e-10, 
    -1.028453e-10, -1.029146e-10, -1.032506e-10, -1.028665e-10, 
    -1.037067e-10, -1.03137e-10, -1.041953e-10, -1.036263e-10, -1.04231e-10, 
    -1.041212e-10, -1.04303e-10, -1.044658e-10, -1.046706e-10, -1.050486e-10, 
    -1.049611e-10, -1.052772e-10, -1.02049e-10, -1.022425e-10, -1.022255e-10, 
    -1.024281e-10, -1.025779e-10, -1.029026e-10, -1.034235e-10, 
    -1.032276e-10, -1.035872e-10, -1.036594e-10, -1.031131e-10, 
    -1.034485e-10, -1.023721e-10, -1.02546e-10, -1.024425e-10, -1.020642e-10, 
    -1.032727e-10, -1.026525e-10, -1.037979e-10, -1.034618e-10, 
    -1.044426e-10, -1.039548e-10, -1.049129e-10, -1.053225e-10, -1.05708e-10, 
    -1.061586e-10, -1.023482e-10, -1.022167e-10, -1.024522e-10, -1.02778e-10, 
    -1.030804e-10, -1.034823e-10, -1.035235e-10, -1.035988e-10, 
    -1.037939e-10, -1.039579e-10, -1.036226e-10, -1.03999e-10, -1.025863e-10, 
    -1.033266e-10, -1.021669e-10, -1.025161e-10, -1.027588e-10, 
    -1.026523e-10, -1.032052e-10, -1.033356e-10, -1.038651e-10, 
    -1.035914e-10, -1.052214e-10, -1.045002e-10, -1.065017e-10, 
    -1.059423e-10, -1.021707e-10, -1.023477e-10, -1.029639e-10, 
    -1.026707e-10, -1.035092e-10, -1.037156e-10, -1.038834e-10, 
    -1.040978e-10, -1.04121e-10, -1.042481e-10, -1.040399e-10, -1.042399e-10, 
    -1.034832e-10, -1.038213e-10, -1.028935e-10, -1.031193e-10, 
    -1.030154e-10, -1.029014e-10, -1.032531e-10, -1.036278e-10, 
    -1.036359e-10, -1.03756e-10, -1.040946e-10, -1.035126e-10, -1.053144e-10, 
    -1.042016e-10, -1.025408e-10, -1.028818e-10, -1.029305e-10, 
    -1.027984e-10, -1.036949e-10, -1.0337e-10, -1.04245e-10, -1.040085e-10, 
    -1.04396e-10, -1.042035e-10, -1.041751e-10, -1.039278e-10, -1.037739e-10, 
    -1.033849e-10, -1.030685e-10, -1.028176e-10, -1.028759e-10, 
    -1.031515e-10, -1.036508e-10, -1.041231e-10, -1.040196e-10, 
    -1.043666e-10, -1.034484e-10, -1.038334e-10, -1.036846e-10, 
    -1.040726e-10, -1.032224e-10, -1.039463e-10, -1.030374e-10, 
    -1.031171e-10, -1.033636e-10, -1.038595e-10, -1.039692e-10, 
    -1.040863e-10, -1.040141e-10, -1.036635e-10, -1.03606e-10, -1.033576e-10, 
    -1.03289e-10, -1.030997e-10, -1.02943e-10, -1.030862e-10, -1.032366e-10, 
    -1.036636e-10, -1.040485e-10, -1.044681e-10, -1.045708e-10, 
    -1.050611e-10, -1.04662e-10, -1.053206e-10, -1.047606e-10, -1.057301e-10, 
    -1.039883e-10, -1.047442e-10, -1.033748e-10, -1.035223e-10, 
    -1.037891e-10, -1.044011e-10, -1.040708e-10, -1.044571e-10, 
    -1.036038e-10, -1.03161e-10, -1.030465e-10, -1.028328e-10, -1.030514e-10, 
    -1.030336e-10, -1.032428e-10, -1.031756e-10, -1.036778e-10, -1.03408e-10, 
    -1.041744e-10, -1.044541e-10, -1.05244e-10, -1.057283e-10, -1.062214e-10, 
    -1.06439e-10, -1.065053e-10, -1.06533e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.393943e-12, -8.430986e-12, -8.423785e-12, -8.453663e-12, -8.43709e-12, 
    -8.456654e-12, -8.401453e-12, -8.432456e-12, -8.412665e-12, 
    -8.397279e-12, -8.511647e-12, -8.454997e-12, -8.570507e-12, 
    -8.534372e-12, -8.625153e-12, -8.564883e-12, -8.637306e-12, 
    -8.623416e-12, -8.665228e-12, -8.653249e-12, -8.706728e-12, 
    -8.670757e-12, -8.734456e-12, -8.698139e-12, -8.703819e-12, -8.66957e-12, 
    -8.466399e-12, -8.504594e-12, -8.464136e-12, -8.469582e-12, 
    -8.467138e-12, -8.437431e-12, -8.42246e-12, -8.391112e-12, -8.396804e-12, 
    -8.419828e-12, -8.472031e-12, -8.454312e-12, -8.498974e-12, 
    -8.497965e-12, -8.54769e-12, -8.52527e-12, -8.608852e-12, -8.585096e-12, 
    -8.65375e-12, -8.636483e-12, -8.652938e-12, -8.647949e-12, -8.653003e-12, 
    -8.62768e-12, -8.638529e-12, -8.616248e-12, -8.529468e-12, -8.55497e-12, 
    -8.478913e-12, -8.433181e-12, -8.402813e-12, -8.381263e-12, 
    -8.384309e-12, -8.390117e-12, -8.419964e-12, -8.448028e-12, 
    -8.469416e-12, -8.483723e-12, -8.497821e-12, -8.540489e-12, 
    -8.563077e-12, -8.613656e-12, -8.604529e-12, -8.619991e-12, 
    -8.634766e-12, -8.659568e-12, -8.655486e-12, -8.666413e-12, 
    -8.619585e-12, -8.650706e-12, -8.59933e-12, -8.613382e-12, -8.501646e-12, 
    -8.459092e-12, -8.441e-12, -8.425169e-12, -8.386652e-12, -8.41325e-12, 
    -8.402765e-12, -8.427713e-12, -8.443564e-12, -8.435724e-12, 
    -8.484114e-12, -8.465301e-12, -8.564416e-12, -8.521722e-12, 
    -8.633042e-12, -8.606403e-12, -8.639428e-12, -8.622576e-12, -8.65145e-12, 
    -8.625464e-12, -8.670481e-12, -8.680283e-12, -8.673584e-12, 
    -8.699318e-12, -8.624023e-12, -8.652938e-12, -8.435505e-12, 
    -8.436783e-12, -8.44274e-12, -8.416553e-12, -8.414952e-12, -8.390956e-12, 
    -8.412308e-12, -8.4214e-12, -8.444484e-12, -8.458137e-12, -8.471117e-12, 
    -8.499656e-12, -8.531529e-12, -8.576103e-12, -8.60813e-12, -8.629598e-12, 
    -8.616434e-12, -8.628056e-12, -8.615064e-12, -8.608975e-12, -8.67661e-12, 
    -8.638631e-12, -8.695617e-12, -8.692464e-12, -8.666673e-12, 
    -8.692819e-12, -8.437681e-12, -8.430323e-12, -8.404775e-12, 
    -8.424769e-12, -8.388344e-12, -8.408731e-12, -8.420454e-12, 
    -8.465693e-12, -8.475634e-12, -8.48485e-12, -8.503055e-12, -8.526417e-12, 
    -8.567402e-12, -8.603066e-12, -8.635625e-12, -8.63324e-12, -8.63408e-12, 
    -8.641352e-12, -8.623336e-12, -8.64431e-12, -8.64783e-12, -8.638626e-12, 
    -8.692042e-12, -8.676782e-12, -8.692397e-12, -8.682461e-12, 
    -8.432715e-12, -8.445096e-12, -8.438406e-12, -8.450986e-12, 
    -8.442123e-12, -8.481535e-12, -8.493352e-12, -8.548651e-12, 
    -8.525957e-12, -8.562076e-12, -8.529627e-12, -8.535376e-12, 
    -8.563252e-12, -8.53138e-12, -8.601098e-12, -8.553829e-12, -8.641635e-12, 
    -8.594426e-12, -8.644594e-12, -8.635485e-12, -8.650567e-12, 
    -8.664075e-12, -8.68107e-12, -8.712427e-12, -8.705166e-12, -8.731391e-12, 
    -8.463555e-12, -8.479614e-12, -8.478202e-12, -8.495009e-12, 
    -8.507439e-12, -8.534382e-12, -8.577597e-12, -8.561346e-12, 
    -8.591182e-12, -8.597171e-12, -8.551845e-12, -8.579673e-12, 
    -8.490363e-12, -8.50479e-12, -8.496201e-12, -8.464821e-12, -8.565089e-12, 
    -8.513629e-12, -8.608658e-12, -8.580778e-12, -8.662148e-12, -8.62168e-12, 
    -8.701169e-12, -8.735149e-12, -8.767138e-12, -8.804515e-12, -8.48838e-12, 
    -8.477468e-12, -8.497008e-12, -8.524041e-12, -8.549128e-12, 
    -8.582478e-12, -8.585892e-12, -8.59214e-12, -8.608326e-12, -8.621934e-12, 
    -8.594114e-12, -8.625345e-12, -8.508133e-12, -8.569557e-12, 
    -8.473341e-12, -8.502311e-12, -8.522448e-12, -8.513615e-12, 
    -8.559489e-12, -8.570302e-12, -8.614239e-12, -8.591526e-12, 
    -8.726761e-12, -8.666926e-12, -8.83298e-12, -8.78657e-12, -8.473655e-12, 
    -8.488343e-12, -8.539463e-12, -8.51514e-12, -8.584706e-12, -8.60183e-12, 
    -8.615752e-12, -8.633547e-12, -8.635469e-12, -8.646013e-12, 
    -8.628735e-12, -8.645331e-12, -8.58255e-12, -8.610605e-12, -8.533622e-12, 
    -8.552357e-12, -8.543739e-12, -8.534284e-12, -8.563464e-12, 
    -8.594551e-12, -8.595218e-12, -8.605186e-12, -8.633273e-12, 
    -8.584988e-12, -8.73448e-12, -8.64215e-12, -8.50436e-12, -8.53265e-12, 
    -8.536694e-12, -8.525734e-12, -8.600113e-12, -8.573162e-12, 
    -8.645757e-12, -8.626136e-12, -8.658284e-12, -8.642309e-12, 
    -8.639959e-12, -8.619442e-12, -8.606668e-12, -8.574397e-12, 
    -8.548141e-12, -8.527324e-12, -8.532165e-12, -8.555033e-12, 
    -8.596454e-12, -8.635643e-12, -8.627057e-12, -8.655841e-12, 
    -8.579662e-12, -8.611603e-12, -8.599257e-12, -8.63145e-12, -8.560914e-12, 
    -8.620973e-12, -8.545563e-12, -8.552175e-12, -8.572627e-12, 
    -8.613768e-12, -8.622874e-12, -8.632592e-12, -8.626596e-12, 
    -8.597506e-12, -8.592741e-12, -8.57213e-12, -8.566438e-12, -8.550735e-12, 
    -8.537733e-12, -8.549612e-12, -8.562087e-12, -8.597519e-12, -8.62945e-12, 
    -8.664266e-12, -8.672788e-12, -8.713465e-12, -8.680349e-12, 
    -8.734994e-12, -8.688532e-12, -8.768966e-12, -8.624456e-12, 
    -8.687169e-12, -8.573559e-12, -8.585797e-12, -8.607933e-12, 
    -8.658709e-12, -8.631299e-12, -8.663356e-12, -8.592555e-12, 
    -8.555821e-12, -8.54632e-12, -8.528589e-12, -8.546725e-12, -8.54525e-12, 
    -8.562605e-12, -8.557027e-12, -8.598696e-12, -8.576313e-12, -8.6399e-12, 
    -8.663104e-12, -8.728643e-12, -8.768822e-12, -8.809726e-12, 
    -8.827786e-12, -8.833282e-12, -8.83558e-12 ;

 SMIN_NH4 =
  0.000435042, 0.0004368748, 0.0004365185, 0.0004379967, 0.0004371766, 
    0.0004381445, 0.0004354134, 0.0004369472, 0.000435968, 0.0004352066, 
    0.0004408649, 0.0004380622, 0.0004437764, 0.0004419888, 0.0004464791, 
    0.000443498, 0.0004470801, 0.000446393, 0.000448461, 0.0004478684, 
    0.0004505132, 0.0004487342, 0.0004518842, 0.0004500883, 0.0004503691, 
    0.0004486753, 0.0004386267, 0.0004405163, 0.0004385146, 0.0004387841, 
    0.0004386631, 0.0004371933, 0.0004364526, 0.0004349015, 0.000435183, 
    0.0004363222, 0.0004389049, 0.0004380281, 0.0004402376, 0.0004401877, 
    0.0004426474, 0.0004415383, 0.0004456727, 0.0004444975, 0.0004478931, 
    0.0004470391, 0.0004478529, 0.000447606, 0.0004478559, 0.0004466035, 
    0.00044714, 0.000446038, 0.0004417467, 0.0004430081, 0.0004392456, 
    0.000436983, 0.0004354804, 0.0004344141, 0.0004345647, 0.0004348521, 
    0.0004363288, 0.0004377172, 0.0004387753, 0.000439483, 0.0004401804, 
    0.0004422911, 0.0004434084, 0.0004459101, 0.0004454587, 0.0004462234, 
    0.000446954, 0.0004481807, 0.0004479787, 0.0004485191, 0.0004462029, 
    0.0004477422, 0.000445201, 0.000445896, 0.0004403702, 0.0004382649, 
    0.0004373698, 0.0004365864, 0.0004346806, 0.0004359967, 0.0004354778, 
    0.0004367121, 0.0004374963, 0.0004371084, 0.0004395023, 0.0004385715, 
    0.0004434746, 0.0004413627, 0.0004468689, 0.0004455512, 0.0004471845, 
    0.0004463511, 0.000447779, 0.0004464938, 0.0004487201, 0.0004492049, 
    0.0004488735, 0.0004501462, 0.0004464222, 0.0004478523, 0.0004370978, 
    0.0004371611, 0.0004374557, 0.00043616, 0.0004360808, 0.0004348934, 
    0.0004359498, 0.0004363997, 0.0004375417, 0.0004382171, 0.0004388591, 
    0.000440271, 0.0004418477, 0.0004440525, 0.0004456365, 0.0004466983, 
    0.0004460472, 0.0004466219, 0.0004459793, 0.0004456781, 0.0004490231, 
    0.0004471448, 0.000449963, 0.0004498071, 0.0004485315, 0.0004498245, 
    0.0004372054, 0.0004368413, 0.0004355772, 0.0004365663, 0.000434764, 
    0.0004357728, 0.0004363528, 0.0004385908, 0.0004390826, 0.0004395385, 
    0.000440439, 0.0004415947, 0.000443622, 0.000445386, 0.0004469963, 
    0.0004468783, 0.0004469198, 0.0004472794, 0.0004463883, 0.0004474256, 
    0.0004475996, 0.0004471444, 0.000449786, 0.0004490313, 0.0004498035, 
    0.0004493121, 0.0004369596, 0.000437572, 0.0004372409, 0.0004378634, 
    0.0004374247, 0.0004393746, 0.0004399591, 0.0004426946, 0.0004415719, 
    0.0004433586, 0.0004417533, 0.0004420377, 0.0004434166, 0.0004418399, 
    0.0004452885, 0.0004429503, 0.0004472933, 0.0004449583, 0.0004474396, 
    0.0004469889, 0.0004477348, 0.0004484029, 0.0004492433, 0.000450794, 
    0.0004504348, 0.0004517318, 0.0004384852, 0.0004392796, 0.0004392097, 
    0.000440041, 0.0004406559, 0.0004419888, 0.0004441263, 0.0004433224, 
    0.0004447981, 0.0004450943, 0.0004428522, 0.0004442287, 0.0004398108, 
    0.0004405244, 0.0004400995, 0.000438547, 0.0004435071, 0.0004409614, 
    0.0004456621, 0.000444283, 0.0004483075, 0.000446306, 0.0004502371, 
    0.0004519175, 0.0004534992, 0.0004553474, 0.0004397132, 0.0004391733, 
    0.0004401398, 0.0004414772, 0.000442718, 0.0004443677, 0.0004445365, 
    0.0004448454, 0.0004456459, 0.000446319, 0.000444943, 0.0004464876, 
    0.0004406898, 0.0004437281, 0.0004389684, 0.0004404015, 0.0004413976, 
    0.0004409607, 0.0004432299, 0.0004437646, 0.0004459378, 0.0004448144, 
    0.0004515026, 0.0004485435, 0.0004567546, 0.00045446, 0.0004389846, 
    0.0004397111, 0.0004422399, 0.0004410367, 0.0004444777, 0.0004453248, 
    0.0004460132, 0.0004468934, 0.0004469883, 0.0004475098, 0.0004466551, 
    0.000447476, 0.0004443707, 0.0004457583, 0.0004419503, 0.000442877, 
    0.0004424507, 0.0004419829, 0.0004434263, 0.000444964, 0.0004449969, 
    0.0004454899, 0.000446879, 0.0004444907, 0.0004518841, 0.0004473179, 
    0.0004405034, 0.0004419028, 0.0004421028, 0.0004415606, 0.0004452397, 
    0.0004439066, 0.0004474971, 0.0004465267, 0.0004481166, 0.0004473265, 
    0.0004472101, 0.0004461954, 0.0004455634, 0.0004439673, 0.0004426684, 
    0.0004416386, 0.000441878, 0.0004430092, 0.0004450579, 0.0004469962, 
    0.0004465716, 0.000447995, 0.0004442271, 0.000445807, 0.0004451962, 
    0.0004467885, 0.0004433008, 0.0004462715, 0.0004425414, 0.0004428684, 
    0.00044388, 0.0004459149, 0.0004463652, 0.0004468459, 0.0004465492, 
    0.0004451104, 0.0004448746, 0.000443855, 0.0004435734, 0.0004427967, 
    0.0004421534, 0.000442741, 0.0004433579, 0.0004451106, 0.0004466899, 
    0.0004484117, 0.0004488331, 0.0004508447, 0.000449207, 0.0004519093, 
    0.0004496115, 0.000453589, 0.0004464436, 0.0004495452, 0.0004439261, 
    0.0004445314, 0.0004456262, 0.0004481375, 0.0004467817, 0.0004483673, 
    0.0004448653, 0.0004430483, 0.0004425782, 0.0004417012, 0.0004425982, 
    0.0004425252, 0.0004433836, 0.0004431076, 0.0004451686, 0.0004440615, 
    0.0004472064, 0.0004483541, 0.0004515952, 0.0004535819, 0.0004556045, 
    0.0004564972, 0.000456769, 0.0004568826 ;

 SMIN_NH4_vr =
  0.002842044, 0.002846979, 0.002846014, 0.002849991, 0.002847782, 
    0.00285038, 0.00284303, 0.002847152, 0.002844517, 0.002842463, 
    0.002857672, 0.002850143, 0.002865491, 0.002860689, 0.002872731, 
    0.002864735, 0.002874339, 0.002872495, 0.002878035, 0.002876444, 
    0.002883517, 0.00287876, 0.00288718, 0.002882377, 0.002883123, 
    0.002878587, 0.002851683, 0.002856757, 0.002851376, 0.002852101, 
    0.002851772, 0.002847813, 0.002845817, 0.00284164, 0.002842393, 
    0.00284546, 0.002852404, 0.002850043, 0.00285598, 0.002855846, 
    0.002862446, 0.002859469, 0.00287056, 0.002867404, 0.002876506, 
    0.002874213, 0.002876392, 0.002875727, 0.002876392, 0.002873036, 
    0.002874468, 0.002871515, 0.002860063, 0.002863445, 0.002853336, 
    0.002847242, 0.002843197, 0.002840327, 0.002840726, 0.0028415, 
    0.002845471, 0.002849204, 0.002852049, 0.002853947, 0.002855818, 
    0.002861483, 0.002864481, 0.002871189, 0.002869979, 0.002872023, 
    0.002873982, 0.002877264, 0.002876722, 0.002878164, 0.002871954, 
    0.002876079, 0.002869262, 0.002871126, 0.00285635, 0.002850693, 
    0.00284828, 0.00284617, 0.002841036, 0.00284458, 0.002843179, 
    0.002846498, 0.002848607, 0.002847559, 0.002853996, 0.002851488, 
    0.002864654, 0.002858985, 0.002873757, 0.00287022, 0.002874595, 
    0.002872362, 0.002876181, 0.002872739, 0.002878697, 0.002879994, 
    0.002879101, 0.002882509, 0.002872528, 0.00287636, 0.002847547, 
    0.002847718, 0.002848507, 0.002845014, 0.0028448, 0.002841599, 
    0.00284444, 0.002845651, 0.002848721, 0.002850533, 0.002852255, 
    0.002856051, 0.002860282, 0.002866196, 0.002870446, 0.002873288, 
    0.002871542, 0.002873078, 0.002871353, 0.002870541, 0.002879499, 
    0.002874468, 0.00288201, 0.002881594, 0.002878174, 0.002881632, 
    0.002847831, 0.002846847, 0.002843443, 0.002846102, 0.002841245, 
    0.002843961, 0.002845517, 0.002851534, 0.002852855, 0.00285408, 
    0.002856497, 0.002859597, 0.002865038, 0.002869766, 0.002874084, 
    0.002873763, 0.002873873, 0.002874831, 0.002872442, 0.002875217, 
    0.002875679, 0.002874461, 0.002881529, 0.002879509, 0.002881573, 
    0.002880253, 0.002847162, 0.002848805, 0.002847911, 0.002849585, 
    0.002848399, 0.002853642, 0.002855209, 0.002862552, 0.002859535, 
    0.002864333, 0.002860017, 0.002860781, 0.002864475, 0.002860243, 
    0.002869494, 0.002863214, 0.002874865, 0.002868596, 0.002875251, 
    0.00287404, 0.002876034, 0.002877824, 0.002880068, 0.002884218, 
    0.002883251, 0.002886721, 0.002851258, 0.002853388, 0.002853201, 
    0.002855431, 0.002857079, 0.00286066, 0.002866394, 0.002864233, 
    0.002868189, 0.002868983, 0.002862961, 0.002866654, 0.002854786, 
    0.002856698, 0.002855557, 0.002851378, 0.002864701, 0.00285786, 
    0.002870478, 0.002866775, 0.002877559, 0.002872195, 0.00288272, 
    0.002887212, 0.00289144, 0.002896368, 0.002854552, 0.002853096, 
    0.002855691, 0.002859282, 0.002862609, 0.002867038, 0.002867487, 
    0.002868311, 0.002870455, 0.00287226, 0.002868564, 0.002872703, 
    0.002857135, 0.002865294, 0.002852505, 0.002856356, 0.002859027, 
    0.002857855, 0.002863946, 0.002865376, 0.0028712, 0.00286819, 
    0.002886093, 0.002878176, 0.00290012, 0.002893994, 0.002852585, 
    0.002854534, 0.002861323, 0.002858093, 0.002867325, 0.002869597, 
    0.002871437, 0.002873796, 0.002874045, 0.002875443, 0.002873146, 
    0.002875347, 0.002867013, 0.002870737, 0.002860514, 0.002862997, 
    0.002861852, 0.002860591, 0.002864462, 0.002868586, 0.002868673, 
    0.002869989, 0.002873705, 0.002867305, 0.002887098, 0.002874871, 
    0.00285666, 0.002860412, 0.002860948, 0.002859493, 0.00286936, 
    0.002865785, 0.002875409, 0.002872804, 0.00287706, 0.002874944, 
    0.002874625, 0.002871907, 0.002870205, 0.002865923, 0.002862431, 
    0.002859667, 0.002860304, 0.00286334, 0.00286883, 0.002874029, 
    0.002872886, 0.002876698, 0.002866592, 0.002870829, 0.002869184, 
    0.002873455, 0.002864162, 0.002872124, 0.002862121, 0.002862994, 
    0.002865704, 0.002871161, 0.002872365, 0.002873653, 0.002872852, 
    0.002868993, 0.002868358, 0.002865619, 0.002864858, 0.002862775, 
    0.002861041, 0.002862619, 0.002864267, 0.002868972, 0.002873201, 
    0.002877811, 0.002878939, 0.002884313, 0.002879929, 0.00288715, 
    0.002881001, 0.002891637, 0.00287258, 0.002880889, 0.00286583, 
    0.002867449, 0.002870382, 0.002877107, 0.002873473, 0.00287772, 
    0.002868331, 0.002863449, 0.002862185, 0.002859831, 0.002862233, 
    0.002862038, 0.002864338, 0.002863593, 0.002869118, 0.00286615, 
    0.002874576, 0.00287765, 0.002886321, 0.002891626, 0.002897029, 
    0.002899407, 0.002900131, 0.00290043,
  0.001592138, 0.001598168, 0.001596997, 0.001601856, 0.001599161, 
    0.001602342, 0.001593362, 0.001598407, 0.001595187, 0.001592682, 
    0.001611274, 0.001602073, 0.001620824, 0.001614965, 0.001629674, 
    0.001619912, 0.001631641, 0.001629394, 0.001636157, 0.00163422, 
    0.001642859, 0.001637051, 0.001647335, 0.001641473, 0.00164239, 
    0.001636859, 0.001603927, 0.001610129, 0.001603559, 0.001604444, 
    0.001604047, 0.001599217, 0.00159678, 0.001591678, 0.001592605, 
    0.001596352, 0.001604842, 0.001601962, 0.00160922, 0.001609056, 
    0.001617125, 0.001613489, 0.001627037, 0.001623189, 0.001634301, 
    0.001631508, 0.00163417, 0.001633363, 0.00163418, 0.001630084, 
    0.001631839, 0.001628234, 0.00161417, 0.001618306, 0.001605961, 
    0.001598524, 0.001593583, 0.001590073, 0.00159057, 0.001591515, 
    0.001596374, 0.001600941, 0.001604418, 0.001606743, 0.001609033, 
    0.001615955, 0.001619619, 0.001627813, 0.001626337, 0.001628839, 
    0.001631231, 0.001635242, 0.001634582, 0.001636348, 0.001628774, 
    0.001633808, 0.001625495, 0.00162777, 0.00160965, 0.00160274, 
    0.001599796, 0.001597222, 0.001590951, 0.001595282, 0.001593575, 
    0.001597636, 0.001600215, 0.00159894, 0.001606806, 0.001603749, 
    0.001619837, 0.001612912, 0.001630952, 0.00162664, 0.001631985, 
    0.001629258, 0.001633929, 0.001629726, 0.001637006, 0.001638589, 
    0.001637507, 0.001641665, 0.001629492, 0.001634169, 0.001598904, 
    0.001599112, 0.001600081, 0.001595819, 0.001595559, 0.001591652, 
    0.001595129, 0.001596608, 0.001600364, 0.001602584, 0.001604694, 
    0.00160933, 0.001614503, 0.001621731, 0.00162692, 0.001630395, 
    0.001628264, 0.001630145, 0.001628042, 0.001627057, 0.001637996, 
    0.001631855, 0.001641067, 0.001640558, 0.00163639, 0.001640615, 
    0.001599258, 0.001598061, 0.001593902, 0.001597157, 0.001591227, 
    0.001594546, 0.001596454, 0.001603812, 0.001605428, 0.001606926, 
    0.001609882, 0.001613675, 0.001620321, 0.001626099, 0.00163137, 
    0.001630984, 0.00163112, 0.001632296, 0.001629381, 0.001632775, 
    0.001633343, 0.001631855, 0.001640489, 0.001638024, 0.001640547, 
    0.001638942, 0.00159845, 0.001600464, 0.001599376, 0.001601421, 
    0.00159998, 0.001606386, 0.001608305, 0.00161728, 0.0016136, 0.001619458, 
    0.001614196, 0.001615128, 0.001619647, 0.00161448, 0.00162578, 
    0.00161812, 0.001632342, 0.001624698, 0.00163282, 0.001631347, 
    0.001633787, 0.00163597, 0.001638717, 0.00164378, 0.001642608, 
    0.001646841, 0.001603465, 0.001606074, 0.001605846, 0.001608576, 
    0.001610594, 0.001614967, 0.001621974, 0.00161934, 0.001624175, 
    0.001625145, 0.0016178, 0.00162231, 0.001607821, 0.001610163, 
    0.001608769, 0.00160367, 0.001619946, 0.001611598, 0.001627005, 
    0.00162249, 0.001635659, 0.001629112, 0.001641963, 0.001647446, 
    0.001652605, 0.001658624, 0.001607499, 0.001605726, 0.001608901, 
    0.001613288, 0.001617359, 0.001622765, 0.001623318, 0.00162433, 
    0.001626952, 0.001629154, 0.001624649, 0.001629706, 0.001610704, 
    0.00162067, 0.001605055, 0.00160976, 0.00161303, 0.001611597, 
    0.001619039, 0.001620792, 0.001627908, 0.001624231, 0.001646092, 
    0.00163643, 0.001663206, 0.001655735, 0.001605107, 0.001607493, 
    0.001615791, 0.001611844, 0.001623126, 0.001625899, 0.001628154, 
    0.001631033, 0.001631345, 0.00163305, 0.001630255, 0.00163294, 
    0.001622776, 0.00162732, 0.001614844, 0.001617883, 0.001616485, 
    0.001614951, 0.001619684, 0.00162472, 0.001624829, 0.001626443, 
    0.001630985, 0.001623172, 0.001647335, 0.001632421, 0.001610095, 
    0.001614685, 0.001615342, 0.001613564, 0.001625621, 0.001621255, 
    0.001633008, 0.001629835, 0.001635034, 0.001632451, 0.001632071, 
    0.001628751, 0.001626683, 0.001621455, 0.001617199, 0.001613822, 
    0.001614608, 0.001618316, 0.001625028, 0.001631372, 0.001629983, 
    0.001634639, 0.001622309, 0.001627482, 0.001625482, 0.001630694, 
    0.00161927, 0.001628995, 0.001616781, 0.001617853, 0.001621169, 
    0.001627831, 0.001629306, 0.001630879, 0.001629909, 0.001625199, 
    0.001624427, 0.001621088, 0.001620165, 0.00161762, 0.001615511, 
    0.001617438, 0.00161946, 0.001625201, 0.00163037, 0.001636001, 
    0.001637379, 0.001643946, 0.001638598, 0.001647418, 0.001639917, 
    0.001652897, 0.00162956, 0.0016397, 0.00162132, 0.001623303, 0.001626887, 
    0.001635102, 0.00163067, 0.001635853, 0.001624397, 0.001618443, 
    0.001616904, 0.001614027, 0.00161697, 0.00161673, 0.001619544, 
    0.00161864, 0.001625392, 0.001621766, 0.001632061, 0.001635813, 
    0.001646397, 0.001652875, 0.001659465, 0.001662371, 0.001663255, 
    0.001663624,
  0.001500654, 0.00150729, 0.001506, 0.001511349, 0.001508383, 0.001511885, 
    0.001502, 0.001507553, 0.001504009, 0.001501252, 0.001521721, 
    0.001511588, 0.001532239, 0.001525784, 0.001541992, 0.001531234, 
    0.00154416, 0.001541683, 0.001549138, 0.001547003, 0.001556531, 
    0.001550124, 0.001561468, 0.001555002, 0.001556013, 0.001549912, 
    0.001513629, 0.00152046, 0.001513224, 0.001514198, 0.001513761, 
    0.001508444, 0.001505762, 0.001500147, 0.001501167, 0.001505291, 
    0.001514636, 0.001511466, 0.001519456, 0.001519276, 0.001528163, 
    0.001524157, 0.001539084, 0.001534844, 0.001547092, 0.001544013, 
    0.001546948, 0.001546058, 0.001546959, 0.001542443, 0.001544378, 
    0.001540404, 0.001524907, 0.001529464, 0.001515868, 0.001507682, 
    0.001502244, 0.001498382, 0.001498928, 0.001499969, 0.001505316, 
    0.001510341, 0.001514169, 0.001516728, 0.00151925, 0.001526876, 
    0.001530912, 0.001539941, 0.001538313, 0.001541071, 0.001543707, 
    0.001548129, 0.001547402, 0.00154935, 0.001540999, 0.001546549, 
    0.001537385, 0.001539892, 0.001519933, 0.001512321, 0.001509082, 
    0.001506248, 0.001499348, 0.001504113, 0.001502235, 0.001506704, 
    0.001509542, 0.001508138, 0.001516798, 0.001513432, 0.001531151, 
    0.001523523, 0.0015434, 0.001538647, 0.001544539, 0.001541533, 
    0.001546682, 0.001542048, 0.001550074, 0.001551821, 0.001550628, 
    0.001555212, 0.001541791, 0.001546947, 0.001508099, 0.001508328, 
    0.001509394, 0.001504705, 0.001504418, 0.001500119, 0.001503945, 
    0.001505573, 0.001509706, 0.00151215, 0.001514473, 0.001519578, 
    0.001525276, 0.001533238, 0.001538955, 0.001542785, 0.001540437, 
    0.00154251, 0.001540193, 0.001539106, 0.001551166, 0.001544396, 
    0.001554553, 0.001553991, 0.001549396, 0.001554055, 0.001508489, 
    0.001507171, 0.001502595, 0.001506176, 0.001499651, 0.001503304, 
    0.001505403, 0.001513502, 0.001515281, 0.00151693, 0.001520186, 
    0.001524362, 0.001531685, 0.001538051, 0.00154386, 0.001543435, 
    0.001543585, 0.001544882, 0.001541668, 0.001545409, 0.001546037, 
    0.001544396, 0.001553916, 0.001551197, 0.001553979, 0.001552209, 
    0.001507599, 0.001509816, 0.001508618, 0.00151087, 0.001509284, 
    0.001516336, 0.00151845, 0.001528335, 0.00152428, 0.001530733, 
    0.001524936, 0.001525963, 0.001530943, 0.001525249, 0.0015377, 
    0.00152926, 0.001544932, 0.001536509, 0.00154546, 0.001543835, 
    0.001546525, 0.001548933, 0.001551961, 0.001557547, 0.001556254, 
    0.001560923, 0.00151312, 0.001515993, 0.001515741, 0.001518747, 
    0.001520969, 0.001525786, 0.001533505, 0.001530603, 0.00153593, 
    0.001536999, 0.001528906, 0.001533876, 0.001517916, 0.001520496, 
    0.00151896, 0.001513346, 0.001531271, 0.001522076, 0.00153905, 
    0.001534073, 0.001548589, 0.001541373, 0.001555542, 0.001561591, 
    0.001567283, 0.001573928, 0.001517561, 0.001515609, 0.001519104, 
    0.001523937, 0.00152842, 0.001534377, 0.001534986, 0.001536101, 
    0.00153899, 0.001541418, 0.001536454, 0.001542027, 0.001521093, 
    0.001532069, 0.001514871, 0.001520052, 0.001523652, 0.001522074, 
    0.001530271, 0.001532202, 0.001540045, 0.001535992, 0.001560098, 
    0.00154944, 0.001578985, 0.001570738, 0.001514927, 0.001517555, 
    0.001526693, 0.001522346, 0.001534775, 0.001537831, 0.001540315, 
    0.00154349, 0.001543833, 0.001545713, 0.001542632, 0.001545591, 
    0.001534389, 0.001539397, 0.00152565, 0.001528997, 0.001527458, 
    0.001525768, 0.001530982, 0.001536532, 0.001536651, 0.00153843, 
    0.001543439, 0.001534825, 0.001561471, 0.001545023, 0.001520419, 
    0.001525476, 0.001526199, 0.00152424, 0.001537525, 0.001532713, 
    0.001545667, 0.001542168, 0.001547901, 0.001545052, 0.001544633, 
    0.001540974, 0.001538694, 0.001532934, 0.001528244, 0.001524524, 
    0.001525389, 0.001529475, 0.001536871, 0.001543863, 0.001542332, 
    0.001547465, 0.001533874, 0.001539575, 0.001537372, 0.001543116, 
    0.001530526, 0.001541245, 0.001527784, 0.001528965, 0.001532618, 
    0.001539961, 0.001541586, 0.001543319, 0.00154225, 0.001537059, 
    0.001536209, 0.001532529, 0.001531512, 0.001528708, 0.001526385, 
    0.001528507, 0.001530735, 0.001537062, 0.001542759, 0.001548967, 
    0.001550486, 0.001557731, 0.001551832, 0.001561563, 0.001553289, 
    0.001567607, 0.001541868, 0.001553047, 0.001532784, 0.001534969, 
    0.00153892, 0.001547976, 0.001543089, 0.001548804, 0.001536175, 
    0.001529616, 0.001527919, 0.00152475, 0.001527991, 0.001527728, 
    0.001530828, 0.001529832, 0.001537272, 0.001533276, 0.001544622, 
    0.001548759, 0.001560433, 0.001567582, 0.001574854, 0.001578063, 
    0.001579039, 0.001579447,
  0.001428957, 0.001435722, 0.001434407, 0.001439863, 0.001436836, 
    0.001440409, 0.001430328, 0.00143599, 0.001432376, 0.001429566, 
    0.001450447, 0.001440106, 0.001461187, 0.001454594, 0.001471154, 
    0.001460161, 0.00147337, 0.001470837, 0.001478461, 0.001476277, 
    0.001486026, 0.001479469, 0.001491079, 0.00148446, 0.001485496, 
    0.001479253, 0.001442187, 0.00144916, 0.001441774, 0.001442769, 
    0.001442323, 0.001436899, 0.001434165, 0.00142844, 0.001429479, 
    0.001433684, 0.001443216, 0.001439981, 0.001448134, 0.00144795, 
    0.001457024, 0.001452933, 0.001468181, 0.001463848, 0.001476368, 
    0.00147322, 0.00147622, 0.001475311, 0.001476232, 0.001471615, 
    0.001473593, 0.00146953, 0.001453699, 0.001458352, 0.001444472, 
    0.001436123, 0.001430577, 0.001426641, 0.001427197, 0.001428258, 
    0.001433709, 0.001438834, 0.001442738, 0.00144535, 0.001447923, 
    0.00145571, 0.001459832, 0.001469057, 0.001467393, 0.001470213, 
    0.001472907, 0.001477429, 0.001476685, 0.001478677, 0.001470139, 
    0.001475814, 0.001466444, 0.001469007, 0.001448622, 0.001440854, 
    0.001437551, 0.00143466, 0.001427625, 0.001432483, 0.001430568, 
    0.001435124, 0.001438019, 0.001436587, 0.001445421, 0.001441987, 
    0.001460076, 0.001452286, 0.001472593, 0.001467734, 0.001473757, 
    0.001470684, 0.001475949, 0.001471211, 0.001479419, 0.001481206, 
    0.001479984, 0.001484675, 0.001470948, 0.00147622, 0.001436547, 
    0.00143678, 0.001437868, 0.001433086, 0.001432794, 0.001428411, 
    0.001432311, 0.001433971, 0.001438186, 0.001440679, 0.001443049, 
    0.001448258, 0.001454075, 0.001462208, 0.001468049, 0.001471964, 
    0.001469564, 0.001471683, 0.001469314, 0.001468203, 0.001480536, 
    0.001473612, 0.001484001, 0.001483426, 0.001478725, 0.001483491, 
    0.001436944, 0.001435601, 0.001430935, 0.001434586, 0.001427934, 
    0.001431658, 0.001433799, 0.001442059, 0.001443873, 0.001445556, 
    0.001448878, 0.001453142, 0.001460621, 0.001467126, 0.001473064, 
    0.001472629, 0.001472782, 0.001474108, 0.001470823, 0.001474647, 
    0.001475289, 0.001473611, 0.001483349, 0.001480567, 0.001483414, 
    0.001481603, 0.001436037, 0.001438298, 0.001437077, 0.001439374, 
    0.001437755, 0.001444951, 0.001447108, 0.001457199, 0.001453058, 
    0.001459649, 0.001453728, 0.001454777, 0.001459864, 0.001454048, 
    0.001466767, 0.001458144, 0.00147416, 0.00146555, 0.001474699, 
    0.001473038, 0.001475788, 0.001478251, 0.001481349, 0.001487065, 
    0.001485741, 0.001490521, 0.001441668, 0.0014446, 0.001444342, 
    0.00144741, 0.001449679, 0.001454596, 0.00146248, 0.001459516, 
    0.001464958, 0.001466051, 0.001457782, 0.001462859, 0.001446562, 
    0.001449195, 0.001447628, 0.001441899, 0.001460199, 0.001450809, 
    0.001468146, 0.001463061, 0.0014779, 0.001470521, 0.001485013, 
    0.001491206, 0.001497033, 0.001503842, 0.0014462, 0.001444208, 
    0.001447775, 0.001452709, 0.001457286, 0.001463371, 0.001463993, 
    0.001465133, 0.001468085, 0.001470567, 0.001465493, 0.001471189, 
    0.001449806, 0.001461014, 0.001443455, 0.001448743, 0.001452418, 
    0.001450806, 0.001459177, 0.001461149, 0.001469164, 0.001465021, 
    0.001489677, 0.001478771, 0.001509025, 0.001500573, 0.001443512, 
    0.001446193, 0.001455523, 0.001451084, 0.001463777, 0.0014669, 
    0.001469439, 0.001472685, 0.001473035, 0.001474958, 0.001471807, 
    0.001474833, 0.001463384, 0.001468501, 0.001454457, 0.001457875, 
    0.001456303, 0.001454578, 0.001459902, 0.001465573, 0.001465694, 
    0.001467513, 0.001472636, 0.001463828, 0.001491084, 0.001474254, 
    0.001449117, 0.00145428, 0.001455017, 0.001453017, 0.001466587, 
    0.001461671, 0.001474911, 0.001471333, 0.001477195, 0.001474282, 
    0.001473854, 0.001470112, 0.001467783, 0.001461896, 0.001457106, 
    0.001453308, 0.001454191, 0.001458364, 0.00146592, 0.001473067, 
    0.001471501, 0.00147675, 0.001462857, 0.001468683, 0.001466431, 
    0.001472302, 0.001459437, 0.001470392, 0.001456636, 0.001457842, 
    0.001461574, 0.001469078, 0.001470738, 0.001472511, 0.001471417, 
    0.001466112, 0.001465243, 0.001461483, 0.001460445, 0.001457579, 
    0.001455207, 0.001457375, 0.001459651, 0.001466114, 0.001471938, 
    0.001478286, 0.001479839, 0.001487254, 0.001481218, 0.001491178, 
    0.00148271, 0.001497367, 0.001471027, 0.001482461, 0.001461743, 
    0.001463976, 0.001468014, 0.001477273, 0.001472275, 0.00147812, 
    0.001465209, 0.001458508, 0.001456774, 0.001453539, 0.001456848, 
    0.001456579, 0.001459745, 0.001458728, 0.001466329, 0.001462246, 
    0.001473843, 0.001478074, 0.00149002, 0.00149734, 0.001504791, 
    0.001508079, 0.00150908, 0.001509498,
  0.001343041, 0.00134928, 0.001348067, 0.001353102, 0.001350309, 
    0.001353606, 0.001344305, 0.001349528, 0.001346194, 0.001343602, 
    0.001362882, 0.001353327, 0.001372816, 0.001366715, 0.001382048, 
    0.001371866, 0.001384103, 0.001381754, 0.001388824, 0.001386798, 
    0.001395847, 0.001389759, 0.001400542, 0.001394393, 0.001395355, 
    0.001389558, 0.001355249, 0.001361692, 0.001354867, 0.001355786, 
    0.001355373, 0.001350366, 0.001347844, 0.001342564, 0.001343522, 
    0.001347401, 0.001356199, 0.001353211, 0.001360742, 0.001360572, 
    0.001368963, 0.001365178, 0.001379293, 0.001375279, 0.001386883, 
    0.001383963, 0.001386745, 0.001385902, 0.001386756, 0.001382475, 
    0.001384309, 0.001380543, 0.001365887, 0.001370192, 0.001357359, 
    0.001349651, 0.001344534, 0.001340905, 0.001341418, 0.001342396, 
    0.001347423, 0.001352152, 0.001355757, 0.00135817, 0.001360547, 
    0.001367748, 0.001371561, 0.001380105, 0.001378562, 0.001381176, 
    0.001383673, 0.001387867, 0.001387176, 0.001389025, 0.001381106, 
    0.001386368, 0.001377684, 0.001380058, 0.001361195, 0.001354017, 
    0.001350968, 0.0013483, 0.001341813, 0.001346292, 0.001344526, 
    0.001348728, 0.0013514, 0.001350078, 0.001358235, 0.001355063, 
    0.001371787, 0.00136458, 0.001383381, 0.001378879, 0.001384461, 
    0.001381612, 0.001386494, 0.0013821, 0.001389713, 0.001391371, 
    0.001390238, 0.001394592, 0.001381857, 0.001386745, 0.001350041, 
    0.001350257, 0.001351261, 0.001346849, 0.001346579, 0.001342537, 
    0.001346133, 0.001347665, 0.001351554, 0.001353856, 0.001356044, 
    0.001360857, 0.001366235, 0.001373761, 0.001379171, 0.001382799, 
    0.001380574, 0.001382538, 0.001380342, 0.001379313, 0.00139075, 
    0.001384326, 0.001393966, 0.001393432, 0.001389069, 0.001393492, 
    0.001350408, 0.001349168, 0.001344865, 0.001348232, 0.001342097, 
    0.001345531, 0.001347506, 0.00135513, 0.001356806, 0.00135836, 
    0.00136143, 0.001365372, 0.001372291, 0.001378315, 0.001383818, 
    0.001383414, 0.001383557, 0.001384786, 0.001381741, 0.001385286, 
    0.001385882, 0.001384325, 0.001393361, 0.001390778, 0.001393421, 
    0.001391739, 0.001349571, 0.001351658, 0.00135053, 0.001352651, 
    0.001351157, 0.001357801, 0.001359794, 0.001369125, 0.001365294, 
    0.001371392, 0.001365914, 0.001366884, 0.001371591, 0.001366209, 
    0.001377983, 0.00137, 0.001384834, 0.001376856, 0.001385334, 0.001383794, 
    0.001386344, 0.001388629, 0.001391504, 0.001396811, 0.001395582, 
    0.001400022, 0.001354769, 0.001357477, 0.001357238, 0.001360073, 
    0.00136217, 0.001366716, 0.001374012, 0.001371268, 0.001376307, 
    0.001377319, 0.001369664, 0.001374363, 0.00135929, 0.001361724, 
    0.001360274, 0.001354983, 0.001371901, 0.001363215, 0.00137926, 
    0.00137455, 0.001388303, 0.001381461, 0.001394905, 0.00140066, 
    0.001406078, 0.001412415, 0.001358955, 0.001357115, 0.00136041, 
    0.001364972, 0.001369205, 0.001374837, 0.001375413, 0.001376469, 
    0.001379204, 0.001381503, 0.001376803, 0.00138208, 0.001362289, 
    0.001372655, 0.001356419, 0.001361305, 0.001364702, 0.001363212, 
    0.001370954, 0.00137278, 0.001380203, 0.001376365, 0.001399239, 
    0.001389112, 0.001417242, 0.001409372, 0.001356472, 0.001358949, 
    0.001367574, 0.001363469, 0.001375213, 0.001378106, 0.001380459, 
    0.001383467, 0.001383792, 0.001385574, 0.001382653, 0.001385459, 
    0.001374849, 0.001379589, 0.001366588, 0.00136975, 0.001368295, 
    0.001366699, 0.001371626, 0.001376877, 0.001376989, 0.001378673, 
    0.001383423, 0.001375261, 0.001400548, 0.001384923, 0.00136165, 
    0.001366425, 0.001367106, 0.001365256, 0.001377816, 0.001373263, 
    0.001385531, 0.001382214, 0.001387649, 0.001384948, 0.001384551, 
    0.001381082, 0.001378924, 0.001373472, 0.001369039, 0.001365525, 
    0.001366342, 0.001370202, 0.001377198, 0.001383821, 0.00138237, 
    0.001387236, 0.001374361, 0.001379758, 0.001377672, 0.001383112, 
    0.001371195, 0.001381343, 0.001368603, 0.001369719, 0.001373173, 
    0.001380124, 0.001381662, 0.001383306, 0.001382291, 0.001377376, 
    0.001376571, 0.001373089, 0.001372128, 0.001369476, 0.001367282, 
    0.001369287, 0.001371393, 0.001377378, 0.001382774, 0.001388662, 
    0.001390103, 0.001396988, 0.001391383, 0.001400635, 0.00139277, 
    0.001406389, 0.001381931, 0.001392537, 0.00137333, 0.001375397, 
    0.001379138, 0.001387722, 0.001383087, 0.001388508, 0.001376539, 
    0.001370336, 0.001368731, 0.001365738, 0.001368799, 0.00136855, 
    0.00137148, 0.001370539, 0.001377576, 0.001373795, 0.001384541, 
    0.001388465, 0.001399557, 0.001406364, 0.001413297, 0.00141636, 
    0.001417293, 0.001417683,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.212406e-06, 1.222874e-06, 1.220835e-06, 1.229305e-06, 1.224603e-06, 
    1.230154e-06, 1.214524e-06, 1.22329e-06, 1.21769e-06, 1.213346e-06, 
    1.245827e-06, 1.229683e-06, 1.262715e-06, 1.252333e-06, 1.278499e-06, 
    1.261096e-06, 1.282023e-06, 1.277995e-06, 1.290139e-06, 1.286654e-06, 
    1.30225e-06, 1.291749e-06, 1.310374e-06, 1.299738e-06, 1.301398e-06, 
    1.291402e-06, 1.232924e-06, 1.243812e-06, 1.23228e-06, 1.233829e-06, 
    1.233134e-06, 1.224699e-06, 1.22046e-06, 1.211607e-06, 1.213212e-06, 
    1.219715e-06, 1.234525e-06, 1.229487e-06, 1.242205e-06, 1.241917e-06, 
    1.256153e-06, 1.249724e-06, 1.27378e-06, 1.266918e-06, 1.286799e-06, 
    1.281784e-06, 1.286563e-06, 1.285112e-06, 1.286581e-06, 1.27923e-06, 
    1.282377e-06, 1.275918e-06, 1.250928e-06, 1.258246e-06, 1.236485e-06, 
    1.223495e-06, 1.214907e-06, 1.208833e-06, 1.20969e-06, 1.211326e-06, 
    1.219753e-06, 1.227704e-06, 1.233781e-06, 1.237854e-06, 1.241875e-06, 
    1.254086e-06, 1.260576e-06, 1.275169e-06, 1.272529e-06, 1.277003e-06, 
    1.281285e-06, 1.288491e-06, 1.287303e-06, 1.290483e-06, 1.276884e-06, 
    1.285913e-06, 1.271026e-06, 1.275088e-06, 1.242969e-06, 1.230846e-06, 
    1.225711e-06, 1.221226e-06, 1.21035e-06, 1.217855e-06, 1.214893e-06, 
    1.221945e-06, 1.226437e-06, 1.224214e-06, 1.237966e-06, 1.23261e-06, 
    1.260961e-06, 1.248708e-06, 1.280785e-06, 1.273071e-06, 1.282638e-06, 
    1.277751e-06, 1.28613e-06, 1.278588e-06, 1.291667e-06, 1.294524e-06, 
    1.292571e-06, 1.300081e-06, 1.278169e-06, 1.286561e-06, 1.224153e-06, 
    1.224515e-06, 1.226204e-06, 1.218788e-06, 1.218336e-06, 1.211562e-06, 
    1.217588e-06, 1.220159e-06, 1.226697e-06, 1.230573e-06, 1.234264e-06, 
    1.242399e-06, 1.251516e-06, 1.264325e-06, 1.27357e-06, 1.279786e-06, 
    1.275972e-06, 1.279339e-06, 1.275575e-06, 1.273813e-06, 1.293453e-06, 
    1.282405e-06, 1.298999e-06, 1.298078e-06, 1.290557e-06, 1.298182e-06, 
    1.224769e-06, 1.222684e-06, 1.215461e-06, 1.221112e-06, 1.210826e-06, 
    1.216578e-06, 1.219891e-06, 1.232721e-06, 1.235549e-06, 1.238175e-06, 
    1.243369e-06, 1.250051e-06, 1.261819e-06, 1.272105e-06, 1.281534e-06, 
    1.280842e-06, 1.281085e-06, 1.283196e-06, 1.27797e-06, 1.284054e-06, 
    1.285076e-06, 1.282404e-06, 1.297955e-06, 1.293502e-06, 1.298058e-06, 
    1.295158e-06, 1.223362e-06, 1.226871e-06, 1.224974e-06, 1.228543e-06, 
    1.226028e-06, 1.23723e-06, 1.240599e-06, 1.256429e-06, 1.24992e-06, 
    1.260287e-06, 1.250971e-06, 1.252619e-06, 1.260625e-06, 1.251473e-06, 
    1.271536e-06, 1.257915e-06, 1.283277e-06, 1.269609e-06, 1.284136e-06, 
    1.281492e-06, 1.285871e-06, 1.2898e-06, 1.294752e-06, 1.303915e-06, 
    1.30179e-06, 1.309472e-06, 1.232113e-06, 1.236683e-06, 1.236281e-06, 
    1.241072e-06, 1.244622e-06, 1.252334e-06, 1.264755e-06, 1.260077e-06, 
    1.268673e-06, 1.270402e-06, 1.257345e-06, 1.265353e-06, 1.239746e-06, 
    1.243864e-06, 1.241411e-06, 1.232471e-06, 1.261152e-06, 1.24639e-06, 
    1.273721e-06, 1.265671e-06, 1.289239e-06, 1.277489e-06, 1.300621e-06, 
    1.310574e-06, 1.31998e-06, 1.331014e-06, 1.239181e-06, 1.236072e-06, 
    1.241642e-06, 1.249371e-06, 1.256565e-06, 1.266162e-06, 1.267147e-06, 
    1.268949e-06, 1.273626e-06, 1.277564e-06, 1.269519e-06, 1.278552e-06, 
    1.244819e-06, 1.262438e-06, 1.234895e-06, 1.243155e-06, 1.248913e-06, 
    1.246386e-06, 1.259541e-06, 1.262652e-06, 1.275335e-06, 1.26877e-06, 
    1.308113e-06, 1.290629e-06, 1.339449e-06, 1.325711e-06, 1.234986e-06, 
    1.23917e-06, 1.253791e-06, 1.246823e-06, 1.266804e-06, 1.271748e-06, 
    1.275774e-06, 1.280931e-06, 1.281488e-06, 1.284549e-06, 1.279535e-06, 
    1.28435e-06, 1.266181e-06, 1.274284e-06, 1.252114e-06, 1.257491e-06, 
    1.255016e-06, 1.252303e-06, 1.260684e-06, 1.269644e-06, 1.269836e-06, 
    1.272716e-06, 1.280849e-06, 1.266883e-06, 1.310377e-06, 1.283425e-06, 
    1.243742e-06, 1.251837e-06, 1.252996e-06, 1.249855e-06, 1.271251e-06, 
    1.263477e-06, 1.284474e-06, 1.278781e-06, 1.288115e-06, 1.283473e-06, 
    1.28279e-06, 1.276842e-06, 1.273145e-06, 1.263831e-06, 1.25628e-06, 
    1.250309e-06, 1.251696e-06, 1.258259e-06, 1.270192e-06, 1.281536e-06, 
    1.279047e-06, 1.287403e-06, 1.265347e-06, 1.274571e-06, 1.271001e-06, 
    1.280319e-06, 1.259952e-06, 1.277286e-06, 1.255541e-06, 1.257439e-06, 
    1.263322e-06, 1.2752e-06, 1.277836e-06, 1.280653e-06, 1.278914e-06, 
    1.270497e-06, 1.269121e-06, 1.263178e-06, 1.26154e-06, 1.257024e-06, 
    1.253292e-06, 1.256702e-06, 1.260287e-06, 1.2705e-06, 1.27974e-06, 
    1.289854e-06, 1.292336e-06, 1.304217e-06, 1.29454e-06, 1.310528e-06, 
    1.296927e-06, 1.320517e-06, 1.278295e-06, 1.296532e-06, 1.263591e-06, 
    1.267118e-06, 1.273511e-06, 1.288239e-06, 1.280277e-06, 1.289591e-06, 
    1.269067e-06, 1.258486e-06, 1.255756e-06, 1.250671e-06, 1.255872e-06, 
    1.255449e-06, 1.260436e-06, 1.258832e-06, 1.270839e-06, 1.264382e-06, 
    1.282771e-06, 1.289516e-06, 1.308664e-06, 1.320475e-06, 1.332555e-06, 
    1.337906e-06, 1.339537e-06, 1.340219e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.529265e-06, 7.563329e-06, 7.55669e-06, 7.584184e-06, 7.568925e-06, 
    7.586915e-06, 7.536134e-06, 7.56462e-06, 7.546424e-06, 7.532271e-06, 
    7.637537e-06, 7.585349e-06, 7.691932e-06, 7.658536e-06, 7.742495e-06, 
    7.686703e-06, 7.753753e-06, 7.740879e-06, 7.779649e-06, 7.768524e-06, 
    7.818129e-06, 7.784757e-06, 7.843899e-06, 7.810151e-06, 7.81541e-06, 
    7.783614e-06, 7.595916e-06, 7.631089e-06, 7.593813e-06, 7.598828e-06, 
    7.596572e-06, 7.569199e-06, 7.555409e-06, 7.526601e-06, 7.531818e-06, 
    7.552978e-06, 7.601024e-06, 7.584699e-06, 7.625855e-06, 7.624927e-06, 
    7.670808e-06, 7.650105e-06, 7.72738e-06, 7.705381e-06, 7.768978e-06, 
    7.752953e-06, 7.768206e-06, 7.763569e-06, 7.768243e-06, 7.744767e-06, 
    7.754804e-06, 7.734161e-06, 7.654074e-06, 7.677619e-06, 7.607413e-06, 
    7.565262e-06, 7.537345e-06, 7.517553e-06, 7.520332e-06, 7.525664e-06, 
    7.553085e-06, 7.578908e-06, 7.598606e-06, 7.611779e-06, 7.624769e-06, 
    7.664122e-06, 7.685003e-06, 7.731802e-06, 7.723358e-06, 7.737656e-06, 
    7.751352e-06, 7.774336e-06, 7.770549e-06, 7.780669e-06, 7.737246e-06, 
    7.766086e-06, 7.718477e-06, 7.731484e-06, 7.628328e-06, 7.589138e-06, 
    7.572452e-06, 7.55789e-06, 7.522477e-06, 7.546918e-06, 7.537269e-06, 
    7.560206e-06, 7.574788e-06, 7.567563e-06, 7.612131e-06, 7.594778e-06, 
    7.686228e-06, 7.646793e-06, 7.749764e-06, 7.725073e-06, 7.755661e-06, 
    7.740048e-06, 7.766787e-06, 7.742707e-06, 7.78443e-06, 7.793522e-06, 
    7.78729e-06, 7.811191e-06, 7.741321e-06, 7.768119e-06, 7.567406e-06, 
    7.568583e-06, 7.574058e-06, 7.549941e-06, 7.548467e-06, 7.526406e-06, 
    7.546019e-06, 7.554377e-06, 7.575617e-06, 7.588172e-06, 7.600118e-06, 
    7.626431e-06, 7.655829e-06, 7.697016e-06, 7.726662e-06, 7.746541e-06, 
    7.734343e-06, 7.745096e-06, 7.733055e-06, 7.727405e-06, 7.790088e-06, 
    7.754863e-06, 7.807728e-06, 7.804803e-06, 7.780844e-06, 7.805109e-06, 
    7.569394e-06, 7.562614e-06, 7.53911e-06, 7.557487e-06, 7.52399e-06, 
    7.542723e-06, 7.553484e-06, 7.595116e-06, 7.604279e-06, 7.612772e-06, 
    7.629554e-06, 7.651101e-06, 7.688962e-06, 7.72195e-06, 7.752119e-06, 
    7.749895e-06, 7.750669e-06, 7.757395e-06, 7.740695e-06, 7.760122e-06, 
    7.763369e-06, 7.754844e-06, 7.804387e-06, 7.79022e-06, 7.804708e-06, 
    7.795471e-06, 7.564806e-06, 7.576185e-06, 7.570017e-06, 7.581596e-06, 
    7.573417e-06, 7.609714e-06, 7.620596e-06, 7.671633e-06, 7.650673e-06, 
    7.684041e-06, 7.654049e-06, 7.659356e-06, 7.685077e-06, 7.65565e-06, 
    7.720093e-06, 7.676347e-06, 7.757648e-06, 7.713875e-06, 7.760375e-06, 
    7.751921e-06, 7.765894e-06, 7.77842e-06, 7.794177e-06, 7.823293e-06, 
    7.816533e-06, 7.840911e-06, 7.593176e-06, 7.607953e-06, 7.606658e-06, 
    7.622139e-06, 7.633592e-06, 7.658471e-06, 7.6984e-06, 7.683364e-06, 
    7.710952e-06, 7.716494e-06, 7.674556e-06, 7.700278e-06, 7.617781e-06, 
    7.631065e-06, 7.623152e-06, 7.594211e-06, 7.686742e-06, 7.63919e-06, 
    7.727052e-06, 7.701236e-06, 7.776608e-06, 7.739081e-06, 7.812814e-06, 
    7.844376e-06, 7.874155e-06, 7.908933e-06, 7.616031e-06, 7.605964e-06, 
    7.62397e-06, 7.6489e-06, 7.672066e-06, 7.702905e-06, 7.706059e-06, 
    7.711824e-06, 7.726802e-06, 7.739407e-06, 7.713621e-06, 7.742546e-06, 
    7.634118e-06, 7.690875e-06, 7.602046e-06, 7.628745e-06, 7.647321e-06, 
    7.639175e-06, 7.681545e-06, 7.691527e-06, 7.732169e-06, 7.711154e-06, 
    7.836549e-06, 7.78099e-06, 7.935474e-06, 7.892205e-06, 7.60244e-06, 
    7.615968e-06, 7.663125e-06, 7.640675e-06, 7.704947e-06, 7.720795e-06, 
    7.733675e-06, 7.750156e-06, 7.751926e-06, 7.761699e-06, 7.74567e-06, 
    7.761054e-06, 7.702883e-06, 7.728858e-06, 7.657653e-06, 7.674943e-06, 
    7.666982e-06, 7.658236e-06, 7.685189e-06, 7.713932e-06, 7.714554e-06, 
    7.723761e-06, 7.749724e-06, 7.705058e-06, 7.843664e-06, 7.757932e-06, 
    7.630731e-06, 7.656812e-06, 7.660552e-06, 7.650438e-06, 7.719182e-06, 
    7.694244e-06, 7.761462e-06, 7.743267e-06, 7.77306e-06, 7.758246e-06, 
    7.756048e-06, 7.737039e-06, 7.725187e-06, 7.695319e-06, 7.671029e-06, 
    7.65181e-06, 7.656262e-06, 7.677382e-06, 7.715672e-06, 7.751979e-06, 
    7.744008e-06, 7.770691e-06, 7.700112e-06, 7.729672e-06, 7.71822e-06, 
    7.748049e-06, 7.682927e-06, 7.738465e-06, 7.668737e-06, 7.674833e-06, 
    7.693726e-06, 7.73179e-06, 7.740226e-06, 7.749227e-06, 7.74366e-06, 
    7.716709e-06, 7.712293e-06, 7.693217e-06, 7.687936e-06, 7.67343e-06, 
    7.6614e-06, 7.672373e-06, 7.683878e-06, 7.716663e-06, 7.746223e-06, 
    7.778494e-06, 7.786404e-06, 7.824129e-06, 7.793376e-06, 7.844098e-06, 
    7.800917e-06, 7.875709e-06, 7.741689e-06, 7.799853e-06, 7.694594e-06, 
    7.705904e-06, 7.726373e-06, 7.773416e-06, 7.748009e-06, 7.777722e-06, 
    7.712117e-06, 7.678116e-06, 7.669341e-06, 7.652964e-06, 7.6697e-06, 
    7.668339e-06, 7.68437e-06, 7.679202e-06, 7.717729e-06, 7.697024e-06, 
    7.75588e-06, 7.777395e-06, 7.838255e-06, 7.875613e-06, 7.913733e-06, 
    7.930556e-06, 7.935681e-06, 7.937815e-06,
  3.965582e-06, 3.995709e-06, 3.989847e-06, 4.014192e-06, 4.000683e-06, 
    4.016632e-06, 3.971687e-06, 3.996904e-06, 3.980801e-06, 3.968295e-06, 
    4.061586e-06, 4.01528e-06, 4.109927e-06, 4.080236e-06, 4.154983e-06, 
    4.105297e-06, 4.16503e-06, 4.153555e-06, 4.188147e-06, 4.178226e-06, 
    4.222569e-06, 4.192728e-06, 4.245635e-06, 4.21544e-06, 4.220155e-06, 
    4.191744e-06, 4.02459e-06, 4.055808e-06, 4.022742e-06, 4.027188e-06, 
    4.025194e-06, 4.00096e-06, 3.988763e-06, 3.963288e-06, 3.96791e-06, 
    3.986625e-06, 4.029187e-06, 4.014726e-06, 4.051225e-06, 4.0504e-06, 
    4.091172e-06, 4.07277e-06, 4.141531e-06, 4.121946e-06, 4.17864e-06, 
    4.164354e-06, 4.177968e-06, 4.173839e-06, 4.178021e-06, 4.157077e-06, 
    4.166046e-06, 4.147636e-06, 4.076212e-06, 4.097153e-06, 4.034813e-06, 
    3.997489e-06, 3.97279e-06, 3.955292e-06, 3.957764e-06, 3.962477e-06, 
    3.986735e-06, 4.009601e-06, 4.027057e-06, 4.038748e-06, 4.050281e-06, 
    4.085246e-06, 4.103815e-06, 4.145492e-06, 4.137965e-06, 4.150724e-06, 
    4.162935e-06, 4.183456e-06, 4.180077e-06, 4.189126e-06, 4.150392e-06, 
    4.176118e-06, 4.133679e-06, 4.14527e-06, 4.053393e-06, 4.018626e-06, 
    4.003861e-06, 3.990973e-06, 3.959665e-06, 3.981274e-06, 3.97275e-06, 
    3.993047e-06, 4.005961e-06, 3.999573e-06, 4.039068e-06, 4.023695e-06, 
    4.104917e-06, 4.069857e-06, 4.16151e-06, 4.139511e-06, 4.16679e-06, 
    4.152863e-06, 4.176734e-06, 4.155248e-06, 4.192498e-06, 4.200622e-06, 
    4.195069e-06, 4.216423e-06, 4.154057e-06, 4.177965e-06, 3.999393e-06, 
    4.000434e-06, 4.00529e-06, 3.983961e-06, 3.982659e-06, 3.96316e-06, 
    3.98051e-06, 3.987906e-06, 4.006712e-06, 4.017847e-06, 4.028444e-06, 
    4.051782e-06, 4.0779e-06, 4.114536e-06, 4.140935e-06, 4.158664e-06, 
    4.147791e-06, 4.15739e-06, 4.146659e-06, 4.141634e-06, 4.197575e-06, 
    4.166128e-06, 4.21335e-06, 4.210733e-06, 4.18934e-06, 4.211027e-06, 
    4.001166e-06, 3.995173e-06, 3.974385e-06, 3.99065e-06, 3.961039e-06, 
    3.9776e-06, 3.987133e-06, 4.024011e-06, 4.032136e-06, 4.039668e-06, 
    4.054565e-06, 4.073711e-06, 4.107376e-06, 4.136756e-06, 4.163647e-06, 
    4.161674e-06, 4.162368e-06, 4.168381e-06, 4.15349e-06, 4.170828e-06, 
    4.173738e-06, 4.166127e-06, 4.210382e-06, 4.197721e-06, 4.210677e-06, 
    4.202433e-06, 3.997121e-06, 4.00721e-06, 4.001757e-06, 4.012012e-06, 
    4.004784e-06, 4.036953e-06, 4.046617e-06, 4.091956e-06, 4.073332e-06, 
    4.102995e-06, 4.076344e-06, 4.08106e-06, 4.103953e-06, 4.077784e-06, 
    4.135129e-06, 4.096209e-06, 4.168615e-06, 4.129623e-06, 4.171062e-06, 
    4.16353e-06, 4.176006e-06, 4.187189e-06, 4.201278e-06, 4.227311e-06, 
    4.221279e-06, 4.243087e-06, 4.022269e-06, 4.035385e-06, 4.034234e-06, 
    4.047979e-06, 4.058154e-06, 4.080247e-06, 4.115768e-06, 4.102399e-06, 
    4.12696e-06, 4.131896e-06, 4.094588e-06, 4.117475e-06, 4.044176e-06, 
    4.05598e-06, 4.048954e-06, 4.023301e-06, 4.105471e-06, 4.063221e-06, 
    4.141371e-06, 4.118389e-06, 4.185593e-06, 4.152116e-06, 4.217958e-06, 
    4.246207e-06, 4.272878e-06, 4.304096e-06, 4.042555e-06, 4.033635e-06, 
    4.049616e-06, 4.071757e-06, 4.092354e-06, 4.119789e-06, 4.122602e-06, 
    4.127749e-06, 4.141098e-06, 4.152332e-06, 4.129372e-06, 4.15515e-06, 
    4.05871e-06, 4.109148e-06, 4.03026e-06, 4.053949e-06, 4.070453e-06, 
    4.063214e-06, 4.100873e-06, 4.109766e-06, 4.145974e-06, 4.127245e-06, 
    4.239223e-06, 4.189546e-06, 4.327937e-06, 4.289097e-06, 4.030519e-06, 
    4.042527e-06, 4.084414e-06, 4.064465e-06, 4.121625e-06, 4.135738e-06, 
    4.147228e-06, 4.161926e-06, 4.163517e-06, 4.172236e-06, 4.157951e-06, 
    4.171673e-06, 4.119847e-06, 4.142978e-06, 4.079624e-06, 4.095008e-06, 
    4.087929e-06, 4.080167e-06, 4.104141e-06, 4.129732e-06, 4.130287e-06, 
    4.138505e-06, 4.161679e-06, 4.121857e-06, 4.245636e-06, 4.169022e-06, 
    4.055635e-06, 4.078818e-06, 4.082143e-06, 4.073152e-06, 4.134322e-06, 
    4.112118e-06, 4.172024e-06, 4.155804e-06, 4.182395e-06, 4.169173e-06, 
    4.167228e-06, 4.150274e-06, 4.139729e-06, 4.113133e-06, 4.091543e-06, 
    4.074457e-06, 4.078428e-06, 4.097205e-06, 4.131301e-06, 4.163658e-06, 
    4.156561e-06, 4.180372e-06, 4.11747e-06, 4.143799e-06, 4.133613e-06, 
    4.160194e-06, 4.102042e-06, 4.151519e-06, 4.089428e-06, 4.094859e-06, 
    4.111678e-06, 4.145582e-06, 4.153108e-06, 4.161136e-06, 4.156183e-06, 
    4.13217e-06, 4.128244e-06, 4.111271e-06, 4.106585e-06, 4.093677e-06, 
    4.082999e-06, 4.092753e-06, 4.103004e-06, 4.132183e-06, 4.158539e-06, 
    4.187347e-06, 4.194411e-06, 4.228163e-06, 4.200669e-06, 4.246062e-06, 
    4.207442e-06, 4.274385e-06, 4.154404e-06, 4.206324e-06, 4.112446e-06, 
    4.122524e-06, 4.140767e-06, 4.182738e-06, 4.160069e-06, 4.186589e-06, 
    4.12809e-06, 4.09785e-06, 4.090049e-06, 4.075494e-06, 4.090382e-06, 
    4.089171e-06, 4.103435e-06, 4.098849e-06, 4.133153e-06, 4.114714e-06, 
    4.167177e-06, 4.186381e-06, 4.240797e-06, 4.274276e-06, 4.308466e-06, 
    4.323586e-06, 4.328193e-06, 4.330118e-06,
  3.780337e-06, 3.813905e-06, 3.80737e-06, 3.834516e-06, 3.819449e-06, 
    3.837237e-06, 3.787134e-06, 3.815238e-06, 3.797288e-06, 3.783356e-06, 
    3.887426e-06, 3.835729e-06, 3.941455e-06, 3.908253e-06, 3.99189e-06, 
    3.936279e-06, 4.003145e-06, 3.990286e-06, 4.029051e-06, 4.01793e-06, 
    4.067675e-06, 4.034189e-06, 4.09357e-06, 4.05967e-06, 4.064964e-06, 
    4.033085e-06, 3.846113e-06, 3.880972e-06, 3.844051e-06, 3.849013e-06, 
    3.846787e-06, 3.819758e-06, 3.806166e-06, 3.777779e-06, 3.782927e-06, 
    3.803781e-06, 3.851245e-06, 3.835107e-06, 3.875841e-06, 3.874919e-06, 
    3.920477e-06, 3.899908e-06, 3.976821e-06, 3.954897e-06, 4.018394e-06, 
    4.002384e-06, 4.017641e-06, 4.013013e-06, 4.017701e-06, 3.994232e-06, 
    4.00428e-06, 3.983656e-06, 3.903756e-06, 3.927165e-06, 3.857521e-06, 
    3.815895e-06, 3.788364e-06, 3.768876e-06, 3.771629e-06, 3.776877e-06, 
    3.803903e-06, 3.829391e-06, 3.848863e-06, 3.861911e-06, 3.874787e-06, 
    3.913861e-06, 3.934618e-06, 3.981258e-06, 3.972828e-06, 3.987117e-06, 
    4.000794e-06, 4.023794e-06, 4.020005e-06, 4.030152e-06, 3.986742e-06, 
    4.015569e-06, 3.968028e-06, 3.981007e-06, 3.878277e-06, 3.839459e-06, 
    3.822998e-06, 3.808625e-06, 3.773745e-06, 3.797817e-06, 3.78832e-06, 
    3.810934e-06, 3.825332e-06, 3.818209e-06, 3.862268e-06, 3.845113e-06, 
    3.93585e-06, 3.896656e-06, 3.999197e-06, 3.974558e-06, 4.005113e-06, 
    3.98951e-06, 4.016259e-06, 3.992182e-06, 4.033931e-06, 4.043045e-06, 
    4.036816e-06, 4.060771e-06, 3.990848e-06, 4.017639e-06, 3.818009e-06, 
    3.81917e-06, 3.824584e-06, 3.800811e-06, 3.79936e-06, 3.777637e-06, 
    3.796964e-06, 3.805206e-06, 3.826169e-06, 3.838589e-06, 3.850413e-06, 
    3.876464e-06, 3.905644e-06, 3.946609e-06, 3.976153e-06, 3.996008e-06, 
    3.983829e-06, 3.994581e-06, 3.982562e-06, 3.976935e-06, 4.039628e-06, 
    4.004373e-06, 4.057322e-06, 4.054385e-06, 4.030393e-06, 4.054716e-06, 
    3.819986e-06, 3.813304e-06, 3.790141e-06, 3.808263e-06, 3.775275e-06, 
    3.793723e-06, 3.804348e-06, 3.845468e-06, 3.854532e-06, 3.86294e-06, 
    3.879572e-06, 3.90096e-06, 3.938599e-06, 3.971475e-06, 4.00159e-06, 
    3.999381e-06, 4.000158e-06, 4.006897e-06, 3.990212e-06, 4.009638e-06, 
    4.012901e-06, 4.004371e-06, 4.053991e-06, 4.039789e-06, 4.054322e-06, 
    4.045073e-06, 3.815476e-06, 3.826725e-06, 3.820645e-06, 3.832081e-06, 
    3.824022e-06, 3.859912e-06, 3.870701e-06, 3.921357e-06, 3.900537e-06, 
    3.933699e-06, 3.903901e-06, 3.909173e-06, 3.934776e-06, 3.90551e-06, 
    3.969657e-06, 3.926114e-06, 4.007158e-06, 3.963497e-06, 4.009901e-06, 
    4.00146e-06, 4.015441e-06, 4.027979e-06, 4.043778e-06, 4.072994e-06, 
    4.066221e-06, 4.090707e-06, 3.843523e-06, 3.858161e-06, 3.856873e-06, 
    3.872217e-06, 3.883581e-06, 3.908263e-06, 3.947986e-06, 3.933029e-06, 
    3.960508e-06, 3.966034e-06, 3.924295e-06, 3.949897e-06, 3.867972e-06, 
    3.881156e-06, 3.873306e-06, 3.844675e-06, 3.93647e-06, 3.889244e-06, 
    3.976641e-06, 3.950917e-06, 4.02619e-06, 3.988678e-06, 4.062495e-06, 
    4.094216e-06, 4.124178e-06, 4.159292e-06, 3.866162e-06, 3.856204e-06, 
    3.874044e-06, 3.89878e-06, 3.921798e-06, 3.952484e-06, 3.955631e-06, 
    3.961392e-06, 3.976334e-06, 3.988916e-06, 3.963212e-06, 3.992072e-06, 
    3.884211e-06, 3.940581e-06, 3.85244e-06, 3.878888e-06, 3.897321e-06, 
    3.889233e-06, 3.931322e-06, 3.941268e-06, 3.981797e-06, 3.960826e-06, 
    4.086375e-06, 4.030626e-06, 4.18612e-06, 4.142418e-06, 3.852727e-06, 
    3.866129e-06, 3.912923e-06, 3.890629e-06, 3.954537e-06, 3.970335e-06, 
    3.983199e-06, 3.999664e-06, 4.001446e-06, 4.011217e-06, 3.99521e-06, 
    4.010585e-06, 3.952549e-06, 3.97844e-06, 3.907566e-06, 3.924765e-06, 
    3.916849e-06, 3.908173e-06, 3.934977e-06, 3.963615e-06, 3.964232e-06, 
    3.973433e-06, 3.999403e-06, 3.954797e-06, 4.093586e-06, 4.007629e-06, 
    3.880766e-06, 3.906672e-06, 3.910383e-06, 3.900334e-06, 3.968749e-06, 
    3.943901e-06, 4.010979e-06, 3.992804e-06, 4.022603e-06, 4.007783e-06, 
    4.005605e-06, 3.98661e-06, 3.974803e-06, 3.945038e-06, 3.920892e-06, 
    3.901791e-06, 3.906229e-06, 3.927224e-06, 3.965371e-06, 4.001605e-06, 
    3.993655e-06, 4.020335e-06, 3.949889e-06, 3.979362e-06, 3.967958e-06, 
    3.997723e-06, 3.932631e-06, 3.988019e-06, 3.918524e-06, 3.924597e-06, 
    3.943409e-06, 3.981361e-06, 3.989785e-06, 3.99878e-06, 3.993229e-06, 
    3.966342e-06, 3.961946e-06, 3.942952e-06, 3.937713e-06, 3.923275e-06, 
    3.911338e-06, 3.922243e-06, 3.933709e-06, 3.966355e-06, 3.99587e-06, 
    4.028157e-06, 4.036076e-06, 4.073958e-06, 4.043104e-06, 4.094066e-06, 
    4.050713e-06, 4.125886e-06, 3.991245e-06, 4.049449e-06, 3.944267e-06, 
    3.955543e-06, 3.975969e-06, 4.022994e-06, 3.997583e-06, 4.02731e-06, 
    3.961774e-06, 3.927947e-06, 3.91922e-06, 3.902951e-06, 3.919592e-06, 
    3.918237e-06, 3.934187e-06, 3.929058e-06, 3.967441e-06, 3.946804e-06, 
    4.005549e-06, 4.027076e-06, 4.088136e-06, 4.125754e-06, 4.164202e-06, 
    4.18122e-06, 4.186406e-06, 4.188575e-06,
  3.868289e-06, 3.905089e-06, 3.897922e-06, 3.927699e-06, 3.911168e-06, 
    3.930686e-06, 3.875737e-06, 3.906553e-06, 3.886867e-06, 3.871596e-06, 
    3.985798e-06, 3.929031e-06, 4.045185e-06, 4.008674e-06, 4.100695e-06, 
    4.039493e-06, 4.11309e-06, 4.098924e-06, 4.141632e-06, 4.129376e-06, 
    4.184231e-06, 4.147295e-06, 4.212805e-06, 4.175396e-06, 4.181238e-06, 
    4.146079e-06, 3.940424e-06, 3.978709e-06, 3.938161e-06, 3.943608e-06, 
    3.941163e-06, 3.911509e-06, 3.896605e-06, 3.865484e-06, 3.871125e-06, 
    3.893987e-06, 3.946059e-06, 3.928346e-06, 3.973062e-06, 3.972049e-06, 
    4.022112e-06, 3.999502e-06, 4.084099e-06, 4.059968e-06, 4.129887e-06, 
    4.112249e-06, 4.129057e-06, 4.123957e-06, 4.129124e-06, 4.103271e-06, 
    4.114338e-06, 4.091624e-06, 4.003732e-06, 4.029467e-06, 3.952947e-06, 
    3.907276e-06, 3.877085e-06, 3.85573e-06, 3.858745e-06, 3.864497e-06, 
    3.894121e-06, 3.922074e-06, 3.943442e-06, 3.957765e-06, 3.971904e-06, 
    4.014845e-06, 4.037665e-06, 4.088986e-06, 4.079702e-06, 4.095436e-06, 
    4.110496e-06, 4.135839e-06, 4.131663e-06, 4.142846e-06, 4.095021e-06, 
    4.126776e-06, 4.074418e-06, 4.088706e-06, 3.975748e-06, 3.933121e-06, 
    3.915066e-06, 3.899299e-06, 3.861065e-06, 3.887449e-06, 3.877038e-06, 
    3.90183e-06, 3.917622e-06, 3.909808e-06, 3.958157e-06, 3.939326e-06, 
    4.03902e-06, 3.995931e-06, 4.108738e-06, 4.081607e-06, 4.115254e-06, 
    4.098069e-06, 4.127536e-06, 4.101011e-06, 4.147013e-06, 4.157062e-06, 
    4.150193e-06, 4.176608e-06, 4.099543e-06, 4.129057e-06, 3.909588e-06, 
    3.910863e-06, 3.9168e-06, 3.890731e-06, 3.889139e-06, 3.865329e-06, 
    3.886512e-06, 3.89555e-06, 3.918539e-06, 3.932167e-06, 3.945143e-06, 
    3.973747e-06, 4.005809e-06, 4.050852e-06, 4.083363e-06, 4.105225e-06, 
    4.091813e-06, 4.103653e-06, 4.090418e-06, 4.084222e-06, 4.153294e-06, 
    4.114441e-06, 4.172804e-06, 4.169564e-06, 4.143112e-06, 4.16993e-06, 
    3.911757e-06, 3.904428e-06, 3.879033e-06, 3.8989e-06, 3.86274e-06, 
    3.88296e-06, 3.89461e-06, 3.939719e-06, 3.949664e-06, 3.958895e-06, 
    3.977159e-06, 4.000658e-06, 4.042041e-06, 4.078215e-06, 4.111373e-06, 
    4.108939e-06, 4.109796e-06, 4.117219e-06, 4.098843e-06, 4.12024e-06, 
    4.123836e-06, 4.114437e-06, 4.169131e-06, 4.153469e-06, 4.169496e-06, 
    4.159295e-06, 3.90681e-06, 3.91915e-06, 3.912479e-06, 3.925027e-06, 
    3.916185e-06, 3.955574e-06, 3.967421e-06, 4.023083e-06, 4.000195e-06, 
    4.036652e-06, 4.003891e-06, 4.009687e-06, 4.037843e-06, 4.005658e-06, 
    4.076216e-06, 4.028314e-06, 4.117508e-06, 4.069439e-06, 4.120529e-06, 
    4.111229e-06, 4.126633e-06, 4.140451e-06, 4.157868e-06, 4.190095e-06, 
    4.182622e-06, 4.209643e-06, 3.93758e-06, 3.953649e-06, 3.952234e-06, 
    3.969082e-06, 3.981564e-06, 4.008684e-06, 4.052365e-06, 4.035913e-06, 
    4.066143e-06, 4.072224e-06, 4.026308e-06, 4.054469e-06, 3.964422e-06, 
    3.978904e-06, 3.970279e-06, 3.938847e-06, 4.0397e-06, 3.987788e-06, 
    4.083901e-06, 4.05559e-06, 4.13848e-06, 4.097156e-06, 4.178511e-06, 
    4.213522e-06, 4.246604e-06, 4.285418e-06, 3.962434e-06, 3.9515e-06, 
    3.971088e-06, 3.998266e-06, 4.023564e-06, 4.057314e-06, 4.060775e-06, 
    4.067116e-06, 4.083562e-06, 4.097414e-06, 4.069121e-06, 4.10089e-06, 
    3.982265e-06, 4.044221e-06, 3.947369e-06, 3.976414e-06, 3.996661e-06, 
    3.987774e-06, 4.034035e-06, 4.044975e-06, 4.089579e-06, 4.066492e-06, 
    4.204867e-06, 4.143372e-06, 4.315087e-06, 4.266763e-06, 3.947683e-06, 
    3.962396e-06, 4.013809e-06, 3.989307e-06, 4.059572e-06, 4.076958e-06, 
    4.091119e-06, 4.109253e-06, 4.111214e-06, 4.12198e-06, 4.104346e-06, 
    4.121282e-06, 4.057386e-06, 4.085881e-06, 4.007917e-06, 4.026826e-06, 
    4.018122e-06, 4.008585e-06, 4.038055e-06, 4.069565e-06, 4.070241e-06, 
    4.08037e-06, 4.108978e-06, 4.059858e-06, 4.212834e-06, 4.118038e-06, 
    3.97847e-06, 4.006939e-06, 4.011015e-06, 3.99997e-06, 4.075214e-06, 
    4.047872e-06, 4.121717e-06, 4.101697e-06, 4.134525e-06, 4.118196e-06, 
    4.115796e-06, 4.094876e-06, 4.081876e-06, 4.049124e-06, 4.022568e-06, 
    4.001571e-06, 4.006449e-06, 4.02953e-06, 4.071497e-06, 4.111391e-06, 
    4.102636e-06, 4.132025e-06, 4.054458e-06, 4.086897e-06, 4.074344e-06, 
    4.107114e-06, 4.035476e-06, 4.096438e-06, 4.019963e-06, 4.026641e-06, 
    4.04733e-06, 4.089101e-06, 4.098372e-06, 4.10828e-06, 4.102165e-06, 
    4.072565e-06, 4.067726e-06, 4.046827e-06, 4.041065e-06, 4.025187e-06, 
    4.012063e-06, 4.024052e-06, 4.036662e-06, 4.072578e-06, 4.105076e-06, 
    4.140648e-06, 4.149376e-06, 4.191166e-06, 4.157131e-06, 4.213365e-06, 
    4.165531e-06, 4.248501e-06, 4.099987e-06, 4.164129e-06, 4.048273e-06, 
    4.060679e-06, 4.083164e-06, 4.134961e-06, 4.10696e-06, 4.139717e-06, 
    4.067537e-06, 4.030327e-06, 4.020728e-06, 4.002846e-06, 4.021137e-06, 
    4.019648e-06, 4.037185e-06, 4.031546e-06, 4.073773e-06, 4.051064e-06, 
    4.115736e-06, 4.139458e-06, 4.206807e-06, 4.24835e-06, 4.290841e-06, 
    4.309664e-06, 4.315401e-06, 4.3178e-06,
  4.120485e-06, 4.158958e-06, 4.151462e-06, 4.182611e-06, 4.165315e-06, 
    4.185736e-06, 4.128268e-06, 4.16049e-06, 4.139903e-06, 4.12394e-06, 
    4.243444e-06, 4.184004e-06, 4.305692e-06, 4.267408e-06, 4.363952e-06, 
    4.299723e-06, 4.37697e-06, 4.36209e-06, 4.40696e-06, 4.394078e-06, 
    4.451765e-06, 4.412913e-06, 4.481837e-06, 4.442467e-06, 4.448614e-06, 
    4.411635e-06, 4.195926e-06, 4.236018e-06, 4.193557e-06, 4.199259e-06, 
    4.1967e-06, 4.165673e-06, 4.150088e-06, 4.117552e-06, 4.123448e-06, 
    4.147349e-06, 4.201825e-06, 4.183285e-06, 4.230095e-06, 4.229034e-06, 
    4.281494e-06, 4.257795e-06, 4.346524e-06, 4.321197e-06, 4.394616e-06, 
    4.376085e-06, 4.393744e-06, 4.388385e-06, 4.393814e-06, 4.366655e-06, 
    4.378279e-06, 4.354424e-06, 4.262228e-06, 4.289206e-06, 4.209035e-06, 
    4.161249e-06, 4.129678e-06, 4.10736e-06, 4.110511e-06, 4.116522e-06, 
    4.147489e-06, 4.176724e-06, 4.199083e-06, 4.214078e-06, 4.228882e-06, 
    4.273881e-06, 4.297805e-06, 4.351656e-06, 4.341908e-06, 4.358429e-06, 
    4.374243e-06, 4.400872e-06, 4.396482e-06, 4.408238e-06, 4.357991e-06, 
    4.391348e-06, 4.336361e-06, 4.351361e-06, 4.232918e-06, 4.188282e-06, 
    4.169397e-06, 4.152903e-06, 4.112935e-06, 4.140513e-06, 4.129629e-06, 
    4.155548e-06, 4.172066e-06, 4.163891e-06, 4.214488e-06, 4.194776e-06, 
    4.299225e-06, 4.254054e-06, 4.372397e-06, 4.343907e-06, 4.379242e-06, 
    4.36119e-06, 4.392147e-06, 4.36428e-06, 4.412617e-06, 4.423184e-06, 
    4.415961e-06, 4.443741e-06, 4.362739e-06, 4.393745e-06, 4.163663e-06, 
    4.164996e-06, 4.171206e-06, 4.143945e-06, 4.14228e-06, 4.117391e-06, 
    4.139532e-06, 4.148982e-06, 4.173024e-06, 4.187284e-06, 4.200865e-06, 
    4.230813e-06, 4.264406e-06, 4.311635e-06, 4.345751e-06, 4.368706e-06, 
    4.354622e-06, 4.367055e-06, 4.353158e-06, 4.346652e-06, 4.419223e-06, 
    4.378388e-06, 4.439739e-06, 4.436331e-06, 4.408518e-06, 4.436715e-06, 
    4.165931e-06, 4.158265e-06, 4.131714e-06, 4.152484e-06, 4.114685e-06, 
    4.13582e-06, 4.148001e-06, 4.195189e-06, 4.205596e-06, 4.215261e-06, 
    4.234387e-06, 4.259006e-06, 4.302392e-06, 4.340348e-06, 4.375164e-06, 
    4.372608e-06, 4.373508e-06, 4.381307e-06, 4.362004e-06, 4.38448e-06, 
    4.388259e-06, 4.378383e-06, 4.435874e-06, 4.419405e-06, 4.436258e-06, 
    4.42553e-06, 4.160756e-06, 4.173664e-06, 4.166686e-06, 4.179813e-06, 
    4.170563e-06, 4.211786e-06, 4.224191e-06, 4.282514e-06, 4.258521e-06, 
    4.296741e-06, 4.262394e-06, 4.268469e-06, 4.297994e-06, 4.264245e-06, 
    4.338251e-06, 4.288e-06, 4.381609e-06, 4.331141e-06, 4.384784e-06, 
    4.375013e-06, 4.391196e-06, 4.40572e-06, 4.42403e-06, 4.457932e-06, 
    4.450068e-06, 4.478506e-06, 4.192949e-06, 4.20977e-06, 4.208287e-06, 
    4.225928e-06, 4.239002e-06, 4.267417e-06, 4.313221e-06, 4.295963e-06, 
    4.327676e-06, 4.334059e-06, 4.285891e-06, 4.31543e-06, 4.221049e-06, 
    4.236217e-06, 4.227181e-06, 4.194275e-06, 4.299938e-06, 4.245524e-06, 
    4.346316e-06, 4.316604e-06, 4.403647e-06, 4.360235e-06, 4.445743e-06, 
    4.482595e-06, 4.517434e-06, 4.558356e-06, 4.218966e-06, 4.207518e-06, 
    4.228028e-06, 4.256501e-06, 4.283015e-06, 4.318413e-06, 4.322044e-06, 
    4.328698e-06, 4.345959e-06, 4.360503e-06, 4.330804e-06, 4.364153e-06, 
    4.239742e-06, 4.30468e-06, 4.203195e-06, 4.23361e-06, 4.254819e-06, 
    4.245506e-06, 4.293993e-06, 4.305467e-06, 4.352278e-06, 4.328043e-06, 
    4.473484e-06, 4.408793e-06, 4.589654e-06, 4.538685e-06, 4.203522e-06, 
    4.218926e-06, 4.272791e-06, 4.247112e-06, 4.320782e-06, 4.339028e-06, 
    4.353893e-06, 4.372939e-06, 4.374997e-06, 4.386308e-06, 4.367783e-06, 
    4.385575e-06, 4.318489e-06, 4.348394e-06, 4.266612e-06, 4.286436e-06, 
    4.277309e-06, 4.267312e-06, 4.29821e-06, 4.331271e-06, 4.331977e-06, 
    4.342611e-06, 4.37266e-06, 4.321082e-06, 4.481878e-06, 4.382176e-06, 
    4.23576e-06, 4.265592e-06, 4.26986e-06, 4.258284e-06, 4.337197e-06, 
    4.308507e-06, 4.386032e-06, 4.365001e-06, 4.39949e-06, 4.382332e-06, 
    4.379811e-06, 4.357838e-06, 4.344191e-06, 4.309821e-06, 4.281972e-06, 
    4.259961e-06, 4.265074e-06, 4.289272e-06, 4.333298e-06, 4.375185e-06, 
    4.36599e-06, 4.396863e-06, 4.315416e-06, 4.349462e-06, 4.336286e-06, 
    4.370691e-06, 4.295506e-06, 4.359489e-06, 4.279239e-06, 4.286241e-06, 
    4.307939e-06, 4.351778e-06, 4.361509e-06, 4.371916e-06, 4.365492e-06, 
    4.334418e-06, 4.329339e-06, 4.307411e-06, 4.301368e-06, 4.284716e-06, 
    4.270958e-06, 4.283527e-06, 4.296751e-06, 4.33443e-06, 4.368551e-06, 
    4.405927e-06, 4.415102e-06, 4.459064e-06, 4.42326e-06, 4.482437e-06, 
    4.432101e-06, 4.519443e-06, 4.36321e-06, 4.430621e-06, 4.308927e-06, 
    4.321943e-06, 4.345545e-06, 4.399953e-06, 4.370529e-06, 4.404951e-06, 
    4.32914e-06, 4.290109e-06, 4.280041e-06, 4.261298e-06, 4.28047e-06, 
    4.278909e-06, 4.297297e-06, 4.291383e-06, 4.335685e-06, 4.311855e-06, 
    4.379749e-06, 4.404678e-06, 4.475522e-06, 4.519278e-06, 4.564071e-06, 
    4.58393e-06, 4.589984e-06, 4.592517e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.778243, 5.778224, 5.778228, 5.778212, 5.778221, 5.778211, 5.778239, 
    5.778223, 5.778234, 5.778241, 5.778182, 5.778212, 5.778152, 5.778171, 
    5.778123, 5.778154, 5.778117, 5.778124, 5.778103, 5.778109, 5.778081, 
    5.7781, 5.778067, 5.778086, 5.778083, 5.7781, 5.778205, 5.778186, 
    5.778207, 5.778204, 5.778205, 5.778221, 5.778228, 5.778244, 5.778242, 
    5.77823, 5.778203, 5.778212, 5.778189, 5.778189, 5.778163, 5.778175, 
    5.778132, 5.778144, 5.778109, 5.778118, 5.778109, 5.778111, 5.778109, 
    5.778122, 5.778117, 5.778128, 5.778173, 5.77816, 5.778199, 5.778223, 
    5.778238, 5.77825, 5.778248, 5.778245, 5.77823, 5.778215, 5.778204, 
    5.778197, 5.778189, 5.778167, 5.778155, 5.77813, 5.778134, 5.778126, 
    5.778119, 5.778106, 5.778108, 5.778102, 5.778126, 5.77811, 5.778137, 
    5.77813, 5.778187, 5.778209, 5.778219, 5.778227, 5.778247, 5.778233, 
    5.778238, 5.778225, 5.778217, 5.778222, 5.778196, 5.778206, 5.778155, 
    5.778177, 5.778119, 5.778133, 5.778116, 5.778125, 5.77811, 5.778123, 
    5.7781, 5.778095, 5.778098, 5.778085, 5.778124, 5.778109, 5.778222, 
    5.778221, 5.778218, 5.778232, 5.778232, 5.778244, 5.778234, 5.778229, 
    5.778217, 5.77821, 5.778203, 5.778188, 5.778172, 5.778149, 5.778132, 
    5.778121, 5.778128, 5.778122, 5.778129, 5.778132, 5.778097, 5.778116, 
    5.778087, 5.778089, 5.778102, 5.778089, 5.778221, 5.778224, 5.778237, 
    5.778227, 5.778246, 5.778235, 5.778229, 5.778206, 5.778201, 5.778196, 
    5.778187, 5.778174, 5.778153, 5.778135, 5.778118, 5.778119, 5.778119, 
    5.778115, 5.778124, 5.778113, 5.778111, 5.778116, 5.778089, 5.778097, 
    5.778089, 5.778094, 5.778223, 5.778217, 5.77822, 5.778214, 5.778218, 
    5.778198, 5.778192, 5.778163, 5.778175, 5.778156, 5.778173, 5.77817, 
    5.778155, 5.778172, 5.778136, 5.77816, 5.778115, 5.778139, 5.778113, 
    5.778118, 5.77811, 5.778103, 5.778094, 5.778078, 5.778082, 5.778069, 
    5.778207, 5.778199, 5.7782, 5.778191, 5.778184, 5.778171, 5.778148, 
    5.778156, 5.778141, 5.778138, 5.778162, 5.778147, 5.778193, 5.778186, 
    5.77819, 5.778206, 5.778154, 5.778181, 5.778132, 5.778146, 5.778104, 
    5.778125, 5.778084, 5.778067, 5.77805, 5.77803, 5.778194, 5.7782, 
    5.77819, 5.778176, 5.778163, 5.778145, 5.778144, 5.778141, 5.778132, 
    5.778125, 5.77814, 5.778123, 5.778184, 5.778152, 5.778202, 5.778187, 
    5.778177, 5.778181, 5.778157, 5.778152, 5.778129, 5.778141, 5.778071, 
    5.778102, 5.778016, 5.77804, 5.778202, 5.778194, 5.778168, 5.77818, 
    5.778144, 5.778135, 5.778128, 5.778119, 5.778118, 5.778112, 5.778121, 
    5.778113, 5.778145, 5.778131, 5.778171, 5.778161, 5.778165, 5.778171, 
    5.778155, 5.778139, 5.778139, 5.778134, 5.778119, 5.778144, 5.778067, 
    5.778115, 5.778186, 5.778171, 5.778169, 5.778175, 5.778136, 5.77815, 
    5.778113, 5.778123, 5.778106, 5.778114, 5.778116, 5.778126, 5.778133, 
    5.77815, 5.778163, 5.778174, 5.778172, 5.77816, 5.778138, 5.778118, 
    5.778122, 5.778108, 5.778147, 5.778131, 5.778137, 5.77812, 5.778157, 
    5.778126, 5.778164, 5.778161, 5.778151, 5.778129, 5.778125, 5.77812, 
    5.778122, 5.778138, 5.77814, 5.778151, 5.778154, 5.778162, 5.778169, 
    5.778162, 5.778156, 5.778138, 5.778121, 5.778103, 5.778099, 5.778078, 
    5.778095, 5.778067, 5.77809, 5.778049, 5.778124, 5.778091, 5.77815, 
    5.778144, 5.778132, 5.778106, 5.77812, 5.778104, 5.77814, 5.778159, 
    5.778164, 5.778173, 5.778164, 5.778165, 5.778156, 5.778159, 5.778137, 
    5.778149, 5.778116, 5.778104, 5.77807, 5.778049, 5.778028, 5.778018, 
    5.778016, 5.778015 ;

 SOIL1C_TO_SOIL2C =
  3.09681e-08, 3.110459e-08, 3.107806e-08, 3.118815e-08, 3.112708e-08, 
    3.119917e-08, 3.099577e-08, 3.111001e-08, 3.103709e-08, 3.098039e-08, 
    3.140179e-08, 3.119306e-08, 3.161866e-08, 3.148552e-08, 3.181999e-08, 
    3.159794e-08, 3.186477e-08, 3.181359e-08, 3.196764e-08, 3.192351e-08, 
    3.212053e-08, 3.198801e-08, 3.222268e-08, 3.208889e-08, 3.210981e-08, 
    3.198364e-08, 3.123507e-08, 3.137581e-08, 3.122673e-08, 3.12468e-08, 
    3.12378e-08, 3.112834e-08, 3.107318e-08, 3.095767e-08, 3.097864e-08, 
    3.106348e-08, 3.125583e-08, 3.119054e-08, 3.13551e-08, 3.135138e-08, 
    3.153459e-08, 3.145199e-08, 3.175994e-08, 3.167241e-08, 3.192535e-08, 
    3.186173e-08, 3.192236e-08, 3.190398e-08, 3.19226e-08, 3.182931e-08, 
    3.186927e-08, 3.178718e-08, 3.146745e-08, 3.156141e-08, 3.128118e-08, 
    3.111268e-08, 3.100078e-08, 3.092138e-08, 3.09326e-08, 3.0954e-08, 
    3.106398e-08, 3.116739e-08, 3.124619e-08, 3.129891e-08, 3.135085e-08, 
    3.150806e-08, 3.159128e-08, 3.177763e-08, 3.174401e-08, 3.180098e-08, 
    3.185541e-08, 3.194679e-08, 3.193175e-08, 3.1972e-08, 3.179948e-08, 
    3.191414e-08, 3.172486e-08, 3.177662e-08, 3.136494e-08, 3.120815e-08, 
    3.114149e-08, 3.108316e-08, 3.094123e-08, 3.103924e-08, 3.10006e-08, 
    3.109253e-08, 3.115094e-08, 3.112205e-08, 3.130035e-08, 3.123103e-08, 
    3.159622e-08, 3.143892e-08, 3.184906e-08, 3.175091e-08, 3.187258e-08, 
    3.18105e-08, 3.191688e-08, 3.182114e-08, 3.198699e-08, 3.20231e-08, 
    3.199843e-08, 3.209323e-08, 3.181583e-08, 3.192236e-08, 3.112124e-08, 
    3.112595e-08, 3.11479e-08, 3.105141e-08, 3.104551e-08, 3.09571e-08, 
    3.103577e-08, 3.106927e-08, 3.115433e-08, 3.120463e-08, 3.125246e-08, 
    3.135761e-08, 3.147505e-08, 3.163927e-08, 3.175727e-08, 3.183637e-08, 
    3.178787e-08, 3.183069e-08, 3.178282e-08, 3.176039e-08, 3.200957e-08, 
    3.186965e-08, 3.20796e-08, 3.206798e-08, 3.197296e-08, 3.206929e-08, 
    3.112926e-08, 3.110215e-08, 3.100801e-08, 3.108168e-08, 3.094747e-08, 
    3.102259e-08, 3.106578e-08, 3.123247e-08, 3.12691e-08, 3.130306e-08, 
    3.137013e-08, 3.145621e-08, 3.160722e-08, 3.173862e-08, 3.185858e-08, 
    3.184979e-08, 3.185288e-08, 3.187968e-08, 3.18133e-08, 3.189057e-08, 
    3.190354e-08, 3.186963e-08, 3.206642e-08, 3.20102e-08, 3.206773e-08, 
    3.203113e-08, 3.111096e-08, 3.115658e-08, 3.113193e-08, 3.117828e-08, 
    3.114563e-08, 3.129084e-08, 3.133438e-08, 3.153813e-08, 3.145452e-08, 
    3.15876e-08, 3.146804e-08, 3.148922e-08, 3.159193e-08, 3.14745e-08, 
    3.173137e-08, 3.155721e-08, 3.188072e-08, 3.170678e-08, 3.189162e-08, 
    3.185806e-08, 3.191363e-08, 3.196339e-08, 3.2026e-08, 3.214152e-08, 
    3.211478e-08, 3.221139e-08, 3.122459e-08, 3.128376e-08, 3.127856e-08, 
    3.134049e-08, 3.138629e-08, 3.148556e-08, 3.164478e-08, 3.158491e-08, 
    3.169483e-08, 3.17169e-08, 3.15499e-08, 3.165243e-08, 3.132337e-08, 
    3.137653e-08, 3.134488e-08, 3.122926e-08, 3.15987e-08, 3.140909e-08, 
    3.175922e-08, 3.16565e-08, 3.195629e-08, 3.180719e-08, 3.210005e-08, 
    3.222524e-08, 3.234308e-08, 3.248078e-08, 3.131607e-08, 3.127586e-08, 
    3.134786e-08, 3.144746e-08, 3.153989e-08, 3.166277e-08, 3.167534e-08, 
    3.169836e-08, 3.1758e-08, 3.180813e-08, 3.170564e-08, 3.18207e-08, 
    3.138885e-08, 3.161515e-08, 3.126065e-08, 3.136739e-08, 3.144159e-08, 
    3.140904e-08, 3.157806e-08, 3.16179e-08, 3.177978e-08, 3.16961e-08, 
    3.219433e-08, 3.197389e-08, 3.258564e-08, 3.241468e-08, 3.126181e-08, 
    3.131593e-08, 3.150428e-08, 3.141466e-08, 3.167097e-08, 3.173406e-08, 
    3.178536e-08, 3.185092e-08, 3.1858e-08, 3.189685e-08, 3.183319e-08, 
    3.189433e-08, 3.166303e-08, 3.176639e-08, 3.148276e-08, 3.155179e-08, 
    3.152003e-08, 3.14852e-08, 3.159271e-08, 3.170725e-08, 3.17097e-08, 
    3.174643e-08, 3.184991e-08, 3.167201e-08, 3.222277e-08, 3.188261e-08, 
    3.137494e-08, 3.147918e-08, 3.149407e-08, 3.145369e-08, 3.172774e-08, 
    3.162844e-08, 3.18959e-08, 3.182361e-08, 3.194205e-08, 3.18832e-08, 
    3.187454e-08, 3.179895e-08, 3.175189e-08, 3.163299e-08, 3.153626e-08, 
    3.145955e-08, 3.147739e-08, 3.156165e-08, 3.171426e-08, 3.185864e-08, 
    3.182701e-08, 3.193306e-08, 3.165239e-08, 3.177007e-08, 3.172458e-08, 
    3.184319e-08, 3.158332e-08, 3.180459e-08, 3.152675e-08, 3.155111e-08, 
    3.162647e-08, 3.177805e-08, 3.18116e-08, 3.18474e-08, 3.182531e-08, 
    3.171813e-08, 3.170058e-08, 3.162464e-08, 3.160367e-08, 3.154581e-08, 
    3.149791e-08, 3.154167e-08, 3.158764e-08, 3.171818e-08, 3.183582e-08, 
    3.19641e-08, 3.199549e-08, 3.214535e-08, 3.202335e-08, 3.222467e-08, 
    3.205349e-08, 3.234982e-08, 3.181743e-08, 3.204847e-08, 3.16299e-08, 
    3.167499e-08, 3.175655e-08, 3.194362e-08, 3.184264e-08, 3.196074e-08, 
    3.169989e-08, 3.156455e-08, 3.152954e-08, 3.146421e-08, 3.153104e-08, 
    3.15256e-08, 3.158954e-08, 3.156899e-08, 3.172251e-08, 3.164005e-08, 
    3.187432e-08, 3.195981e-08, 3.220127e-08, 3.234928e-08, 3.249998e-08, 
    3.256651e-08, 3.258675e-08, 3.259522e-08 ;

 SOIL1C_TO_SOIL3C =
  3.673164e-10, 3.689359e-10, 3.686211e-10, 3.699273e-10, 3.692028e-10, 
    3.700581e-10, 3.676447e-10, 3.690002e-10, 3.681349e-10, 3.674622e-10, 
    3.724624e-10, 3.699857e-10, 3.750357e-10, 3.734559e-10, 3.774246e-10, 
    3.747898e-10, 3.77956e-10, 3.773487e-10, 3.791767e-10, 3.78653e-10, 
    3.80991e-10, 3.794184e-10, 3.822031e-10, 3.806155e-10, 3.808638e-10, 
    3.793665e-10, 3.704841e-10, 3.72154e-10, 3.703852e-10, 3.706233e-10, 
    3.705165e-10, 3.692177e-10, 3.685632e-10, 3.671926e-10, 3.674415e-10, 
    3.684481e-10, 3.707304e-10, 3.699557e-10, 3.719083e-10, 3.718642e-10, 
    3.740381e-10, 3.730579e-10, 3.767121e-10, 3.756735e-10, 3.786749e-10, 
    3.7792e-10, 3.786394e-10, 3.784213e-10, 3.786422e-10, 3.775352e-10, 
    3.780095e-10, 3.770354e-10, 3.732415e-10, 3.743564e-10, 3.710312e-10, 
    3.690319e-10, 3.677042e-10, 3.66762e-10, 3.668952e-10, 3.671491e-10, 
    3.68454e-10, 3.69681e-10, 3.706161e-10, 3.712415e-10, 3.718579e-10, 
    3.737233e-10, 3.747108e-10, 3.76922e-10, 3.765231e-10, 3.77199e-10, 
    3.778449e-10, 3.789292e-10, 3.787508e-10, 3.792285e-10, 3.771813e-10, 
    3.785418e-10, 3.762958e-10, 3.769101e-10, 3.720251e-10, 3.701647e-10, 
    3.693737e-10, 3.686816e-10, 3.669976e-10, 3.681605e-10, 3.677021e-10, 
    3.687928e-10, 3.694858e-10, 3.691431e-10, 3.712586e-10, 3.704362e-10, 
    3.747694e-10, 3.729028e-10, 3.777696e-10, 3.766049e-10, 3.780487e-10, 
    3.77312e-10, 3.785743e-10, 3.774383e-10, 3.794063e-10, 3.798348e-10, 
    3.79542e-10, 3.80667e-10, 3.773753e-10, 3.786393e-10, 3.691334e-10, 
    3.691893e-10, 3.694498e-10, 3.683049e-10, 3.682349e-10, 3.671858e-10, 
    3.681193e-10, 3.685168e-10, 3.69526e-10, 3.701229e-10, 3.706904e-10, 
    3.719381e-10, 3.733316e-10, 3.752803e-10, 3.766804e-10, 3.77619e-10, 
    3.770435e-10, 3.775516e-10, 3.769836e-10, 3.767174e-10, 3.796742e-10, 
    3.780139e-10, 3.805052e-10, 3.803674e-10, 3.792399e-10, 3.803829e-10, 
    3.692286e-10, 3.689069e-10, 3.6779e-10, 3.686641e-10, 3.670716e-10, 
    3.679629e-10, 3.684754e-10, 3.704533e-10, 3.708879e-10, 3.712908e-10, 
    3.720867e-10, 3.731081e-10, 3.748999e-10, 3.764591e-10, 3.778825e-10, 
    3.777782e-10, 3.778149e-10, 3.781329e-10, 3.773452e-10, 3.782622e-10, 
    3.784161e-10, 3.780137e-10, 3.803489e-10, 3.796817e-10, 3.803644e-10, 
    3.799301e-10, 3.690115e-10, 3.695528e-10, 3.692603e-10, 3.698103e-10, 
    3.694228e-10, 3.711459e-10, 3.716625e-10, 3.740801e-10, 3.73088e-10, 
    3.746671e-10, 3.732484e-10, 3.734998e-10, 3.747185e-10, 3.733251e-10, 
    3.76373e-10, 3.743065e-10, 3.781452e-10, 3.760813e-10, 3.782746e-10, 
    3.778763e-10, 3.785357e-10, 3.791263e-10, 3.798692e-10, 3.812401e-10, 
    3.809227e-10, 3.820692e-10, 3.703598e-10, 3.710619e-10, 3.710001e-10, 
    3.717349e-10, 3.722784e-10, 3.734563e-10, 3.753456e-10, 3.746352e-10, 
    3.759395e-10, 3.762013e-10, 3.742197e-10, 3.754363e-10, 3.715318e-10, 
    3.721626e-10, 3.717871e-10, 3.704152e-10, 3.747988e-10, 3.72549e-10, 
    3.767036e-10, 3.754847e-10, 3.79042e-10, 3.772728e-10, 3.807479e-10, 
    3.822334e-10, 3.836319e-10, 3.852659e-10, 3.714452e-10, 3.709681e-10, 
    3.718224e-10, 3.730042e-10, 3.74101e-10, 3.75559e-10, 3.757083e-10, 
    3.759814e-10, 3.76689e-10, 3.772839e-10, 3.760677e-10, 3.774331e-10, 
    3.723087e-10, 3.749941e-10, 3.707877e-10, 3.720542e-10, 3.729345e-10, 
    3.725484e-10, 3.74554e-10, 3.750266e-10, 3.769475e-10, 3.759546e-10, 
    3.818667e-10, 3.792509e-10, 3.865103e-10, 3.844814e-10, 3.708014e-10, 
    3.714435e-10, 3.736784e-10, 3.726151e-10, 3.756564e-10, 3.76405e-10, 
    3.770137e-10, 3.777917e-10, 3.778757e-10, 3.783366e-10, 3.775813e-10, 
    3.783068e-10, 3.755621e-10, 3.767887e-10, 3.73423e-10, 3.742422e-10, 
    3.738654e-10, 3.73452e-10, 3.747277e-10, 3.760869e-10, 3.76116e-10, 
    3.765518e-10, 3.777797e-10, 3.756687e-10, 3.822042e-10, 3.781678e-10, 
    3.721438e-10, 3.733806e-10, 3.735574e-10, 3.730782e-10, 3.7633e-10, 
    3.751517e-10, 3.783254e-10, 3.774677e-10, 3.788731e-10, 3.781747e-10, 
    3.78072e-10, 3.77175e-10, 3.766165e-10, 3.752057e-10, 3.740579e-10, 
    3.731477e-10, 3.733594e-10, 3.743592e-10, 3.7617e-10, 3.778833e-10, 
    3.775079e-10, 3.787663e-10, 3.754359e-10, 3.768323e-10, 3.762926e-10, 
    3.777e-10, 3.746163e-10, 3.772419e-10, 3.739451e-10, 3.742342e-10, 
    3.751283e-10, 3.76927e-10, 3.77325e-10, 3.777499e-10, 3.774878e-10, 
    3.76216e-10, 3.760077e-10, 3.751066e-10, 3.748578e-10, 3.741712e-10, 
    3.736028e-10, 3.741221e-10, 3.746675e-10, 3.762166e-10, 3.776126e-10, 
    3.791346e-10, 3.795072e-10, 3.812854e-10, 3.798377e-10, 3.822267e-10, 
    3.801954e-10, 3.837118e-10, 3.773942e-10, 3.801359e-10, 3.75169e-10, 
    3.757041e-10, 3.766719e-10, 3.788917e-10, 3.776933e-10, 3.790948e-10, 
    3.759995e-10, 3.743936e-10, 3.739782e-10, 3.732031e-10, 3.739959e-10, 
    3.739314e-10, 3.746902e-10, 3.744464e-10, 3.76268e-10, 3.752895e-10, 
    3.780694e-10, 3.790838e-10, 3.81949e-10, 3.837055e-10, 3.854937e-10, 
    3.862832e-10, 3.865235e-10, 3.866239e-10 ;

 SOIL1C_vr =
  19.98125, 19.98119, 19.9812, 19.98116, 19.98118, 19.98116, 19.98124, 
    19.98119, 19.98122, 19.98124, 19.98108, 19.98116, 19.981, 19.98105, 
    19.98092, 19.98101, 19.98091, 19.98093, 19.98087, 19.98088, 19.98081, 
    19.98086, 19.98077, 19.98082, 19.98081, 19.98086, 19.98114, 19.98109, 
    19.98115, 19.98114, 19.98114, 19.98118, 19.9812, 19.98125, 19.98124, 
    19.98121, 19.98114, 19.98116, 19.9811, 19.9811, 19.98103, 19.98106, 
    19.98095, 19.98098, 19.98088, 19.98091, 19.98088, 19.98089, 19.98088, 
    19.98092, 19.98091, 19.98094, 19.98106, 19.98102, 19.98113, 19.98119, 
    19.98123, 19.98126, 19.98126, 19.98125, 19.98121, 19.98117, 19.98114, 
    19.98112, 19.9811, 19.98104, 19.98101, 19.98094, 19.98095, 19.98093, 
    19.98091, 19.98088, 19.98088, 19.98087, 19.98093, 19.98089, 19.98096, 
    19.98094, 19.98109, 19.98115, 19.98118, 19.9812, 19.98125, 19.98122, 
    19.98123, 19.9812, 19.98118, 19.98119, 19.98112, 19.98115, 19.98101, 
    19.98107, 19.98091, 19.98095, 19.9809, 19.98093, 19.98089, 19.98092, 
    19.98086, 19.98085, 19.98086, 19.98082, 19.98092, 19.98088, 19.98119, 
    19.98119, 19.98118, 19.98121, 19.98122, 19.98125, 19.98122, 19.98121, 
    19.98117, 19.98116, 19.98114, 19.9811, 19.98105, 19.98099, 19.98095, 
    19.98092, 19.98094, 19.98092, 19.98094, 19.98095, 19.98085, 19.98091, 
    19.98083, 19.98083, 19.98087, 19.98083, 19.98118, 19.98119, 19.98123, 
    19.9812, 19.98125, 19.98122, 19.98121, 19.98115, 19.98113, 19.98112, 
    19.98109, 19.98106, 19.981, 19.98095, 19.98091, 19.98091, 19.98091, 
    19.9809, 19.98093, 19.9809, 19.98089, 19.98091, 19.98083, 19.98085, 
    19.98083, 19.98084, 19.98119, 19.98117, 19.98118, 19.98116, 19.98118, 
    19.98112, 19.98111, 19.98103, 19.98106, 19.98101, 19.98106, 19.98105, 
    19.98101, 19.98105, 19.98096, 19.98102, 19.9809, 19.98097, 19.9809, 
    19.98091, 19.98089, 19.98087, 19.98085, 19.9808, 19.98081, 19.98078, 
    19.98115, 19.98112, 19.98113, 19.9811, 19.98109, 19.98105, 19.98099, 
    19.98101, 19.98097, 19.98096, 19.98103, 19.98099, 19.98111, 19.98109, 
    19.9811, 19.98115, 19.98101, 19.98108, 19.98095, 19.98099, 19.98087, 
    19.98093, 19.98082, 19.98077, 19.98073, 19.98067, 19.98111, 19.98113, 
    19.9811, 19.98106, 19.98103, 19.98098, 19.98098, 19.98097, 19.98095, 
    19.98093, 19.98097, 19.98092, 19.98109, 19.981, 19.98113, 19.98109, 
    19.98107, 19.98108, 19.98101, 19.981, 19.98094, 19.98097, 19.98078, 
    19.98087, 19.98063, 19.9807, 19.98113, 19.98111, 19.98104, 19.98108, 
    19.98098, 19.98096, 19.98094, 19.98091, 19.98091, 19.98089, 19.98092, 
    19.9809, 19.98098, 19.98094, 19.98105, 19.98102, 19.98104, 19.98105, 
    19.98101, 19.98097, 19.98096, 19.98095, 19.98091, 19.98098, 19.98077, 
    19.9809, 19.98109, 19.98105, 19.98105, 19.98106, 19.98096, 19.981, 
    19.98089, 19.98092, 19.98088, 19.9809, 19.9809, 19.98093, 19.98095, 
    19.98099, 19.98103, 19.98106, 19.98105, 19.98102, 19.98096, 19.98091, 
    19.98092, 19.98088, 19.98099, 19.98094, 19.98096, 19.98092, 19.98101, 
    19.98093, 19.98103, 19.98102, 19.981, 19.98094, 19.98093, 19.98091, 
    19.98092, 19.98096, 19.98097, 19.981, 19.981, 19.98103, 19.98104, 
    19.98103, 19.98101, 19.98096, 19.98092, 19.98087, 19.98086, 19.9808, 
    19.98085, 19.98077, 19.98083, 19.98072, 19.98092, 19.98084, 19.981, 
    19.98098, 19.98095, 19.98088, 19.98092, 19.98087, 19.98097, 19.98102, 
    19.98103, 19.98106, 19.98103, 19.98104, 19.98101, 19.98102, 19.98096, 
    19.98099, 19.9809, 19.98087, 19.98078, 19.98072, 19.98067, 19.98064, 
    19.98063, 19.98063,
  19.9833, 19.98323, 19.98325, 19.9832, 19.98322, 19.98319, 19.98329, 
    19.98323, 19.98326, 19.98329, 19.9831, 19.98319, 19.983, 19.98306, 
    19.9829, 19.98301, 19.98288, 19.98291, 19.98284, 19.98285, 19.98277, 
    19.98283, 19.98272, 19.98278, 19.98277, 19.98283, 19.98317, 19.98311, 
    19.98318, 19.98317, 19.98317, 19.98322, 19.98325, 19.9833, 19.98329, 
    19.98325, 19.98316, 19.98319, 19.98312, 19.98312, 19.98303, 19.98307, 
    19.98293, 19.98297, 19.98285, 19.98288, 19.98285, 19.98286, 19.98285, 
    19.9829, 19.98288, 19.98292, 19.98307, 19.98302, 19.98315, 19.98323, 
    19.98328, 19.98332, 19.98331, 19.9833, 19.98325, 19.98321, 19.98317, 
    19.98314, 19.98312, 19.98305, 19.98301, 19.98292, 19.98294, 19.98291, 
    19.98289, 19.98285, 19.98285, 19.98283, 19.98291, 19.98286, 19.98295, 
    19.98292, 19.98311, 19.98319, 19.98322, 19.98324, 19.98331, 19.98326, 
    19.98328, 19.98324, 19.98321, 19.98323, 19.98314, 19.98318, 19.98301, 
    19.98308, 19.98289, 19.98293, 19.98288, 19.98291, 19.98286, 19.9829, 
    19.98283, 19.98281, 19.98282, 19.98278, 19.9829, 19.98285, 19.98323, 
    19.98322, 19.98321, 19.98326, 19.98326, 19.9833, 19.98327, 19.98325, 
    19.98321, 19.98319, 19.98317, 19.98312, 19.98306, 19.98299, 19.98293, 
    19.98289, 19.98292, 19.9829, 19.98292, 19.98293, 19.98281, 19.98288, 
    19.98278, 19.98279, 19.98283, 19.98279, 19.98322, 19.98324, 19.98328, 
    19.98325, 19.98331, 19.98327, 19.98325, 19.98318, 19.98316, 19.98314, 
    19.98311, 19.98307, 19.983, 19.98294, 19.98289, 19.98289, 19.98289, 
    19.98288, 19.98291, 19.98287, 19.98286, 19.98288, 19.98279, 19.98281, 
    19.98279, 19.98281, 19.98323, 19.98321, 19.98322, 19.9832, 19.98322, 
    19.98315, 19.98313, 19.98303, 19.98307, 19.98301, 19.98307, 19.98306, 
    19.98301, 19.98306, 19.98294, 19.98302, 19.98288, 19.98296, 19.98287, 
    19.98289, 19.98286, 19.98284, 19.98281, 19.98276, 19.98277, 19.98272, 
    19.98318, 19.98315, 19.98315, 19.98313, 19.9831, 19.98306, 19.98298, 
    19.98301, 19.98296, 19.98295, 19.98303, 19.98298, 19.98313, 19.98311, 
    19.98312, 19.98318, 19.98301, 19.98309, 19.98293, 19.98298, 19.98284, 
    19.98291, 19.98277, 19.98272, 19.98266, 19.9826, 19.98314, 19.98315, 
    19.98312, 19.98308, 19.98303, 19.98298, 19.98297, 19.98296, 19.98293, 
    19.98291, 19.98296, 19.9829, 19.9831, 19.983, 19.98316, 19.98311, 
    19.98308, 19.98309, 19.98302, 19.983, 19.98292, 19.98296, 19.98273, 
    19.98283, 19.98255, 19.98263, 19.98316, 19.98314, 19.98305, 19.98309, 
    19.98297, 19.98294, 19.98292, 19.98289, 19.98289, 19.98287, 19.9829, 
    19.98287, 19.98298, 19.98293, 19.98306, 19.98303, 19.98304, 19.98306, 
    19.98301, 19.98296, 19.98295, 19.98294, 19.98289, 19.98297, 19.98272, 
    19.98287, 19.98311, 19.98306, 19.98305, 19.98307, 19.98295, 19.98299, 
    19.98287, 19.9829, 19.98285, 19.98287, 19.98288, 19.98291, 19.98293, 
    19.98299, 19.98303, 19.98307, 19.98306, 19.98302, 19.98295, 19.98289, 
    19.9829, 19.98285, 19.98298, 19.98293, 19.98295, 19.98289, 19.98301, 
    19.98291, 19.98304, 19.98303, 19.98299, 19.98292, 19.98291, 19.98289, 
    19.9829, 19.98295, 19.98296, 19.98299, 19.983, 19.98303, 19.98305, 
    19.98303, 19.98301, 19.98295, 19.98289, 19.98284, 19.98282, 19.98275, 
    19.98281, 19.98272, 19.9828, 19.98266, 19.9829, 19.9828, 19.98299, 
    19.98297, 19.98293, 19.98285, 19.98289, 19.98284, 19.98296, 19.98302, 
    19.98304, 19.98307, 19.98304, 19.98304, 19.98301, 19.98302, 19.98295, 
    19.98299, 19.98288, 19.98284, 19.98273, 19.98266, 19.98259, 19.98256, 
    19.98255, 19.98255,
  19.98426, 19.98419, 19.9842, 19.98414, 19.98418, 19.98414, 19.98424, 
    19.98418, 19.98422, 19.98425, 19.98404, 19.98414, 19.98392, 19.98399, 
    19.98382, 19.98394, 19.9838, 19.98383, 19.98375, 19.98377, 19.98367, 
    19.98374, 19.98362, 19.98368, 19.98368, 19.98374, 19.98412, 19.98405, 
    19.98413, 19.98411, 19.98412, 19.98417, 19.9842, 19.98426, 19.98425, 
    19.98421, 19.98411, 19.98414, 19.98406, 19.98406, 19.98397, 19.98401, 
    19.98385, 19.9839, 19.98377, 19.9838, 19.98377, 19.98378, 19.98377, 
    19.98382, 19.9838, 19.98384, 19.984, 19.98395, 19.9841, 19.98418, 
    19.98424, 19.98428, 19.98428, 19.98426, 19.98421, 19.98416, 19.98412, 
    19.98409, 19.98406, 19.98398, 19.98394, 19.98384, 19.98386, 19.98383, 
    19.9838, 19.98376, 19.98376, 19.98375, 19.98383, 19.98377, 19.98387, 
    19.98384, 19.98405, 19.98413, 19.98417, 19.9842, 19.98427, 19.98422, 
    19.98424, 19.98419, 19.98416, 19.98418, 19.98409, 19.98412, 19.98394, 
    19.98402, 19.98381, 19.98386, 19.9838, 19.98383, 19.98377, 19.98382, 
    19.98374, 19.98372, 19.98373, 19.98368, 19.98382, 19.98377, 19.98418, 
    19.98418, 19.98417, 19.98421, 19.98422, 19.98426, 19.98422, 19.98421, 
    19.98416, 19.98414, 19.98411, 19.98406, 19.984, 19.98392, 19.98385, 
    19.98381, 19.98384, 19.98382, 19.98384, 19.98385, 19.98373, 19.9838, 
    19.98369, 19.9837, 19.98374, 19.9837, 19.98417, 19.98419, 19.98424, 
    19.9842, 19.98427, 19.98423, 19.98421, 19.98412, 19.9841, 19.98409, 
    19.98405, 19.98401, 19.98393, 19.98386, 19.9838, 19.98381, 19.9838, 
    19.98379, 19.98383, 19.98379, 19.98378, 19.9838, 19.9837, 19.98372, 
    19.9837, 19.98372, 19.98418, 19.98416, 19.98417, 19.98415, 19.98417, 
    19.98409, 19.98407, 19.98397, 19.98401, 19.98394, 19.984, 19.98399, 
    19.98394, 19.984, 19.98387, 19.98396, 19.98379, 19.98388, 19.98379, 
    19.9838, 19.98377, 19.98375, 19.98372, 19.98366, 19.98367, 19.98362, 
    19.98413, 19.9841, 19.9841, 19.98407, 19.98404, 19.98399, 19.98391, 
    19.98394, 19.98389, 19.98388, 19.98396, 19.98391, 19.98408, 19.98405, 
    19.98406, 19.98412, 19.98393, 19.98403, 19.98385, 19.98391, 19.98375, 
    19.98383, 19.98368, 19.98362, 19.98356, 19.98349, 19.98408, 19.9841, 
    19.98406, 19.98401, 19.98396, 19.9839, 19.9839, 19.98388, 19.98385, 
    19.98383, 19.98388, 19.98382, 19.98404, 19.98393, 19.98411, 19.98405, 
    19.98401, 19.98403, 19.98395, 19.98392, 19.98384, 19.98388, 19.98363, 
    19.98374, 19.98343, 19.98352, 19.98411, 19.98408, 19.98398, 19.98403, 
    19.9839, 19.98387, 19.98384, 19.98381, 19.9838, 19.98378, 19.98382, 
    19.98378, 19.9839, 19.98385, 19.98399, 19.98396, 19.98397, 19.98399, 
    19.98394, 19.98388, 19.98388, 19.98386, 19.98381, 19.9839, 19.98362, 
    19.98379, 19.98405, 19.984, 19.98399, 19.98401, 19.98387, 19.98392, 
    19.98378, 19.98382, 19.98376, 19.98379, 19.9838, 19.98383, 19.98386, 
    19.98392, 19.98397, 19.98401, 19.984, 19.98395, 19.98388, 19.9838, 
    19.98382, 19.98376, 19.98391, 19.98385, 19.98387, 19.98381, 19.98394, 
    19.98383, 19.98397, 19.98396, 19.98392, 19.98384, 19.98383, 19.98381, 
    19.98382, 19.98387, 19.98388, 19.98392, 19.98393, 19.98396, 19.98399, 
    19.98396, 19.98394, 19.98387, 19.98381, 19.98375, 19.98373, 19.98366, 
    19.98372, 19.98362, 19.9837, 19.98355, 19.98382, 19.98371, 19.98392, 
    19.9839, 19.98385, 19.98376, 19.98381, 19.98375, 19.98388, 19.98395, 
    19.98397, 19.984, 19.98397, 19.98397, 19.98394, 19.98395, 19.98387, 
    19.98391, 19.9838, 19.98375, 19.98363, 19.98355, 19.98348, 19.98344, 
    19.98343, 19.98343,
  19.98501, 19.98494, 19.98495, 19.98489, 19.98492, 19.98489, 19.98499, 
    19.98493, 19.98497, 19.985, 19.98478, 19.98489, 19.98467, 19.98474, 
    19.98456, 19.98468, 19.98454, 19.98457, 19.98449, 19.98451, 19.98441, 
    19.98447, 19.98435, 19.98442, 19.98441, 19.98448, 19.98487, 19.98479, 
    19.98487, 19.98486, 19.98487, 19.98492, 19.98495, 19.98501, 19.985, 
    19.98496, 19.98486, 19.98489, 19.9848, 19.98481, 19.98471, 19.98475, 
    19.98459, 19.98464, 19.98451, 19.98454, 19.98451, 19.98452, 19.98451, 
    19.98456, 19.98454, 19.98458, 19.98475, 19.9847, 19.98484, 19.98493, 
    19.98499, 19.98503, 19.98503, 19.98501, 19.98496, 19.9849, 19.98486, 
    19.98483, 19.98481, 19.98472, 19.98468, 19.98458, 19.9846, 19.98457, 
    19.98454, 19.9845, 19.9845, 19.98448, 19.98457, 19.98451, 19.98461, 
    19.98458, 19.9848, 19.98488, 19.98492, 19.98495, 19.98502, 19.98497, 
    19.98499, 19.98494, 19.98491, 19.98493, 19.98483, 19.98487, 19.98468, 
    19.98476, 19.98455, 19.9846, 19.98454, 19.98457, 19.98451, 19.98456, 
    19.98448, 19.98446, 19.98447, 19.98442, 19.98456, 19.98451, 19.98493, 
    19.98492, 19.98491, 19.98496, 19.98497, 19.98501, 19.98497, 19.98495, 
    19.98491, 19.98488, 19.98486, 19.9848, 19.98474, 19.98466, 19.98459, 
    19.98455, 19.98458, 19.98456, 19.98458, 19.98459, 19.98446, 19.98454, 
    19.98443, 19.98443, 19.98448, 19.98443, 19.98492, 19.98494, 19.98499, 
    19.98495, 19.98502, 19.98498, 19.98495, 19.98487, 19.98485, 19.98483, 
    19.9848, 19.98475, 19.98467, 19.9846, 19.98454, 19.98455, 19.98454, 
    19.98453, 19.98457, 19.98453, 19.98452, 19.98454, 19.98443, 19.98446, 
    19.98443, 19.98445, 19.98493, 19.98491, 19.98492, 19.9849, 19.98491, 
    19.98484, 19.98482, 19.98471, 19.98475, 19.98468, 19.98475, 19.98474, 
    19.98468, 19.98474, 19.98461, 19.9847, 19.98453, 19.98462, 19.98453, 
    19.98454, 19.98451, 19.98449, 19.98446, 19.98439, 19.98441, 19.98436, 
    19.98487, 19.98484, 19.98484, 19.98481, 19.98479, 19.98474, 19.98465, 
    19.98468, 19.98463, 19.98462, 19.9847, 19.98465, 19.98482, 19.98479, 
    19.98481, 19.98487, 19.98468, 19.98478, 19.98459, 19.98465, 19.98449, 
    19.98457, 19.98442, 19.98435, 19.98429, 19.98422, 19.98483, 19.98485, 
    19.98481, 19.98476, 19.98471, 19.98464, 19.98464, 19.98462, 19.98459, 
    19.98457, 19.98462, 19.98456, 19.98479, 19.98467, 19.98485, 19.9848, 
    19.98476, 19.98478, 19.98469, 19.98467, 19.98458, 19.98463, 19.98437, 
    19.98448, 19.98416, 19.98425, 19.98485, 19.98483, 19.98473, 19.98477, 
    19.98464, 19.98461, 19.98458, 19.98455, 19.98454, 19.98452, 19.98456, 
    19.98452, 19.98464, 19.98459, 19.98474, 19.9847, 19.98472, 19.98474, 
    19.98468, 19.98462, 19.98462, 19.9846, 19.98455, 19.98464, 19.98435, 
    19.98453, 19.98479, 19.98474, 19.98473, 19.98475, 19.98461, 19.98466, 
    19.98452, 19.98456, 19.9845, 19.98453, 19.98453, 19.98457, 19.9846, 
    19.98466, 19.98471, 19.98475, 19.98474, 19.9847, 19.98462, 19.98454, 
    19.98456, 19.9845, 19.98465, 19.98459, 19.98461, 19.98455, 19.98469, 
    19.98457, 19.98471, 19.9847, 19.98466, 19.98458, 19.98457, 19.98455, 
    19.98456, 19.98462, 19.98462, 19.98466, 19.98467, 19.9847, 19.98473, 
    19.98471, 19.98468, 19.98462, 19.98455, 19.98449, 19.98447, 19.98439, 
    19.98446, 19.98435, 19.98444, 19.98429, 19.98456, 19.98444, 19.98466, 
    19.98464, 19.9846, 19.9845, 19.98455, 19.98449, 19.98462, 19.9847, 
    19.98471, 19.98475, 19.98471, 19.98472, 19.98468, 19.98469, 19.98461, 
    19.98466, 19.98453, 19.98449, 19.98436, 19.98429, 19.98421, 19.98417, 
    19.98416, 19.98416,
  19.98609, 19.98602, 19.98603, 19.98598, 19.98601, 19.98598, 19.98607, 
    19.98602, 19.98605, 19.98608, 19.98588, 19.98598, 19.98577, 19.98584, 
    19.98568, 19.98578, 19.98566, 19.98568, 19.98561, 19.98563, 19.98554, 
    19.9856, 19.98549, 19.98555, 19.98554, 19.9856, 19.98596, 19.98589, 
    19.98596, 19.98595, 19.98596, 19.98601, 19.98603, 19.98609, 19.98608, 
    19.98604, 19.98595, 19.98598, 19.9859, 19.9859, 19.98582, 19.98586, 
    19.98571, 19.98575, 19.98563, 19.98566, 19.98563, 19.98564, 19.98563, 
    19.98568, 19.98566, 19.98569, 19.98585, 19.9858, 19.98594, 19.98602, 
    19.98607, 19.98611, 19.9861, 19.98609, 19.98604, 19.98599, 19.98595, 
    19.98593, 19.9859, 19.98583, 19.98579, 19.9857, 19.98572, 19.98569, 
    19.98566, 19.98562, 19.98563, 19.98561, 19.98569, 19.98563, 19.98573, 
    19.9857, 19.9859, 19.98597, 19.986, 19.98603, 19.9861, 19.98605, 
    19.98607, 19.98603, 19.986, 19.98601, 19.98593, 19.98596, 19.98579, 
    19.98586, 19.98567, 19.98571, 19.98565, 19.98568, 19.98563, 19.98568, 
    19.9856, 19.98558, 19.98559, 19.98555, 19.98568, 19.98563, 19.98601, 
    19.98601, 19.986, 19.98605, 19.98605, 19.98609, 19.98605, 19.98604, 
    19.986, 19.98597, 19.98595, 19.9859, 19.98584, 19.98577, 19.98571, 
    19.98567, 19.98569, 19.98567, 19.9857, 19.98571, 19.98559, 19.98566, 
    19.98556, 19.98556, 19.98561, 19.98556, 19.98601, 19.98602, 19.98607, 
    19.98603, 19.9861, 19.98606, 19.98604, 19.98596, 19.98594, 19.98593, 
    19.98589, 19.98585, 19.98578, 19.98572, 19.98566, 19.98567, 19.98566, 
    19.98565, 19.98568, 19.98565, 19.98564, 19.98566, 19.98556, 19.98559, 
    19.98556, 19.98558, 19.98602, 19.986, 19.98601, 19.98598, 19.986, 
    19.98593, 19.98591, 19.98581, 19.98585, 19.98579, 19.98585, 19.98584, 
    19.98579, 19.98584, 19.98572, 19.98581, 19.98565, 19.98573, 19.98565, 
    19.98566, 19.98564, 19.98561, 19.98558, 19.98553, 19.98554, 19.98549, 
    19.98596, 19.98594, 19.98594, 19.98591, 19.98589, 19.98584, 19.98576, 
    19.98579, 19.98574, 19.98573, 19.98581, 19.98576, 19.98592, 19.98589, 
    19.98591, 19.98596, 19.98578, 19.98588, 19.98571, 19.98576, 19.98561, 
    19.98569, 19.98555, 19.98549, 19.98543, 19.98536, 19.98592, 19.98594, 
    19.9859, 19.98586, 19.98581, 19.98575, 19.98575, 19.98574, 19.98571, 
    19.98569, 19.98573, 19.98568, 19.98589, 19.98578, 19.98595, 19.9859, 
    19.98586, 19.98588, 19.98579, 19.98577, 19.9857, 19.98574, 19.9855, 
    19.98561, 19.98531, 19.9854, 19.98594, 19.98592, 19.98583, 19.98587, 
    19.98575, 19.98572, 19.9857, 19.98566, 19.98566, 19.98564, 19.98567, 
    19.98564, 19.98575, 19.9857, 19.98584, 19.98581, 19.98582, 19.98584, 
    19.98579, 19.98573, 19.98573, 19.98571, 19.98566, 19.98575, 19.98549, 
    19.98565, 19.98589, 19.98584, 19.98583, 19.98585, 19.98572, 19.98577, 
    19.98564, 19.98568, 19.98562, 19.98565, 19.98565, 19.98569, 19.98571, 
    19.98577, 19.98582, 19.98585, 19.98584, 19.9858, 19.98573, 19.98566, 
    19.98568, 19.98563, 19.98576, 19.9857, 19.98573, 19.98567, 19.98579, 
    19.98569, 19.98582, 19.98581, 19.98577, 19.9857, 19.98568, 19.98567, 
    19.98568, 19.98573, 19.98574, 19.98577, 19.98578, 19.98581, 19.98583, 
    19.98581, 19.98579, 19.98573, 19.98567, 19.98561, 19.9856, 19.98553, 
    19.98558, 19.98549, 19.98557, 19.98543, 19.98568, 19.98557, 19.98577, 
    19.98575, 19.98571, 19.98562, 19.98567, 19.98561, 19.98574, 19.9858, 
    19.98582, 19.98585, 19.98582, 19.98582, 19.98579, 19.9858, 19.98573, 
    19.98577, 19.98565, 19.98561, 19.9855, 19.98543, 19.98536, 19.98532, 
    19.98531, 19.98531,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222804, 0.722278, 0.7222785, 0.7222765, 0.7222776, 0.7222763, 0.7222799, 
    0.7222779, 0.7222792, 0.7222801, 0.7222728, 0.7222764, 0.7222689, 
    0.7222713, 0.7222654, 0.7222693, 0.7222646, 0.7222655, 0.7222629, 
    0.7222636, 0.7222602, 0.7222625, 0.7222583, 0.7222607, 0.7222604, 
    0.7222626, 0.7222757, 0.7222732, 0.7222759, 0.7222755, 0.7222757, 
    0.7222776, 0.7222785, 0.7222806, 0.7222802, 0.7222787, 0.7222753, 
    0.7222765, 0.7222736, 0.7222736, 0.7222704, 0.7222719, 0.7222665, 
    0.722268, 0.7222636, 0.7222647, 0.7222636, 0.7222639, 0.7222636, 
    0.7222652, 0.7222646, 0.722266, 0.7222716, 0.72227, 0.7222749, 0.7222778, 
    0.7222798, 0.7222812, 0.722281, 0.7222806, 0.7222787, 0.7222769, 
    0.7222755, 0.7222746, 0.7222736, 0.7222709, 0.7222694, 0.7222662, 
    0.7222667, 0.7222658, 0.7222648, 0.7222632, 0.7222635, 0.7222627, 
    0.7222658, 0.7222638, 0.7222671, 0.7222662, 0.7222734, 0.7222762, 
    0.7222773, 0.7222784, 0.7222809, 0.7222791, 0.7222798, 0.7222782, 
    0.7222772, 0.7222777, 0.7222745, 0.7222758, 0.7222694, 0.7222721, 
    0.7222649, 0.7222666, 0.7222645, 0.7222656, 0.7222638, 0.7222654, 
    0.7222625, 0.7222618, 0.7222623, 0.7222607, 0.7222655, 0.7222636, 
    0.7222777, 0.7222776, 0.7222772, 0.722279, 0.722279, 0.7222806, 
    0.7222792, 0.7222786, 0.7222771, 0.7222762, 0.7222754, 0.7222735, 
    0.7222715, 0.7222686, 0.7222666, 0.7222651, 0.722266, 0.7222652, 
    0.7222661, 0.7222665, 0.7222621, 0.7222645, 0.7222609, 0.7222611, 
    0.7222627, 0.7222611, 0.7222776, 0.7222781, 0.7222797, 0.7222784, 
    0.7222807, 0.7222794, 0.7222787, 0.7222757, 0.7222751, 0.7222745, 
    0.7222733, 0.7222718, 0.7222692, 0.7222669, 0.7222648, 0.7222649, 
    0.7222648, 0.7222643, 0.7222655, 0.7222642, 0.7222639, 0.7222645, 
    0.7222611, 0.7222621, 0.7222611, 0.7222617, 0.7222779, 0.7222771, 
    0.7222775, 0.7222767, 0.7222773, 0.7222747, 0.7222739, 0.7222704, 
    0.7222719, 0.7222695, 0.7222716, 0.7222713, 0.7222694, 0.7222715, 
    0.722267, 0.72227, 0.7222643, 0.7222674, 0.7222642, 0.7222648, 0.7222638, 
    0.7222629, 0.7222618, 0.7222598, 0.7222602, 0.7222586, 0.7222759, 
    0.7222748, 0.722275, 0.7222738, 0.7222731, 0.7222713, 0.7222685, 
    0.7222695, 0.7222676, 0.7222672, 0.7222702, 0.7222683, 0.7222741, 
    0.7222732, 0.7222738, 0.7222758, 0.7222693, 0.7222726, 0.7222665, 
    0.7222683, 0.722263, 0.7222657, 0.7222605, 0.7222583, 0.7222562, 
    0.7222538, 0.7222743, 0.722275, 0.7222737, 0.722272, 0.7222704, 
    0.7222682, 0.722268, 0.7222676, 0.7222665, 0.7222657, 0.7222674, 
    0.7222654, 0.722273, 0.722269, 0.7222753, 0.7222733, 0.7222721, 
    0.7222726, 0.7222697, 0.722269, 0.7222661, 0.7222676, 0.7222589, 
    0.7222627, 0.722252, 0.722255, 0.7222753, 0.7222743, 0.722271, 0.7222725, 
    0.722268, 0.7222669, 0.722266, 0.7222649, 0.7222648, 0.7222641, 
    0.7222652, 0.7222641, 0.7222682, 0.7222664, 0.7222713, 0.7222701, 
    0.7222707, 0.7222713, 0.7222694, 0.7222674, 0.7222674, 0.7222667, 
    0.7222649, 0.722268, 0.7222583, 0.7222643, 0.7222732, 0.7222714, 
    0.7222711, 0.7222719, 0.722267, 0.7222688, 0.7222641, 0.7222654, 
    0.7222633, 0.7222643, 0.7222645, 0.7222658, 0.7222666, 0.7222687, 
    0.7222704, 0.7222717, 0.7222714, 0.72227, 0.7222673, 0.7222648, 
    0.7222653, 0.7222635, 0.7222683, 0.7222663, 0.7222671, 0.722265, 
    0.7222696, 0.7222657, 0.7222705, 0.7222701, 0.7222688, 0.7222661, 
    0.7222656, 0.7222649, 0.7222653, 0.7222672, 0.7222675, 0.7222689, 
    0.7222692, 0.7222703, 0.7222711, 0.7222703, 0.7222695, 0.7222672, 
    0.7222651, 0.7222629, 0.7222623, 0.7222597, 0.7222618, 0.7222583, 
    0.7222613, 0.7222561, 0.7222655, 0.7222614, 0.7222688, 0.722268, 
    0.7222666, 0.7222633, 0.722265, 0.722263, 0.7222675, 0.7222699, 
    0.7222705, 0.7222717, 0.7222705, 0.7222706, 0.7222695, 0.7222698, 
    0.7222672, 0.7222686, 0.7222645, 0.722263, 0.7222587, 0.7222561, 
    0.7222535, 0.7222523, 0.722252, 0.7222518 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  3.597945e-20, -1.541976e-20, -2.569961e-20, -2.006177e-36, 5.139921e-21, 
    1.027984e-20, -3.083953e-20, -2.569961e-20, -1.027984e-20, 3.083953e-20, 
    0, 5.139921e-21, 2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -2.006177e-36, -5.139921e-21, 5.139921e-21, -2.055969e-20, 0, 
    -1.027984e-20, -1.541976e-20, -1.541976e-20, -1.027984e-20, 5.139921e-20, 
    -5.139921e-21, -2.006177e-36, 3.083953e-20, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 2.055969e-20, 2.055969e-20, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 2.006177e-36, -3.083953e-20, 
    -1.027984e-20, -5.139921e-21, 0, -4.111937e-20, -3.597945e-20, 
    -1.541976e-20, -1.541976e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -2.055969e-20, 2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    3.597945e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    2.569961e-20, 5.139921e-21, -2.569961e-20, 1.027984e-20, -1.541976e-20, 
    0, -1.027984e-20, 3.597945e-20, 2.006177e-36, -2.006177e-36, 
    -3.597945e-20, 5.139921e-21, -1.027984e-20, -2.569961e-20, 1.027984e-20, 
    -3.083953e-20, -1.027984e-20, 2.055969e-20, 4.111937e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 3.083953e-20, 3.083953e-20, -5.139921e-21, 
    5.139921e-21, -2.006177e-36, -1.541976e-20, 0, 5.139921e-21, 
    1.027984e-20, -5.139921e-20, 0, 0, -5.139921e-21, 2.006177e-36, 
    -5.139921e-21, -2.006177e-36, 2.055969e-20, 0, 5.139921e-21, 
    -3.083953e-20, 1.541976e-20, -5.139921e-21, 3.083953e-20, 1.027984e-20, 
    -2.055969e-20, -1.541976e-20, -4.111937e-20, 2.569961e-20, -2.569961e-20, 
    -1.541976e-20, -2.569961e-20, -2.006177e-36, 2.055969e-20, 5.139921e-21, 
    -1.027984e-20, -6.167906e-20, -1.541976e-20, -1.027984e-20, 0, 
    2.055969e-20, 5.139921e-21, -2.569961e-20, 5.139921e-21, 2.055969e-20, 0, 
    3.083953e-20, 2.006177e-36, -1.541976e-20, 5.139921e-21, 3.083953e-20, 
    5.139921e-21, -2.055969e-20, 0, 1.541976e-20, -3.597945e-20, 
    -1.541976e-20, -3.083953e-20, -2.055969e-20, -1.027984e-20, 1.027984e-20, 
    3.083953e-20, 1.541976e-20, 5.139921e-21, 2.055969e-20, 0, 1.027984e-20, 
    -5.139921e-21, 3.083953e-20, 1.541976e-20, -1.541976e-20, -2.055969e-20, 
    1.541976e-20, 1.541976e-20, 3.597945e-20, -2.006177e-36, 1.027984e-20, 
    -2.055969e-20, 0, 1.027984e-20, -1.027984e-20, 4.111937e-20, 
    1.027984e-20, 5.139921e-21, -2.006177e-36, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 1.027984e-20, -2.569961e-20, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, -2.569961e-20, 1.541976e-20, 3.083953e-20, -2.569961e-20, 
    -2.569961e-20, 2.055969e-20, -4.111937e-20, 0, 5.139921e-21, 
    2.006177e-36, -2.055969e-20, -2.569961e-20, 5.139921e-21, 2.055969e-20, 
    1.541976e-20, 5.139921e-21, 0, 1.541976e-20, 2.055969e-20, -2.569961e-20, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, 3.083953e-20, -2.055969e-20, 5.139921e-21, 
    3.597945e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, 
    1.027984e-20, -1.027984e-20, -2.055969e-20, 2.569961e-20, -1.541976e-20, 
    3.083953e-20, 1.541976e-20, 1.541976e-20, -1.541976e-20, 2.569961e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, -1.027984e-20, -2.055969e-20, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -1.541976e-20, -4.111937e-20, -2.055969e-20, 3.083953e-20, 5.653913e-20, 
    -2.006177e-36, 1.027984e-20, -5.139921e-21, 2.055969e-20, 2.569961e-20, 
    -2.055969e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -2.055969e-20, 0, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 5.139921e-21, 0, -1.541976e-20, 1.027984e-20, 
    1.541976e-20, 5.139921e-21, 2.055969e-20, -5.139921e-21, 1.541976e-20, 
    4.111937e-20, -1.027984e-20, -1.541976e-20, -2.569961e-20, 2.569961e-20, 
    3.083953e-20, -3.597945e-20, -1.541976e-20, 2.055969e-20, -1.541976e-20, 
    1.541976e-20, -3.083953e-20, 5.139921e-21, 2.055969e-20, -1.027984e-20, 
    -2.006177e-36, -3.083953e-20, -4.111937e-20, -2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 2.569961e-20, -2.055969e-20, -2.055969e-20, 5.139921e-21, 
    1.027984e-20, 2.569961e-20, 0, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, 2.055969e-20, 3.083953e-20, 
    5.139921e-21, 1.027984e-20, -2.006177e-36, -4.625929e-20, 1.027984e-20, 
    -1.541976e-20, -2.055969e-20, 2.006177e-36, -1.541976e-20, -1.541976e-20, 
    5.139921e-21, 3.597945e-20, -1.541976e-20, 0, -3.083953e-20, 
    -2.006177e-36, -4.111937e-20, 3.083953e-20, -1.027984e-20, 2.569961e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, -1.541976e-20,
  -1.541976e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, 3.083953e-20, 
    -1.541976e-20, -2.055969e-20, -2.055969e-20, 5.139921e-21, 2.569961e-20, 
    1.027984e-20, 1.541976e-20, 2.006177e-36, -5.139921e-21, 1.027984e-20, 
    3.083953e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    0, -2.569961e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -2.569961e-20, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, -2.055969e-20, 
    -1.541976e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 2.006177e-36, 
    1.541976e-20, -1.027984e-20, 0, 5.139921e-21, -5.139921e-21, 
    1.541976e-20, 0, 2.569961e-20, -1.541976e-20, 0, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 0, 5.139921e-21, -1.541976e-20, 
    -3.083953e-20, 1.541976e-20, 2.055969e-20, 5.139921e-21, 1.027984e-20, 0, 
    3.597945e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 1.541976e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, 0, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 4.625929e-20, -1.027984e-20, 0, 0, -2.569961e-20, 0, 
    -2.569961e-20, -2.055969e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -2.569961e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 0, 2.569961e-20, -1.027984e-20, 2.055969e-20, 2.006177e-36, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 2.006177e-36, 2.006177e-36, 
    2.006177e-36, 2.055969e-20, 2.006177e-36, 1.027984e-20, -5.139921e-21, 0, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-20, 
    0, 5.139921e-21, 0, -3.083953e-20, 1.541976e-20, -3.083953e-20, 
    -5.139921e-21, -3.083953e-20, -1.027984e-20, -2.055969e-20, 
    -1.541976e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.541976e-20, 2.055969e-20, 
    0, -1.541976e-20, -2.055969e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 2.569961e-20, 3.597945e-20, 1.027984e-20, 1.027984e-20, 0, 
    -2.569961e-20, -2.055969e-20, -1.027984e-20, 2.006177e-36, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 2.055969e-20, -1.027984e-20, -2.569961e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, 0, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, -2.006177e-36, -5.139921e-21, 
    0, -1.027984e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -2.006177e-36, -5.139921e-21, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 2.569961e-20, 1.541976e-20, 
    -2.006177e-36, 1.541976e-20, 1.027984e-20, 1.027984e-20, 5.139921e-21, 0, 
    1.027984e-20, 0, 4.111937e-20, 5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 0, 2.569961e-20, 5.139921e-21, 0, 1.027984e-20, 
    -1.541976e-20, 0, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -1.027984e-20, -2.006177e-36, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 1.541976e-20, 2.006177e-36, -1.027984e-20, 
    -1.541976e-20, 0, 2.055969e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 
    2.055969e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 1.541976e-20, 
    2.006177e-36, -1.027984e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    3.597945e-20, 5.139921e-21, -1.541976e-20, 2.569961e-20, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, 3.083953e-20, 4.111937e-20, 
    -2.055969e-20, 2.006177e-36, 0, 5.139921e-21, 1.541976e-20, 
    -2.006177e-36, -5.139921e-21, 2.569961e-20, -1.027984e-20, 2.006177e-36, 
    1.027984e-20, -1.027984e-20, 3.597945e-20, 1.027984e-20, -1.027984e-20, 
    -2.055969e-20, -1.541976e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -3.083953e-20, -1.541976e-20, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, -3.597945e-20, 2.055969e-20, -2.006177e-36, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, 2.006177e-36, -5.139921e-21, 2.569961e-20, 
    -5.139921e-21, -2.055969e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-20, 1.027984e-20, 0, 0, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, 0, -2.569961e-20, 
    1.027984e-20, 1.027984e-20, 3.597945e-20, -3.083953e-20, 1.027984e-20, 0, 
    -2.055969e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 1.541976e-20, 
    -2.055969e-20, -5.139921e-21, 2.055969e-20, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, -1.541976e-20, 2.055969e-20, -2.569961e-20, -3.083953e-20, 
    5.139921e-21, 0, -1.027984e-20, 2.055969e-20, 1.027984e-20, 2.569961e-20, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20,
  -5.139921e-21, -3.597945e-20, 0, 1.027984e-20, -3.597945e-20, 0, 
    -3.597945e-20, 5.139921e-21, 3.083953e-20, 1.027984e-20, 0, 
    -3.597945e-20, -1.541976e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    -1.541976e-20, 3.083953e-20, -1.541976e-20, 2.569961e-20, -1.541976e-20, 
    2.569961e-20, 1.027984e-20, 2.055969e-20, -2.569961e-20, -1.541976e-20, 
    2.569961e-20, -5.139921e-21, -1.541976e-20, -3.597945e-20, 3.083953e-20, 
    5.139921e-21, 1.027984e-20, -2.055969e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, -1.027984e-20, -4.625929e-20, 
    4.111937e-20, -1.027984e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    2.055969e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, -2.569961e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -3.597945e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, -1.541976e-20, -3.083953e-20, 
    1.541976e-20, 1.027984e-20, 5.139921e-21, 3.597945e-20, 2.569961e-20, 
    3.083953e-20, -1.541976e-20, 2.569961e-20, 2.006177e-36, 4.111937e-20, 
    5.139921e-21, 2.055969e-20, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.569961e-20, -5.139921e-21, 2.055969e-20, 
    -5.139921e-21, 5.139921e-21, 0, -2.055969e-20, -1.541976e-20, 
    2.569961e-20, 1.027984e-20, -1.027984e-20, -2.055969e-20, 0, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 0, 
    -2.569961e-20, -1.541976e-20, -5.139921e-21, 2.055969e-20, -1.027984e-20, 
    2.006177e-36, -1.027984e-20, 0, 2.055969e-20, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 
    2.006177e-36, -5.139921e-21, 1.541976e-20, 0, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 4.625929e-20, 3.083953e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, 1.027984e-20, 4.111937e-20, 
    1.027984e-20, 2.006177e-36, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    -2.055969e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 0, 5.139921e-21, -5.139921e-21, -1.027984e-20, 0, 
    2.006177e-36, -2.055969e-20, 3.083953e-20, 1.541976e-20, 0, 
    -2.569961e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    2.569961e-20, -5.139921e-21, -1.541976e-20, 0, 2.006177e-36, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 0, 3.597945e-20, 5.139921e-21, 
    4.625929e-20, 1.541976e-20, 0, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -2.006177e-36, -3.597945e-20, 5.139921e-21, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, 3.083953e-20, -3.597945e-20, 
    -5.139921e-21, 5.139921e-21, 2.569961e-20, 1.541976e-20, -1.541976e-20, 
    1.541976e-20, -5.139921e-21, -2.055969e-20, 0, 2.006177e-36, 
    1.541976e-20, -1.027984e-20, -2.055969e-20, -2.569961e-20, 1.541976e-20, 
    -2.569961e-20, -2.055969e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 4.111937e-20, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-20, -5.139921e-21, 
    -2.006177e-36, 1.027984e-20, 2.006177e-36, 0, 5.139921e-21, 1.541976e-20, 
    -1.027984e-20, 1.027984e-20, -3.083953e-20, 0, -3.083953e-20, 
    -5.139921e-21, -2.569961e-20, 5.139921e-21, 2.569961e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    0, 1.541976e-20, 0, 1.027984e-20, 3.083953e-20, 3.083953e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    0, -2.055969e-20, 5.139921e-21, -1.027984e-20, 3.597945e-20, 
    -5.139921e-21, 2.055969e-20, -2.055969e-20, 0, 3.597945e-20, 
    5.139921e-21, 3.597945e-20, 5.139921e-21, 1.027984e-20, -2.055969e-20, 
    -1.027984e-20, 0, -3.597945e-20, -5.139921e-21, 5.139921e-21, 
    -2.569961e-20, 2.055969e-20, -3.597945e-20, -2.569961e-20, 2.006177e-36, 
    -2.055969e-20, 2.055969e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    3.597945e-20, 1.541976e-20, 1.541976e-20, 0, 1.027984e-20, -2.006177e-36, 
    -1.541976e-20, 5.139921e-21, -2.006177e-36, 1.027984e-20, -1.541976e-20, 
    0, 0, 1.027984e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, 0, 1.027984e-20, -5.139921e-21, 0, 1.541976e-20, 
    2.055969e-20, 5.139921e-21, 5.139921e-21, -4.625929e-20, -2.055969e-20, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -2.006177e-36, 2.006177e-36, 
    3.083953e-20, 0,
  5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -2.055969e-20, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.027984e-20, -2.569961e-20, 
    1.541976e-20, -1.027984e-20, -2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -3.597945e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, -1.027984e-20, 
    0, 0, -5.139921e-21, -1.541976e-20, -2.006177e-36, 1.027984e-20, 
    1.541976e-20, -2.006177e-36, -1.027984e-20, 1.027984e-20, 3.597945e-20, 
    -2.055969e-20, 1.541976e-20, 4.111937e-20, -1.027984e-20, 1.541976e-20, 
    -2.569961e-20, -1.027984e-20, -3.083953e-20, -1.027984e-20, 
    -2.055969e-20, 2.055969e-20, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -4.111937e-20, -5.139921e-21, 1.027984e-20, 2.569961e-20, -2.569961e-20, 
    -5.139921e-21, 1.027984e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, -1.027984e-20, 2.055969e-20, 
    -1.027984e-20, 0, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -3.083953e-20, 2.569961e-20, 2.055969e-20, 3.597945e-20, -2.055969e-20, 
    -1.027984e-20, -2.055969e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, 5.139921e-21, -3.597945e-20, 5.139921e-21, 
    -5.139921e-21, -2.569961e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, 
    3.083953e-20, 1.541976e-20, 0, 0, -5.139921e-21, 1.027984e-20, 
    -4.625929e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    2.055969e-20, 1.027984e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, 
    5.139921e-21, -2.569961e-20, 1.027984e-20, 1.541976e-20, 2.006177e-36, 
    2.055969e-20, -5.139921e-21, 1.027984e-20, 2.006177e-36, -5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, 0, -5.139921e-21, 
    -1.027984e-20, 4.111937e-20, -1.541976e-20, 0, -2.055969e-20, 
    2.569961e-20, -2.569961e-20, -5.139921e-21, -2.569961e-20, -1.027984e-20, 
    -1.027984e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, 0, 
    -1.027984e-20, 5.139921e-21, -3.083953e-20, -4.625929e-20, 3.083953e-20, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, -2.055969e-20, 4.625929e-20, 
    1.027984e-20, -2.055969e-20, 3.083953e-20, -1.027984e-20, -1.027984e-20, 
    -2.006177e-36, -1.027984e-20, 1.027984e-20, 0, -1.027984e-20, 
    -2.006177e-36, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-20, -2.055969e-20, 
    2.006177e-36, -2.006177e-36, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, -2.055969e-20, -1.027984e-20, 
    5.139921e-21, 0, -5.139921e-21, 2.569961e-20, 3.083953e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, 
    -1.027984e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, -2.055969e-20, 
    -5.139921e-21, -3.083953e-20, -3.083953e-20, -1.541976e-20, 2.006177e-36, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, 2.569961e-20, 1.027984e-20, 
    5.139921e-21, -2.055969e-20, 2.569961e-20, -2.055969e-20, -2.055969e-20, 
    -1.027984e-20, -1.027984e-20, -2.055969e-20, -3.597945e-20, 0, 
    -5.139921e-21, 2.055969e-20, -2.006177e-36, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, 2.006177e-36, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, -4.625929e-20, 5.139921e-21, 2.055969e-20, 
    1.027984e-20, 2.055969e-20, -4.111937e-20, 2.055969e-20, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 2.055969e-20, -1.027984e-20, -2.569961e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 0, -2.055969e-20, -2.569961e-20, 
    -5.139921e-21, -2.569961e-20, -2.569961e-20, -5.139921e-21, 0, 
    5.139921e-21, 2.569961e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, -5.139921e-21, 3.083953e-20, 1.027984e-20, 
    2.006177e-36, -1.027984e-20, 1.541976e-20, -5.139921e-21, 3.597945e-20, 
    1.541976e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    2.055969e-20, -1.541976e-20, -1.027984e-20, -2.006177e-36, -2.569961e-20, 
    0, -5.139921e-21, -3.083953e-20, -1.027984e-20, -2.006177e-36, 0, 
    -2.569961e-20, 2.006177e-36, 1.541976e-20, -2.006177e-36, -3.083953e-20, 
    5.139921e-21, -3.083953e-20, 5.139921e-21, 3.083953e-20, 5.139921e-21, 
    3.083953e-20, 2.006177e-36, 5.139921e-21, 2.569961e-20, 5.139921e-21, 0, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    -2.006177e-36, 2.055969e-20, 5.139921e-21, 1.027984e-20, 2.006177e-36, 
    2.055969e-20, -5.139921e-21, 2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -2.569961e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 3.597945e-20, 
    2.055969e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, 2.569961e-20, 
    4.111937e-20, 4.625929e-20, -3.597945e-20, -2.055969e-20, 1.027984e-20, 
    -2.055969e-20, -2.055969e-20, 3.597945e-20, -3.083953e-20, 0, 
    -1.027984e-20, -2.006177e-36, 0, -3.597945e-20, 0,
  1.541976e-20, -5.139921e-21, 2.569961e-20, -5.139921e-21, 2.055969e-20, 
    -1.027984e-20, -2.055969e-20, 2.569961e-20, -1.541976e-20, -2.569961e-20, 
    1.027984e-20, -1.541976e-20, -1.027984e-20, 1.027984e-20, 0, 
    -1.027984e-20, -1.027984e-20, -2.006177e-36, 1.541976e-20, 0, 
    -1.541976e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -1.027984e-20, 2.055969e-20, -1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 3.083953e-20, -3.083953e-20, 0, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, -2.006177e-36, 2.055969e-20, 
    5.139921e-21, -1.027984e-20, 2.006177e-36, 5.139921e-21, 1.541976e-20, 
    -2.055969e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, -1.027984e-20, 
    2.055969e-20, -2.006177e-36, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    0, -1.027984e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, -3.597945e-20, 
    -2.055969e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, -2.569961e-20, 
    -2.055969e-20, 5.139921e-21, 0, -1.027984e-20, 0, -2.569961e-20, 
    1.027984e-20, 3.597945e-20, 1.541976e-20, -2.055969e-20, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, 
    3.083953e-20, 1.027984e-20, -2.569961e-20, 2.569961e-20, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, -2.055969e-20, 3.083953e-20, -1.027984e-20, 
    -2.569961e-20, -1.027984e-20, -2.055969e-20, 1.541976e-20, 0, 
    1.027984e-20, -1.541976e-20, 1.027984e-20, -5.139921e-21, 3.083953e-20, 
    5.139921e-21, -2.569961e-20, -2.569961e-20, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -2.006177e-36, 2.006177e-36, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 1.541976e-20, 2.055969e-20, -1.027984e-20, 3.083953e-20, 
    0, 5.139921e-21, 0, 5.139921e-21, -2.569961e-20, -1.541976e-20, 
    -1.027984e-20, -2.569961e-20, 2.055969e-20, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, -2.569961e-20, -2.055969e-20, -1.027984e-20, 1.541976e-20, 
    2.006177e-36, -2.569961e-20, -2.569961e-20, 1.541976e-20, -1.541976e-20, 
    2.055969e-20, 2.055969e-20, -2.055969e-20, -2.055969e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, -2.006177e-36, 2.055969e-20, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, 2.055969e-20, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, -3.083953e-20, 0, -2.569961e-20, 
    2.055969e-20, 5.139921e-21, -2.569961e-20, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 2.006177e-36, 1.027984e-20, 
    1.027984e-20, 3.597945e-20, 2.006177e-36, 4.111937e-20, -1.541976e-20, 
    -1.027984e-20, 1.541976e-20, 0, -2.055969e-20, 2.055969e-20, 0, 
    5.139921e-21, -2.006177e-36, 1.027984e-20, -2.055969e-20, -3.597945e-20, 
    1.027984e-20, -1.541976e-20, 4.111937e-20, -2.006177e-36, 2.055969e-20, 
    -4.111937e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, 0, 
    -2.055969e-20, -4.111937e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 3.597945e-20, 1.541976e-20, -1.541976e-20, 4.625929e-20, 
    5.139921e-21, 5.139921e-21, -2.055969e-20, 2.055969e-20, 3.083953e-20, 0, 
    1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 2.055969e-20, 
    2.055969e-20, 2.055969e-20, -1.541976e-20, 3.597945e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 4.625929e-20, -1.027984e-20, 0, 
    5.139921e-21, -2.055969e-20, -3.083953e-20, -1.027984e-20, 1.027984e-20, 
    2.055969e-20, 1.541976e-20, -2.569961e-20, -2.055969e-20, 3.597945e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    5.139921e-20, 5.139921e-21, 2.569961e-20, -1.541976e-20, 0, 0, 
    2.055969e-20, -1.541976e-20, -2.569961e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, 
    5.139921e-21, 3.597945e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 0, 1.027984e-20, -1.541976e-20, -2.055969e-20, 
    2.006177e-36, -2.055969e-20, -5.139921e-21, -2.055969e-20, 0, 
    3.083953e-20, -1.027984e-20, -1.027984e-20, -3.083953e-20, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 2.569961e-20, 2.569961e-20, 
    -1.541976e-20, 3.083953e-20, -3.083953e-20, 1.027984e-20, 1.541976e-20, 
    -2.055969e-20, 1.541976e-20, 2.006177e-36, -1.027984e-20, -1.027984e-20, 
    -1.541976e-20, -3.083953e-20, -3.083953e-20, -1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 
    2.055969e-20, -2.569961e-20, -5.139921e-21, -1.541976e-20, -2.569961e-20, 
    2.055969e-20, -5.139921e-21, 0, 1.541976e-20, 5.139921e-21, 1.541976e-20, 
    -1.027984e-20, 0, 2.006177e-36,
  8.598827e-29, 8.598799e-29, 8.598804e-29, 8.598782e-29, 8.598795e-29, 
    8.598779e-29, 8.598821e-29, 8.598798e-29, 8.598813e-29, 8.598825e-29, 
    8.598738e-29, 8.598781e-29, 8.598694e-29, 8.598721e-29, 8.598652e-29, 
    8.598698e-29, 8.598643e-29, 8.598654e-29, 8.598622e-29, 8.598631e-29, 
    8.59859e-29, 8.598618e-29, 8.59857e-29, 8.598597e-29, 8.598593e-29, 
    8.598619e-29, 8.598772e-29, 8.598743e-29, 8.598774e-29, 8.59877e-29, 
    8.598772e-29, 8.598794e-29, 8.598805e-29, 8.598829e-29, 8.598825e-29, 
    8.598807e-29, 8.598768e-29, 8.598781e-29, 8.598748e-29, 8.598749e-29, 
    8.598711e-29, 8.598728e-29, 8.598665e-29, 8.598683e-29, 8.598631e-29, 
    8.598644e-29, 8.598631e-29, 8.598635e-29, 8.598631e-29, 8.598651e-29, 
    8.598642e-29, 8.598659e-29, 8.598725e-29, 8.598705e-29, 8.598763e-29, 
    8.598798e-29, 8.59882e-29, 8.598837e-29, 8.598834e-29, 8.59883e-29, 
    8.598807e-29, 8.598786e-29, 8.59877e-29, 8.598759e-29, 8.598749e-29, 
    8.598716e-29, 8.598699e-29, 8.598661e-29, 8.598668e-29, 8.598656e-29, 
    8.598645e-29, 8.598627e-29, 8.59863e-29, 8.598621e-29, 8.598657e-29, 
    8.598633e-29, 8.598672e-29, 8.598662e-29, 8.598746e-29, 8.598778e-29, 
    8.598792e-29, 8.598804e-29, 8.598832e-29, 8.598813e-29, 8.59882e-29, 
    8.598802e-29, 8.59879e-29, 8.598796e-29, 8.598759e-29, 8.598773e-29, 
    8.598698e-29, 8.598731e-29, 8.598646e-29, 8.598667e-29, 8.598642e-29, 
    8.598654e-29, 8.598633e-29, 8.598652e-29, 8.598618e-29, 8.598611e-29, 
    8.598616e-29, 8.598597e-29, 8.598653e-29, 8.598631e-29, 8.598796e-29, 
    8.598795e-29, 8.59879e-29, 8.59881e-29, 8.598811e-29, 8.598829e-29, 
    8.598813e-29, 8.598806e-29, 8.598789e-29, 8.598778e-29, 8.598769e-29, 
    8.598747e-29, 8.598723e-29, 8.59869e-29, 8.598665e-29, 8.598649e-29, 
    8.598659e-29, 8.59865e-29, 8.59866e-29, 8.598665e-29, 8.598613e-29, 
    8.598642e-29, 8.598599e-29, 8.598601e-29, 8.598621e-29, 8.598601e-29, 
    8.598794e-29, 8.598799e-29, 8.598819e-29, 8.598804e-29, 8.598831e-29, 
    8.598816e-29, 8.598807e-29, 8.598773e-29, 8.598766e-29, 8.598758e-29, 
    8.598745e-29, 8.598727e-29, 8.598696e-29, 8.598669e-29, 8.598645e-29, 
    8.598646e-29, 8.598646e-29, 8.59864e-29, 8.598654e-29, 8.598638e-29, 
    8.598636e-29, 8.598642e-29, 8.598602e-29, 8.598613e-29, 8.598601e-29, 
    8.598609e-29, 8.598798e-29, 8.598788e-29, 8.598793e-29, 8.598784e-29, 
    8.598791e-29, 8.598761e-29, 8.598752e-29, 8.59871e-29, 8.598727e-29, 
    8.5987e-29, 8.598725e-29, 8.59872e-29, 8.598699e-29, 8.598723e-29, 
    8.598671e-29, 8.598707e-29, 8.59864e-29, 8.598676e-29, 8.598638e-29, 
    8.598645e-29, 8.598633e-29, 8.598623e-29, 8.59861e-29, 8.598586e-29, 
    8.598592e-29, 8.598572e-29, 8.598775e-29, 8.598763e-29, 8.598763e-29, 
    8.598751e-29, 8.598742e-29, 8.598721e-29, 8.598689e-29, 8.598701e-29, 
    8.598678e-29, 8.598674e-29, 8.598708e-29, 8.598687e-29, 8.598754e-29, 
    8.598743e-29, 8.59875e-29, 8.598773e-29, 8.598698e-29, 8.598737e-29, 
    8.598665e-29, 8.598686e-29, 8.598625e-29, 8.598655e-29, 8.598595e-29, 
    8.598569e-29, 8.598545e-29, 8.598516e-29, 8.598756e-29, 8.598764e-29, 
    8.598749e-29, 8.598729e-29, 8.59871e-29, 8.598685e-29, 8.598682e-29, 
    8.598677e-29, 8.598665e-29, 8.598655e-29, 8.598676e-29, 8.598652e-29, 
    8.598741e-29, 8.598695e-29, 8.598767e-29, 8.598745e-29, 8.59873e-29, 
    8.598737e-29, 8.598702e-29, 8.598694e-29, 8.598661e-29, 8.598678e-29, 
    8.598575e-29, 8.598621e-29, 8.598495e-29, 8.59853e-29, 8.598767e-29, 
    8.598756e-29, 8.598717e-29, 8.598736e-29, 8.598683e-29, 8.59867e-29, 
    8.59866e-29, 8.598646e-29, 8.598645e-29, 8.598637e-29, 8.598649e-29, 
    8.598637e-29, 8.598684e-29, 8.598663e-29, 8.598722e-29, 8.598707e-29, 
    8.598714e-29, 8.598721e-29, 8.598699e-29, 8.598675e-29, 8.598675e-29, 
    8.598668e-29, 8.598646e-29, 8.598683e-29, 8.59857e-29, 8.59864e-29, 
    8.598744e-29, 8.598722e-29, 8.598719e-29, 8.598728e-29, 8.598671e-29, 
    8.598692e-29, 8.598637e-29, 8.598652e-29, 8.598627e-29, 8.598639e-29, 
    8.598641e-29, 8.598657e-29, 8.598666e-29, 8.598691e-29, 8.598711e-29, 
    8.598727e-29, 8.598723e-29, 8.598705e-29, 8.598674e-29, 8.598645e-29, 
    8.598651e-29, 8.598629e-29, 8.598687e-29, 8.598663e-29, 8.598672e-29, 
    8.598648e-29, 8.598701e-29, 8.598655e-29, 8.598713e-29, 8.598708e-29, 
    8.598692e-29, 8.598661e-29, 8.598654e-29, 8.598647e-29, 8.598651e-29, 
    8.598674e-29, 8.598677e-29, 8.598693e-29, 8.598697e-29, 8.598708e-29, 
    8.598719e-29, 8.59871e-29, 8.5987e-29, 8.598674e-29, 8.598649e-29, 
    8.598623e-29, 8.598616e-29, 8.598586e-29, 8.598611e-29, 8.598569e-29, 
    8.598604e-29, 8.598544e-29, 8.598653e-29, 8.598606e-29, 8.598692e-29, 
    8.598682e-29, 8.598666e-29, 8.598627e-29, 8.598648e-29, 8.598624e-29, 
    8.598677e-29, 8.598705e-29, 8.598712e-29, 8.598725e-29, 8.598711e-29, 
    8.598713e-29, 8.5987e-29, 8.598704e-29, 8.598672e-29, 8.598689e-29, 
    8.598641e-29, 8.598624e-29, 8.598574e-29, 8.598544e-29, 8.598513e-29, 
    8.598499e-29, 8.598495e-29, 8.598493e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.134403e-08, 1.139405e-08, 1.138433e-08, 1.142467e-08, 1.140229e-08, 
    1.142871e-08, 1.135418e-08, 1.139604e-08, 1.136931e-08, 1.134854e-08, 
    1.150296e-08, 1.142647e-08, 1.158243e-08, 1.153364e-08, 1.165621e-08, 
    1.157484e-08, 1.167262e-08, 1.165387e-08, 1.171032e-08, 1.169415e-08, 
    1.176635e-08, 1.171779e-08, 1.180379e-08, 1.175476e-08, 1.176242e-08, 
    1.171618e-08, 1.144187e-08, 1.149344e-08, 1.143881e-08, 1.144616e-08, 
    1.144286e-08, 1.140275e-08, 1.138254e-08, 1.134021e-08, 1.13479e-08, 
    1.137899e-08, 1.144947e-08, 1.142554e-08, 1.148585e-08, 1.148449e-08, 
    1.155162e-08, 1.152135e-08, 1.163421e-08, 1.160213e-08, 1.169482e-08, 
    1.167151e-08, 1.169373e-08, 1.168699e-08, 1.169381e-08, 1.165963e-08, 
    1.167427e-08, 1.164419e-08, 1.152702e-08, 1.156145e-08, 1.145876e-08, 
    1.139701e-08, 1.135601e-08, 1.132691e-08, 1.133103e-08, 1.133887e-08, 
    1.137917e-08, 1.141706e-08, 1.144594e-08, 1.146526e-08, 1.148429e-08, 
    1.15419e-08, 1.15724e-08, 1.164069e-08, 1.162837e-08, 1.164924e-08, 
    1.166919e-08, 1.170268e-08, 1.169717e-08, 1.171192e-08, 1.16487e-08, 
    1.169071e-08, 1.162135e-08, 1.164032e-08, 1.148946e-08, 1.1432e-08, 
    1.140757e-08, 1.13862e-08, 1.133419e-08, 1.13701e-08, 1.135595e-08, 
    1.138963e-08, 1.141103e-08, 1.140045e-08, 1.146578e-08, 1.144038e-08, 
    1.157421e-08, 1.151656e-08, 1.166686e-08, 1.16309e-08, 1.167549e-08, 
    1.165273e-08, 1.169172e-08, 1.165663e-08, 1.171741e-08, 1.173065e-08, 
    1.17216e-08, 1.175635e-08, 1.165469e-08, 1.169373e-08, 1.140015e-08, 
    1.140188e-08, 1.140992e-08, 1.137456e-08, 1.13724e-08, 1.134e-08, 
    1.136883e-08, 1.138111e-08, 1.141228e-08, 1.143071e-08, 1.144824e-08, 
    1.148677e-08, 1.15298e-08, 1.158999e-08, 1.163323e-08, 1.166221e-08, 
    1.164444e-08, 1.166013e-08, 1.164259e-08, 1.163437e-08, 1.172569e-08, 
    1.167441e-08, 1.175135e-08, 1.174709e-08, 1.171227e-08, 1.174757e-08, 
    1.140309e-08, 1.139316e-08, 1.135866e-08, 1.138566e-08, 1.133647e-08, 
    1.1364e-08, 1.137983e-08, 1.144091e-08, 1.145434e-08, 1.146678e-08, 
    1.149136e-08, 1.15229e-08, 1.157824e-08, 1.162639e-08, 1.167035e-08, 
    1.166713e-08, 1.166827e-08, 1.167809e-08, 1.165376e-08, 1.168208e-08, 
    1.168683e-08, 1.16744e-08, 1.174652e-08, 1.172592e-08, 1.1747e-08, 
    1.173359e-08, 1.139639e-08, 1.14131e-08, 1.140407e-08, 1.142106e-08, 
    1.140909e-08, 1.14623e-08, 1.147826e-08, 1.155292e-08, 1.152228e-08, 
    1.157105e-08, 1.152724e-08, 1.1535e-08, 1.157264e-08, 1.15296e-08, 
    1.162373e-08, 1.155991e-08, 1.167847e-08, 1.161473e-08, 1.168246e-08, 
    1.167016e-08, 1.169053e-08, 1.170876e-08, 1.173171e-08, 1.177405e-08, 
    1.176424e-08, 1.179965e-08, 1.143803e-08, 1.145971e-08, 1.14578e-08, 
    1.148049e-08, 1.149728e-08, 1.153366e-08, 1.1592e-08, 1.157006e-08, 
    1.161035e-08, 1.161843e-08, 1.155723e-08, 1.159481e-08, 1.147422e-08, 
    1.14937e-08, 1.148211e-08, 1.143974e-08, 1.157512e-08, 1.150564e-08, 
    1.163394e-08, 1.15963e-08, 1.170616e-08, 1.165152e-08, 1.175885e-08, 
    1.180472e-08, 1.184791e-08, 1.189838e-08, 1.147154e-08, 1.145681e-08, 
    1.148319e-08, 1.151969e-08, 1.155357e-08, 1.15986e-08, 1.16032e-08, 
    1.161164e-08, 1.163349e-08, 1.165187e-08, 1.161431e-08, 1.165647e-08, 
    1.149822e-08, 1.158115e-08, 1.145124e-08, 1.149035e-08, 1.151754e-08, 
    1.150562e-08, 1.156756e-08, 1.158215e-08, 1.164148e-08, 1.161081e-08, 
    1.17934e-08, 1.171261e-08, 1.193681e-08, 1.187415e-08, 1.145166e-08, 
    1.147149e-08, 1.154052e-08, 1.150768e-08, 1.16016e-08, 1.162472e-08, 
    1.164352e-08, 1.166755e-08, 1.167014e-08, 1.168438e-08, 1.166105e-08, 
    1.168346e-08, 1.159869e-08, 1.163657e-08, 1.153263e-08, 1.155793e-08, 
    1.154629e-08, 1.153352e-08, 1.157292e-08, 1.16149e-08, 1.16158e-08, 
    1.162925e-08, 1.166718e-08, 1.160198e-08, 1.180382e-08, 1.167916e-08, 
    1.149312e-08, 1.153132e-08, 1.153678e-08, 1.152198e-08, 1.162241e-08, 
    1.158602e-08, 1.168403e-08, 1.165754e-08, 1.170095e-08, 1.167938e-08, 
    1.16762e-08, 1.16485e-08, 1.163126e-08, 1.158768e-08, 1.155223e-08, 
    1.152413e-08, 1.153066e-08, 1.156154e-08, 1.161746e-08, 1.167038e-08, 
    1.165879e-08, 1.169765e-08, 1.159479e-08, 1.163792e-08, 1.162125e-08, 
    1.166472e-08, 1.156948e-08, 1.165057e-08, 1.154875e-08, 1.155768e-08, 
    1.158529e-08, 1.164084e-08, 1.165314e-08, 1.166626e-08, 1.165816e-08, 
    1.161889e-08, 1.161245e-08, 1.158462e-08, 1.157694e-08, 1.155574e-08, 
    1.153818e-08, 1.155422e-08, 1.157106e-08, 1.16189e-08, 1.166202e-08, 
    1.170902e-08, 1.172053e-08, 1.177545e-08, 1.173074e-08, 1.180451e-08, 
    1.174178e-08, 1.185038e-08, 1.165527e-08, 1.173994e-08, 1.158655e-08, 
    1.160308e-08, 1.163296e-08, 1.170152e-08, 1.166451e-08, 1.170779e-08, 
    1.16122e-08, 1.15626e-08, 1.154977e-08, 1.152584e-08, 1.155032e-08, 
    1.154833e-08, 1.157176e-08, 1.156423e-08, 1.162049e-08, 1.159027e-08, 
    1.167612e-08, 1.170745e-08, 1.179594e-08, 1.185019e-08, 1.190541e-08, 
    1.192979e-08, 1.193721e-08, 1.194032e-08 ;

 SOIL1N_TO_SOIL3N =
  1.346024e-10, 1.351961e-10, 1.350807e-10, 1.355595e-10, 1.352939e-10, 
    1.356074e-10, 1.347227e-10, 1.352196e-10, 1.349024e-10, 1.346558e-10, 
    1.364888e-10, 1.355809e-10, 1.374322e-10, 1.36853e-10, 1.38308e-10, 
    1.373421e-10, 1.385028e-10, 1.382802e-10, 1.389503e-10, 1.387583e-10, 
    1.396154e-10, 1.390389e-10, 1.400598e-10, 1.394778e-10, 1.395688e-10, 
    1.390199e-10, 1.357636e-10, 1.363758e-10, 1.357274e-10, 1.358147e-10, 
    1.357755e-10, 1.352994e-10, 1.350594e-10, 1.34557e-10, 1.346482e-10, 
    1.350172e-10, 1.358539e-10, 1.355699e-10, 1.362857e-10, 1.362696e-10, 
    1.370665e-10, 1.367072e-10, 1.380468e-10, 1.37666e-10, 1.387663e-10, 
    1.384896e-10, 1.387533e-10, 1.386734e-10, 1.387544e-10, 1.383485e-10, 
    1.385224e-10, 1.381653e-10, 1.367745e-10, 1.371832e-10, 1.359642e-10, 
    1.352313e-10, 1.347445e-10, 1.343991e-10, 1.34448e-10, 1.34541e-10, 
    1.350194e-10, 1.354692e-10, 1.35812e-10, 1.360413e-10, 1.362672e-10, 
    1.369511e-10, 1.373131e-10, 1.381237e-10, 1.379775e-10, 1.382253e-10, 
    1.384621e-10, 1.388596e-10, 1.387942e-10, 1.389693e-10, 1.382188e-10, 
    1.387176e-10, 1.378942e-10, 1.381193e-10, 1.363285e-10, 1.356465e-10, 
    1.353566e-10, 1.351028e-10, 1.344855e-10, 1.349118e-10, 1.347438e-10, 
    1.351436e-10, 1.353977e-10, 1.35272e-10, 1.360476e-10, 1.35746e-10, 
    1.373346e-10, 1.366503e-10, 1.384345e-10, 1.380075e-10, 1.385368e-10, 
    1.382667e-10, 1.387295e-10, 1.38313e-10, 1.390345e-10, 1.391916e-10, 
    1.390842e-10, 1.394967e-10, 1.382899e-10, 1.387533e-10, 1.352685e-10, 
    1.35289e-10, 1.353845e-10, 1.349648e-10, 1.349391e-10, 1.345545e-10, 
    1.348967e-10, 1.350424e-10, 1.354124e-10, 1.356312e-10, 1.358392e-10, 
    1.362966e-10, 1.368075e-10, 1.375219e-10, 1.380352e-10, 1.383793e-10, 
    1.381683e-10, 1.383545e-10, 1.381463e-10, 1.380487e-10, 1.391327e-10, 
    1.38524e-10, 1.394374e-10, 1.393868e-10, 1.389735e-10, 1.393925e-10, 
    1.353034e-10, 1.351854e-10, 1.34776e-10, 1.350964e-10, 1.345126e-10, 
    1.348394e-10, 1.350273e-10, 1.357523e-10, 1.359116e-10, 1.360594e-10, 
    1.363511e-10, 1.367255e-10, 1.373824e-10, 1.37954e-10, 1.384759e-10, 
    1.384376e-10, 1.384511e-10, 1.385676e-10, 1.382789e-10, 1.38615e-10, 
    1.386715e-10, 1.38524e-10, 1.3938e-10, 1.391355e-10, 1.393858e-10, 
    1.392265e-10, 1.352238e-10, 1.354222e-10, 1.35315e-10, 1.355166e-10, 
    1.353746e-10, 1.360062e-10, 1.361956e-10, 1.370819e-10, 1.367182e-10, 
    1.372971e-10, 1.36777e-10, 1.368691e-10, 1.373159e-10, 1.368051e-10, 
    1.379225e-10, 1.371649e-10, 1.385722e-10, 1.378155e-10, 1.386196e-10, 
    1.384736e-10, 1.387153e-10, 1.389318e-10, 1.392042e-10, 1.397068e-10, 
    1.395904e-10, 1.400107e-10, 1.35718e-10, 1.359754e-10, 1.359528e-10, 
    1.362222e-10, 1.364214e-10, 1.368532e-10, 1.375458e-10, 1.372854e-10, 
    1.377635e-10, 1.378595e-10, 1.371331e-10, 1.375791e-10, 1.361477e-10, 
    1.363789e-10, 1.362413e-10, 1.357384e-10, 1.373454e-10, 1.365206e-10, 
    1.380436e-10, 1.375968e-10, 1.389009e-10, 1.382523e-10, 1.395263e-10, 
    1.40071e-10, 1.405837e-10, 1.411827e-10, 1.361159e-10, 1.35941e-10, 
    1.362542e-10, 1.366875e-10, 1.370895e-10, 1.376241e-10, 1.376788e-10, 
    1.377789e-10, 1.380383e-10, 1.382564e-10, 1.378105e-10, 1.383111e-10, 
    1.364325e-10, 1.37417e-10, 1.358749e-10, 1.363392e-10, 1.366619e-10, 
    1.365204e-10, 1.372556e-10, 1.374289e-10, 1.381331e-10, 1.377691e-10, 
    1.399365e-10, 1.389775e-10, 1.41639e-10, 1.408951e-10, 1.358799e-10, 
    1.361153e-10, 1.369346e-10, 1.365448e-10, 1.376598e-10, 1.379342e-10, 
    1.381573e-10, 1.384425e-10, 1.384734e-10, 1.386423e-10, 1.383654e-10, 
    1.386314e-10, 1.376252e-10, 1.380748e-10, 1.36841e-10, 1.371413e-10, 
    1.370032e-10, 1.368516e-10, 1.373193e-10, 1.378175e-10, 1.378282e-10, 
    1.37988e-10, 1.384382e-10, 1.376643e-10, 1.400602e-10, 1.385804e-10, 
    1.36372e-10, 1.368255e-10, 1.368902e-10, 1.367146e-10, 1.379067e-10, 
    1.374747e-10, 1.386382e-10, 1.383238e-10, 1.38839e-10, 1.38583e-10, 
    1.385453e-10, 1.382165e-10, 1.380117e-10, 1.374945e-10, 1.370737e-10, 
    1.367401e-10, 1.368177e-10, 1.371842e-10, 1.37848e-10, 1.384761e-10, 
    1.383385e-10, 1.387999e-10, 1.375789e-10, 1.380908e-10, 1.37893e-10, 
    1.384089e-10, 1.372784e-10, 1.38241e-10, 1.370324e-10, 1.371384e-10, 
    1.374662e-10, 1.381255e-10, 1.382715e-10, 1.384272e-10, 1.383311e-10, 
    1.378649e-10, 1.377885e-10, 1.374582e-10, 1.37367e-10, 1.371153e-10, 
    1.369069e-10, 1.370973e-10, 1.372972e-10, 1.378651e-10, 1.383769e-10, 
    1.389349e-10, 1.390715e-10, 1.397234e-10, 1.391927e-10, 1.400685e-10, 
    1.393238e-10, 1.40613e-10, 1.382968e-10, 1.39302e-10, 1.374811e-10, 
    1.376772e-10, 1.38032e-10, 1.388458e-10, 1.384065e-10, 1.389203e-10, 
    1.377855e-10, 1.371968e-10, 1.370445e-10, 1.367604e-10, 1.37051e-10, 
    1.370274e-10, 1.373055e-10, 1.372162e-10, 1.37884e-10, 1.375252e-10, 
    1.385444e-10, 1.389163e-10, 1.399667e-10, 1.406106e-10, 1.412662e-10, 
    1.415557e-10, 1.416438e-10, 1.416806e-10 ;

 SOIL1N_vr =
  2.497656, 2.497649, 2.49765, 2.497645, 2.497648, 2.497645, 2.497654, 
    2.497649, 2.497652, 2.497655, 2.497635, 2.497645, 2.497625, 2.497631, 
    2.497615, 2.497626, 2.497613, 2.497616, 2.497608, 2.497611, 2.497601, 
    2.497607, 2.497597, 2.497603, 2.497602, 2.497608, 2.497643, 2.497636, 
    2.497643, 2.497643, 2.497643, 2.497648, 2.497651, 2.497656, 2.497655, 
    2.497651, 2.497642, 2.497645, 2.497637, 2.497638, 2.497629, 2.497633, 
    2.497618, 2.497622, 2.497611, 2.497613, 2.497611, 2.497612, 2.497611, 
    2.497615, 2.497613, 2.497617, 2.497632, 2.497627, 2.497641, 2.497649, 
    2.497654, 2.497658, 2.497657, 2.497656, 2.497651, 2.497646, 2.497643, 
    2.49764, 2.497638, 2.49763, 2.497626, 2.497617, 2.497619, 2.497616, 
    2.497614, 2.497609, 2.49761, 2.497608, 2.497616, 2.497611, 2.49762, 
    2.497617, 2.497637, 2.497644, 2.497648, 2.49765, 2.497657, 2.497652, 
    2.497654, 2.49765, 2.497647, 2.497648, 2.49764, 2.497643, 2.497626, 
    2.497633, 2.497614, 2.497619, 2.497613, 2.497616, 2.497611, 2.497615, 
    2.497607, 2.497606, 2.497607, 2.497602, 2.497616, 2.497611, 2.497648, 
    2.497648, 2.497647, 2.497652, 2.497652, 2.497656, 2.497653, 2.497651, 
    2.497647, 2.497644, 2.497642, 2.497637, 2.497632, 2.497624, 2.497618, 
    2.497615, 2.497617, 2.497615, 2.497617, 2.497618, 2.497607, 2.497613, 
    2.497603, 2.497604, 2.497608, 2.497604, 2.497648, 2.497649, 2.497654, 
    2.49765, 2.497657, 2.497653, 2.497651, 2.497643, 2.497641, 2.49764, 
    2.497637, 2.497633, 2.497625, 2.497619, 2.497614, 2.497614, 2.497614, 
    2.497613, 2.497616, 2.497612, 2.497612, 2.497613, 2.497604, 2.497607, 
    2.497604, 2.497606, 2.497649, 2.497647, 2.497648, 2.497646, 2.497647, 
    2.49764, 2.497638, 2.497629, 2.497633, 2.497626, 2.497632, 2.497631, 
    2.497626, 2.497632, 2.49762, 2.497628, 2.497612, 2.497621, 2.497612, 
    2.497614, 2.497611, 2.497609, 2.497606, 2.4976, 2.497602, 2.497597, 
    2.497643, 2.497641, 2.497641, 2.497638, 2.497636, 2.497631, 2.497624, 
    2.497627, 2.497621, 2.49762, 2.497628, 2.497623, 2.497639, 2.497636, 
    2.497638, 2.497643, 2.497626, 2.497635, 2.497618, 2.497623, 2.497609, 
    2.497616, 2.497602, 2.497596, 2.497591, 2.497584, 2.497639, 2.497641, 
    2.497638, 2.497633, 2.497629, 2.497623, 2.497622, 2.497621, 2.497618, 
    2.497616, 2.497621, 2.497615, 2.497636, 2.497625, 2.497642, 2.497637, 
    2.497633, 2.497635, 2.497627, 2.497625, 2.497617, 2.497621, 2.497598, 
    2.497608, 2.497579, 2.497587, 2.497642, 2.497639, 2.49763, 2.497635, 
    2.497622, 2.497619, 2.497617, 2.497614, 2.497614, 2.497612, 2.497615, 
    2.497612, 2.497623, 2.497618, 2.497631, 2.497628, 2.49763, 2.497631, 
    2.497626, 2.497621, 2.497621, 2.497619, 2.497614, 2.497622, 2.497597, 
    2.497612, 2.497636, 2.497632, 2.497631, 2.497633, 2.49762, 2.497624, 
    2.497612, 2.497615, 2.49761, 2.497612, 2.497613, 2.497617, 2.497619, 
    2.497624, 2.497629, 2.497633, 2.497632, 2.497627, 2.49762, 2.497614, 
    2.497615, 2.49761, 2.497623, 2.497618, 2.49762, 2.497614, 2.497627, 
    2.497616, 2.497629, 2.497628, 2.497625, 2.497617, 2.497616, 2.497614, 
    2.497615, 2.49762, 2.497621, 2.497625, 2.497626, 2.497628, 2.497631, 
    2.497628, 2.497626, 2.49762, 2.497615, 2.497609, 2.497607, 2.4976, 
    2.497606, 2.497597, 2.497604, 2.497591, 2.497616, 2.497605, 2.497624, 
    2.497622, 2.497618, 2.49761, 2.497614, 2.497609, 2.497621, 2.497627, 
    2.497629, 2.497632, 2.497629, 2.497629, 2.497626, 2.497627, 2.49762, 
    2.497624, 2.497613, 2.497609, 2.497597, 2.497591, 2.497583, 2.49758, 
    2.497579, 2.497579,
  2.497912, 2.497904, 2.497906, 2.4979, 2.497903, 2.497899, 2.497911, 
    2.497904, 2.497908, 2.497911, 2.497887, 2.497899, 2.497874, 2.497882, 
    2.497863, 2.497876, 2.49786, 2.497863, 2.497854, 2.497857, 2.497846, 
    2.497853, 2.49784, 2.497847, 2.497846, 2.497854, 2.497897, 2.497889, 
    2.497897, 2.497896, 2.497897, 2.497903, 2.497906, 2.497913, 2.497912, 
    2.497907, 2.497895, 2.497899, 2.49789, 2.49789, 2.497879, 2.497884, 
    2.497866, 2.497871, 2.497857, 2.49786, 2.497857, 2.497858, 2.497857, 
    2.497862, 2.49786, 2.497865, 2.497883, 2.497878, 2.497894, 2.497904, 
    2.49791, 2.497915, 2.497914, 2.497913, 2.497907, 2.497901, 2.497896, 
    2.497893, 2.49789, 2.497881, 2.497876, 2.497865, 2.497867, 2.497864, 
    2.497861, 2.497856, 2.497856, 2.497854, 2.497864, 2.497857, 2.497868, 
    2.497865, 2.497889, 2.497898, 2.497902, 2.497905, 2.497914, 2.497908, 
    2.49791, 2.497905, 2.497902, 2.497903, 2.497893, 2.497897, 2.497876, 
    2.497885, 2.497861, 2.497867, 2.49786, 2.497864, 2.497857, 2.497863, 
    2.497853, 2.497851, 2.497853, 2.497847, 2.497863, 2.497857, 2.497903, 
    2.497903, 2.497902, 2.497907, 2.497908, 2.497913, 2.497908, 2.497906, 
    2.497901, 2.497899, 2.497896, 2.49789, 2.497883, 2.497873, 2.497866, 
    2.497862, 2.497865, 2.497862, 2.497865, 2.497866, 2.497852, 2.49786, 
    2.497848, 2.497849, 2.497854, 2.497849, 2.497903, 2.497905, 2.49791, 
    2.497906, 2.497913, 2.497909, 2.497906, 2.497897, 2.497895, 2.497893, 
    2.497889, 2.497884, 2.497875, 2.497868, 2.497861, 2.497861, 2.497861, 
    2.497859, 2.497863, 2.497859, 2.497858, 2.49786, 2.497849, 2.497852, 
    2.497849, 2.497851, 2.497904, 2.497901, 2.497903, 2.4979, 2.497902, 
    2.497894, 2.497891, 2.497879, 2.497884, 2.497876, 2.497883, 2.497882, 
    2.497876, 2.497883, 2.497868, 2.497878, 2.497859, 2.497869, 2.497859, 
    2.497861, 2.497858, 2.497855, 2.497851, 2.497844, 2.497846, 2.49784, 
    2.497897, 2.497894, 2.497894, 2.497891, 2.497888, 2.497882, 2.497873, 
    2.497876, 2.49787, 2.497869, 2.497879, 2.497873, 2.497892, 2.497889, 
    2.49789, 2.497897, 2.497876, 2.497887, 2.497866, 2.497872, 2.497855, 
    2.497864, 2.497847, 2.497839, 2.497833, 2.497825, 2.497892, 2.497894, 
    2.49789, 2.497885, 2.497879, 2.497872, 2.497871, 2.49787, 2.497866, 
    2.497864, 2.497869, 2.497863, 2.497888, 2.497875, 2.497895, 2.497889, 
    2.497885, 2.497887, 2.497877, 2.497874, 2.497865, 2.49787, 2.497841, 
    2.497854, 2.497819, 2.497829, 2.497895, 2.497892, 2.497881, 2.497886, 
    2.497871, 2.497868, 2.497865, 2.497861, 2.497861, 2.497859, 2.497862, 
    2.497859, 2.497872, 2.497866, 2.497882, 2.497878, 2.49788, 2.497882, 
    2.497876, 2.497869, 2.497869, 2.497867, 2.497861, 2.497871, 2.49784, 
    2.497859, 2.497889, 2.497883, 2.497882, 2.497884, 2.497868, 2.497874, 
    2.497859, 2.497863, 2.497856, 2.497859, 2.49786, 2.497864, 2.497867, 
    2.497874, 2.497879, 2.497884, 2.497883, 2.497878, 2.497869, 2.497861, 
    2.497863, 2.497856, 2.497873, 2.497866, 2.497868, 2.497862, 2.497877, 
    2.497864, 2.49788, 2.497878, 2.497874, 2.497865, 2.497863, 2.497861, 
    2.497863, 2.497869, 2.49787, 2.497874, 2.497875, 2.497879, 2.497881, 
    2.497879, 2.497876, 2.497869, 2.497862, 2.497854, 2.497853, 2.497844, 
    2.497851, 2.497839, 2.497849, 2.497832, 2.497863, 2.49785, 2.497874, 
    2.497871, 2.497867, 2.497856, 2.497862, 2.497855, 2.49787, 2.497878, 
    2.49788, 2.497884, 2.49788, 2.49788, 2.497876, 2.497877, 2.497869, 
    2.497873, 2.49786, 2.497855, 2.497841, 2.497832, 2.497824, 2.49782, 
    2.497819, 2.497818,
  2.498032, 2.498024, 2.498025, 2.498018, 2.498022, 2.498017, 2.49803, 
    2.498023, 2.498028, 2.498031, 2.498004, 2.498018, 2.497991, 2.497999, 
    2.497978, 2.497992, 2.497975, 2.497978, 2.497968, 2.497971, 2.497959, 
    2.497967, 2.497952, 2.497961, 2.497959, 2.497967, 2.498015, 2.498006, 
    2.498016, 2.498014, 2.498015, 2.498022, 2.498025, 2.498033, 2.498031, 
    2.498026, 2.498014, 2.498018, 2.498008, 2.498008, 2.497996, 2.498001, 
    2.497982, 2.497987, 2.497971, 2.497975, 2.497971, 2.497972, 2.497971, 
    2.497977, 2.497975, 2.49798, 2.498, 2.497994, 2.498012, 2.498023, 
    2.49803, 2.498035, 2.498034, 2.498033, 2.498026, 2.498019, 2.498014, 
    2.498011, 2.498008, 2.497998, 2.497992, 2.497981, 2.497983, 2.497979, 
    2.497976, 2.49797, 2.497971, 2.497968, 2.497979, 2.497972, 2.497984, 
    2.497981, 2.498007, 2.498017, 2.498021, 2.498025, 2.498034, 2.498028, 
    2.49803, 2.498024, 2.49802, 2.498022, 2.498011, 2.498015, 2.497992, 
    2.498002, 2.497976, 2.497982, 2.497974, 2.497978, 2.497972, 2.497978, 
    2.497967, 2.497965, 2.497967, 2.49796, 2.497978, 2.497971, 2.498022, 
    2.498022, 2.498021, 2.498027, 2.498027, 2.498033, 2.498028, 2.498026, 
    2.49802, 2.498017, 2.498014, 2.498007, 2.498, 2.497989, 2.497982, 
    2.497977, 2.49798, 2.497977, 2.49798, 2.497982, 2.497966, 2.497975, 
    2.497961, 2.497962, 2.497968, 2.497962, 2.498022, 2.498024, 2.498029, 
    2.498025, 2.498034, 2.498029, 2.498026, 2.498015, 2.498013, 2.498011, 
    2.498006, 2.498001, 2.497991, 2.497983, 2.497975, 2.497976, 2.497976, 
    2.497974, 2.497978, 2.497973, 2.497972, 2.497975, 2.497962, 2.497966, 
    2.497962, 2.497964, 2.498023, 2.49802, 2.498022, 2.498019, 2.498021, 
    2.498012, 2.498009, 2.497996, 2.498001, 2.497993, 2.498, 2.497999, 
    2.497992, 2.498, 2.497983, 2.497994, 2.497974, 2.497985, 2.497973, 
    2.497975, 2.497972, 2.497969, 2.497965, 2.497957, 2.497959, 2.497953, 
    2.498016, 2.498012, 2.498012, 2.498008, 2.498005, 2.497999, 2.497989, 
    2.497993, 2.497986, 2.497984, 2.497995, 2.497988, 2.498009, 2.498006, 
    2.498008, 2.498015, 2.497992, 2.498004, 2.497982, 2.497988, 2.497969, 
    2.497979, 2.49796, 2.497952, 2.497945, 2.497936, 2.49801, 2.498013, 
    2.498008, 2.498002, 2.497996, 2.497988, 2.497987, 2.497986, 2.497982, 
    2.497978, 2.497985, 2.497978, 2.498005, 2.497991, 2.498013, 2.498007, 
    2.498002, 2.498004, 2.497993, 2.497991, 2.49798, 2.497986, 2.497954, 
    2.497968, 2.497929, 2.49794, 2.498013, 2.49801, 2.497998, 2.498004, 
    2.497987, 2.497983, 2.49798, 2.497976, 2.497975, 2.497973, 2.497977, 
    2.497973, 2.497988, 2.497981, 2.497999, 2.497995, 2.497997, 2.497999, 
    2.497992, 2.497985, 2.497985, 2.497983, 2.497976, 2.497987, 2.497952, 
    2.497974, 2.498006, 2.497999, 2.497998, 2.498001, 2.497984, 2.49799, 
    2.497973, 2.497977, 2.49797, 2.497974, 2.497974, 2.497979, 2.497982, 
    2.49799, 2.497996, 2.498001, 2.498, 2.497994, 2.497984, 2.497975, 
    2.497977, 2.497971, 2.497988, 2.497981, 2.497984, 2.497976, 2.497993, 
    2.497979, 2.497997, 2.497995, 2.49799, 2.49798, 2.497978, 2.497976, 
    2.497977, 2.497984, 2.497985, 2.49799, 2.497992, 2.497995, 2.497998, 
    2.497996, 2.497993, 2.497984, 2.497977, 2.497969, 2.497967, 2.497957, 
    2.497965, 2.497952, 2.497963, 2.497944, 2.497978, 2.497963, 2.49799, 
    2.497987, 2.497982, 2.49797, 2.497976, 2.497969, 2.497985, 2.497994, 
    2.497996, 2.498, 2.497996, 2.497997, 2.497993, 2.497994, 2.497984, 
    2.497989, 2.497974, 2.497969, 2.497954, 2.497944, 2.497935, 2.49793, 
    2.497929, 2.497929,
  2.498126, 2.498117, 2.498119, 2.498111, 2.498116, 2.498111, 2.498124, 
    2.498116, 2.498121, 2.498125, 2.498097, 2.498111, 2.498083, 2.498092, 
    2.49807, 2.498085, 2.498067, 2.498071, 2.498061, 2.498064, 2.498051, 
    2.498059, 2.498044, 2.498053, 2.498051, 2.49806, 2.498108, 2.498099, 
    2.498109, 2.498108, 2.498108, 2.498115, 2.498119, 2.498127, 2.498125, 
    2.49812, 2.498107, 2.498111, 2.498101, 2.498101, 2.498089, 2.498094, 
    2.498074, 2.49808, 2.498063, 2.498068, 2.498064, 2.498065, 2.498064, 
    2.49807, 2.498067, 2.498072, 2.498093, 2.498087, 2.498105, 2.498116, 
    2.498124, 2.498129, 2.498128, 2.498127, 2.49812, 2.498113, 2.498108, 
    2.498104, 2.498101, 2.498091, 2.498085, 2.498073, 2.498075, 2.498071, 
    2.498068, 2.498062, 2.498063, 2.49806, 2.498072, 2.498064, 2.498076, 
    2.498073, 2.4981, 2.49811, 2.498115, 2.498118, 2.498127, 2.498121, 
    2.498124, 2.498118, 2.498114, 2.498116, 2.498104, 2.498109, 2.498085, 
    2.498095, 2.498068, 2.498075, 2.498067, 2.498071, 2.498064, 2.49807, 
    2.49806, 2.498057, 2.498059, 2.498053, 2.49807, 2.498064, 2.498116, 
    2.498116, 2.498114, 2.49812, 2.498121, 2.498127, 2.498122, 2.498119, 
    2.498114, 2.49811, 2.498107, 2.498101, 2.498093, 2.498082, 2.498074, 
    2.498069, 2.498072, 2.49807, 2.498073, 2.498074, 2.498058, 2.498067, 
    2.498053, 2.498054, 2.49806, 2.498054, 2.498115, 2.498117, 2.498123, 
    2.498118, 2.498127, 2.498122, 2.498119, 2.498109, 2.498106, 2.498104, 
    2.4981, 2.498094, 2.498084, 2.498075, 2.498068, 2.498068, 2.498068, 
    2.498066, 2.498071, 2.498066, 2.498065, 2.498067, 2.498054, 2.498058, 
    2.498054, 2.498057, 2.498116, 2.498114, 2.498115, 2.498112, 2.498114, 
    2.498105, 2.498102, 2.498089, 2.498094, 2.498085, 2.498093, 2.498092, 
    2.498085, 2.498093, 2.498076, 2.498087, 2.498066, 2.498078, 2.498066, 
    2.498068, 2.498064, 2.498061, 2.498057, 2.498049, 2.498051, 2.498045, 
    2.498109, 2.498105, 2.498106, 2.498101, 2.498099, 2.498092, 2.498082, 
    2.498085, 2.498078, 2.498077, 2.498088, 2.498081, 2.498103, 2.498099, 
    2.498101, 2.498109, 2.498085, 2.498097, 2.498074, 2.498081, 2.498061, 
    2.498071, 2.498052, 2.498044, 2.498036, 2.498027, 2.498103, 2.498106, 
    2.498101, 2.498095, 2.498089, 2.49808, 2.49808, 2.498078, 2.498074, 
    2.498071, 2.498078, 2.49807, 2.498098, 2.498084, 2.498107, 2.4981, 
    2.498095, 2.498097, 2.498086, 2.498083, 2.498073, 2.498078, 2.498046, 
    2.49806, 2.49802, 2.498032, 2.498107, 2.498103, 2.498091, 2.498097, 
    2.49808, 2.498076, 2.498073, 2.498068, 2.498068, 2.498065, 2.49807, 
    2.498065, 2.49808, 2.498074, 2.498092, 2.498088, 2.49809, 2.498092, 
    2.498085, 2.498078, 2.498077, 2.498075, 2.498068, 2.49808, 2.498044, 
    2.498066, 2.498099, 2.498092, 2.498091, 2.498094, 2.498076, 2.498083, 
    2.498065, 2.49807, 2.498062, 2.498066, 2.498067, 2.498072, 2.498075, 
    2.498082, 2.498089, 2.498094, 2.498093, 2.498087, 2.498077, 2.498068, 
    2.49807, 2.498063, 2.498081, 2.498074, 2.498076, 2.498069, 2.498086, 
    2.498071, 2.498089, 2.498088, 2.498083, 2.498073, 2.498071, 2.498069, 
    2.49807, 2.498077, 2.498078, 2.498083, 2.498084, 2.498088, 2.498091, 
    2.498088, 2.498085, 2.498077, 2.498069, 2.498061, 2.498059, 2.498049, 
    2.498057, 2.498044, 2.498055, 2.498036, 2.49807, 2.498055, 2.498083, 
    2.49808, 2.498075, 2.498062, 2.498069, 2.498061, 2.498078, 2.498087, 
    2.498089, 2.498093, 2.498089, 2.49809, 2.498085, 2.498087, 2.498077, 
    2.498082, 2.498067, 2.498061, 2.498045, 2.498036, 2.498026, 2.498022, 
    2.49802, 2.49802,
  2.498261, 2.498253, 2.498254, 2.498248, 2.498251, 2.498247, 2.498259, 
    2.498252, 2.498256, 2.49826, 2.498235, 2.498247, 2.498222, 2.49823, 
    2.49821, 2.498223, 2.498207, 2.49821, 2.498201, 2.498204, 2.498192, 
    2.4982, 2.498186, 2.498194, 2.498193, 2.4982, 2.498245, 2.498236, 
    2.498245, 2.498244, 2.498245, 2.498251, 2.498254, 2.498261, 2.49826, 
    2.498255, 2.498244, 2.498247, 2.498238, 2.498238, 2.498227, 2.498232, 
    2.498214, 2.498219, 2.498204, 2.498208, 2.498204, 2.498205, 2.498204, 
    2.498209, 2.498207, 2.498212, 2.498231, 2.498225, 2.498242, 2.498252, 
    2.498259, 2.498263, 2.498263, 2.498261, 2.498255, 2.498249, 2.498244, 
    2.498241, 2.498238, 2.498229, 2.498224, 2.498213, 2.498214, 2.498211, 
    2.498208, 2.498202, 2.498203, 2.498201, 2.498211, 2.498204, 2.498216, 
    2.498213, 2.498237, 2.498246, 2.49825, 2.498254, 2.498262, 2.498256, 
    2.498259, 2.498253, 2.49825, 2.498251, 2.498241, 2.498245, 2.498223, 
    2.498233, 2.498208, 2.498214, 2.498207, 2.49821, 2.498204, 2.49821, 
    2.4982, 2.498198, 2.498199, 2.498194, 2.49821, 2.498204, 2.498251, 
    2.498251, 2.49825, 2.498256, 2.498256, 2.498261, 2.498257, 2.498255, 
    2.49825, 2.498247, 2.498244, 2.498237, 2.49823, 2.498221, 2.498214, 
    2.498209, 2.498212, 2.498209, 2.498212, 2.498214, 2.498199, 2.498207, 
    2.498194, 2.498195, 2.498201, 2.498195, 2.498251, 2.498253, 2.498258, 
    2.498254, 2.498262, 2.498257, 2.498255, 2.498245, 2.498243, 2.498241, 
    2.498237, 2.498232, 2.498223, 2.498215, 2.498208, 2.498208, 2.498208, 
    2.498206, 2.49821, 2.498206, 2.498205, 2.498207, 2.498195, 2.498199, 
    2.498195, 2.498197, 2.498252, 2.49825, 2.498251, 2.498248, 2.49825, 
    2.498241, 2.498239, 2.498227, 2.498232, 2.498224, 2.498231, 2.49823, 
    2.498224, 2.49823, 2.498215, 2.498226, 2.498206, 2.498217, 2.498206, 
    2.498208, 2.498204, 2.498201, 2.498198, 2.498191, 2.498192, 2.498187, 
    2.498245, 2.498242, 2.498242, 2.498239, 2.498236, 2.49823, 2.49822, 
    2.498224, 2.498217, 2.498216, 2.498226, 2.49822, 2.49824, 2.498236, 
    2.498238, 2.498245, 2.498223, 2.498235, 2.498214, 2.49822, 2.498202, 
    2.498211, 2.498193, 2.498186, 2.498179, 2.49817, 2.49824, 2.498242, 
    2.498238, 2.498232, 2.498227, 2.498219, 2.498219, 2.498217, 2.498214, 
    2.498211, 2.498217, 2.49821, 2.498236, 2.498222, 2.498243, 2.498237, 
    2.498232, 2.498235, 2.498224, 2.498222, 2.498212, 2.498217, 2.498188, 
    2.498201, 2.498164, 2.498174, 2.498243, 2.49824, 2.498229, 2.498234, 
    2.498219, 2.498215, 2.498212, 2.498208, 2.498208, 2.498205, 2.498209, 
    2.498205, 2.498219, 2.498213, 2.49823, 2.498226, 2.498228, 2.49823, 
    2.498224, 2.498217, 2.498217, 2.498214, 2.498208, 2.498219, 2.498186, 
    2.498206, 2.498236, 2.49823, 2.498229, 2.498232, 2.498215, 2.498221, 
    2.498205, 2.49821, 2.498203, 2.498206, 2.498207, 2.498211, 2.498214, 
    2.498221, 2.498227, 2.498231, 2.49823, 2.498225, 2.498216, 2.498208, 
    2.498209, 2.498203, 2.49822, 2.498213, 2.498216, 2.498209, 2.498224, 
    2.498211, 2.498227, 2.498226, 2.498221, 2.498212, 2.49821, 2.498208, 
    2.49821, 2.498216, 2.498217, 2.498222, 2.498223, 2.498226, 2.498229, 
    2.498227, 2.498224, 2.498216, 2.498209, 2.498201, 2.498199, 2.498191, 
    2.498198, 2.498186, 2.498196, 2.498178, 2.49821, 2.498196, 2.498221, 
    2.498219, 2.498214, 2.498203, 2.498209, 2.498202, 2.498217, 2.498225, 
    2.498227, 2.498231, 2.498227, 2.498228, 2.498224, 2.498225, 2.498216, 
    2.498221, 2.498207, 2.498202, 2.498187, 2.498178, 2.498169, 2.498165, 
    2.498164, 2.498164,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  5.978417e-08, 6.004782e-08, 5.999657e-08, 6.020921e-08, 6.009125e-08, 
    6.023049e-08, 5.983763e-08, 6.005828e-08, 5.991742e-08, 5.980792e-08, 
    6.062189e-08, 6.02187e-08, 6.10408e-08, 6.078362e-08, 6.142971e-08, 
    6.100077e-08, 6.15162e-08, 6.141735e-08, 6.171493e-08, 6.162968e-08, 
    6.201029e-08, 6.175428e-08, 6.220762e-08, 6.194915e-08, 6.198958e-08, 
    6.174583e-08, 6.029985e-08, 6.057169e-08, 6.028374e-08, 6.032251e-08, 
    6.030511e-08, 6.009369e-08, 5.998714e-08, 5.976403e-08, 5.980453e-08, 
    5.996841e-08, 6.033994e-08, 6.021382e-08, 6.053169e-08, 6.052451e-08, 
    6.087841e-08, 6.071884e-08, 6.131371e-08, 6.114463e-08, 6.163324e-08, 
    6.151035e-08, 6.162746e-08, 6.159195e-08, 6.162792e-08, 6.14477e-08, 
    6.152491e-08, 6.136634e-08, 6.074872e-08, 6.093022e-08, 6.038891e-08, 
    6.006344e-08, 5.98473e-08, 5.969392e-08, 5.971561e-08, 5.975694e-08, 
    5.996937e-08, 6.016911e-08, 6.032133e-08, 6.042315e-08, 6.052348e-08, 
    6.082715e-08, 6.098792e-08, 6.134788e-08, 6.128293e-08, 6.139297e-08, 
    6.149813e-08, 6.167465e-08, 6.164559e-08, 6.172336e-08, 6.139008e-08, 
    6.161157e-08, 6.124593e-08, 6.134594e-08, 6.055071e-08, 6.024785e-08, 
    6.011908e-08, 6.000641e-08, 5.973228e-08, 5.992159e-08, 5.984696e-08, 
    6.002452e-08, 6.013734e-08, 6.008154e-08, 6.042593e-08, 6.029204e-08, 
    6.099744e-08, 6.069359e-08, 6.148586e-08, 6.129627e-08, 6.153131e-08, 
    6.141137e-08, 6.161687e-08, 6.143193e-08, 6.175231e-08, 6.182207e-08, 
    6.17744e-08, 6.195755e-08, 6.142167e-08, 6.162745e-08, 6.007998e-08, 
    6.008907e-08, 6.013147e-08, 5.994509e-08, 5.99337e-08, 5.976292e-08, 
    5.991488e-08, 5.997959e-08, 6.014388e-08, 6.024105e-08, 6.033343e-08, 
    6.053654e-08, 6.076338e-08, 6.108062e-08, 6.130855e-08, 6.146134e-08, 
    6.136766e-08, 6.145037e-08, 6.135791e-08, 6.131457e-08, 6.179593e-08, 
    6.152563e-08, 6.19312e-08, 6.190876e-08, 6.172521e-08, 6.191129e-08, 
    6.009547e-08, 6.00431e-08, 5.986127e-08, 6.000356e-08, 5.974432e-08, 
    5.988942e-08, 5.997286e-08, 6.029482e-08, 6.036558e-08, 6.043117e-08, 
    6.056074e-08, 6.0727e-08, 6.10187e-08, 6.127252e-08, 6.150425e-08, 
    6.148726e-08, 6.149325e-08, 6.1545e-08, 6.141678e-08, 6.156606e-08, 
    6.159111e-08, 6.15256e-08, 6.190576e-08, 6.179715e-08, 6.190829e-08, 
    6.183758e-08, 6.006012e-08, 6.014824e-08, 6.010062e-08, 6.019016e-08, 
    6.012708e-08, 6.040757e-08, 6.049168e-08, 6.088524e-08, 6.072373e-08, 
    6.09808e-08, 6.074985e-08, 6.079077e-08, 6.098916e-08, 6.076233e-08, 
    6.125851e-08, 6.092209e-08, 6.154701e-08, 6.121103e-08, 6.156807e-08, 
    6.150324e-08, 6.161059e-08, 6.170672e-08, 6.182767e-08, 6.205084e-08, 
    6.199917e-08, 6.218581e-08, 6.027961e-08, 6.03939e-08, 6.038385e-08, 
    6.050347e-08, 6.059194e-08, 6.078369e-08, 6.109126e-08, 6.09756e-08, 
    6.118793e-08, 6.123056e-08, 6.090797e-08, 6.110603e-08, 6.047041e-08, 
    6.057309e-08, 6.051196e-08, 6.028862e-08, 6.100223e-08, 6.063599e-08, 
    6.131232e-08, 6.11139e-08, 6.169301e-08, 6.140499e-08, 6.197072e-08, 
    6.221256e-08, 6.244021e-08, 6.270623e-08, 6.045629e-08, 6.037863e-08, 
    6.05177e-08, 6.071009e-08, 6.088864e-08, 6.1126e-08, 6.115029e-08, 
    6.119475e-08, 6.130995e-08, 6.14068e-08, 6.120881e-08, 6.143108e-08, 
    6.059688e-08, 6.103403e-08, 6.034927e-08, 6.055544e-08, 6.069875e-08, 
    6.06359e-08, 6.096239e-08, 6.103933e-08, 6.135203e-08, 6.119039e-08, 
    6.215286e-08, 6.172701e-08, 6.290882e-08, 6.257852e-08, 6.03515e-08, 
    6.045603e-08, 6.081986e-08, 6.064675e-08, 6.114185e-08, 6.126373e-08, 
    6.13628e-08, 6.148945e-08, 6.150314e-08, 6.157818e-08, 6.145521e-08, 
    6.157332e-08, 6.112651e-08, 6.132618e-08, 6.077828e-08, 6.091162e-08, 
    6.085028e-08, 6.078299e-08, 6.099067e-08, 6.121192e-08, 6.121667e-08, 
    6.128761e-08, 6.14875e-08, 6.114386e-08, 6.22078e-08, 6.155069e-08, 
    6.057002e-08, 6.077136e-08, 6.080015e-08, 6.072214e-08, 6.125151e-08, 
    6.105969e-08, 6.157635e-08, 6.143672e-08, 6.166551e-08, 6.155182e-08, 
    6.153508e-08, 6.138907e-08, 6.129815e-08, 6.106848e-08, 6.088162e-08, 
    6.073346e-08, 6.076791e-08, 6.093067e-08, 6.122546e-08, 6.150437e-08, 
    6.144327e-08, 6.164812e-08, 6.110595e-08, 6.133328e-08, 6.124541e-08, 
    6.147453e-08, 6.097252e-08, 6.139996e-08, 6.086326e-08, 6.091032e-08, 
    6.105589e-08, 6.134869e-08, 6.141349e-08, 6.148266e-08, 6.143998e-08, 
    6.123295e-08, 6.119904e-08, 6.105235e-08, 6.101184e-08, 6.090008e-08, 
    6.080754e-08, 6.089208e-08, 6.098087e-08, 6.123304e-08, 6.14603e-08, 
    6.170809e-08, 6.176873e-08, 6.205823e-08, 6.182255e-08, 6.221146e-08, 
    6.188078e-08, 6.245322e-08, 6.142476e-08, 6.187108e-08, 6.106251e-08, 
    6.114962e-08, 6.130716e-08, 6.166854e-08, 6.147345e-08, 6.170161e-08, 
    6.119771e-08, 6.093627e-08, 6.086865e-08, 6.074247e-08, 6.087154e-08, 
    6.086104e-08, 6.098455e-08, 6.094486e-08, 6.124142e-08, 6.108212e-08, 
    6.153466e-08, 6.169981e-08, 6.216625e-08, 6.24522e-08, 6.274332e-08, 
    6.287184e-08, 6.291096e-08, 6.292732e-08 ;

 SOIL1_HR_S3 =
  7.095026e-10, 7.126326e-10, 7.120242e-10, 7.145488e-10, 7.131484e-10, 
    7.148015e-10, 7.101373e-10, 7.127569e-10, 7.110846e-10, 7.097845e-10, 
    7.194483e-10, 7.146614e-10, 7.244219e-10, 7.213685e-10, 7.290393e-10, 
    7.239466e-10, 7.300663e-10, 7.288926e-10, 7.324258e-10, 7.314136e-10, 
    7.359326e-10, 7.32893e-10, 7.382756e-10, 7.352068e-10, 7.356868e-10, 
    7.327927e-10, 7.156249e-10, 7.188523e-10, 7.154337e-10, 7.158939e-10, 
    7.156874e-10, 7.131772e-10, 7.119123e-10, 7.092635e-10, 7.097444e-10, 
    7.116899e-10, 7.161008e-10, 7.146036e-10, 7.183774e-10, 7.182922e-10, 
    7.224938e-10, 7.205994e-10, 7.27662e-10, 7.256546e-10, 7.314558e-10, 
    7.299968e-10, 7.313873e-10, 7.309657e-10, 7.313927e-10, 7.29253e-10, 
    7.301697e-10, 7.282869e-10, 7.209541e-10, 7.23109e-10, 7.166823e-10, 
    7.128181e-10, 7.102521e-10, 7.084312e-10, 7.086886e-10, 7.091793e-10, 
    7.117013e-10, 7.140726e-10, 7.158799e-10, 7.170888e-10, 7.182799e-10, 
    7.218853e-10, 7.237941e-10, 7.280679e-10, 7.272967e-10, 7.286032e-10, 
    7.298517e-10, 7.319475e-10, 7.316026e-10, 7.325259e-10, 7.285689e-10, 
    7.311987e-10, 7.268574e-10, 7.280447e-10, 7.186032e-10, 7.150076e-10, 
    7.134788e-10, 7.121411e-10, 7.088866e-10, 7.11134e-10, 7.10248e-10, 
    7.123561e-10, 7.136955e-10, 7.13033e-10, 7.171218e-10, 7.155321e-10, 
    7.239072e-10, 7.202996e-10, 7.29706e-10, 7.27455e-10, 7.302456e-10, 
    7.288217e-10, 7.312616e-10, 7.290656e-10, 7.328697e-10, 7.336979e-10, 
    7.331319e-10, 7.353065e-10, 7.289439e-10, 7.313872e-10, 7.130145e-10, 
    7.131225e-10, 7.136259e-10, 7.114132e-10, 7.112778e-10, 7.092503e-10, 
    7.110544e-10, 7.118227e-10, 7.137732e-10, 7.149268e-10, 7.160236e-10, 
    7.18435e-10, 7.211283e-10, 7.248947e-10, 7.276009e-10, 7.29415e-10, 
    7.283026e-10, 7.292847e-10, 7.281868e-10, 7.276724e-10, 7.333875e-10, 
    7.301783e-10, 7.349937e-10, 7.347272e-10, 7.325479e-10, 7.347573e-10, 
    7.131983e-10, 7.125767e-10, 7.104179e-10, 7.121073e-10, 7.090295e-10, 
    7.107522e-10, 7.117428e-10, 7.155652e-10, 7.164053e-10, 7.17184e-10, 
    7.187222e-10, 7.206963e-10, 7.241595e-10, 7.27173e-10, 7.299243e-10, 
    7.297227e-10, 7.297937e-10, 7.304083e-10, 7.288859e-10, 7.306582e-10, 
    7.309556e-10, 7.301779e-10, 7.346915e-10, 7.33402e-10, 7.347216e-10, 
    7.33882e-10, 7.127787e-10, 7.138249e-10, 7.132596e-10, 7.143226e-10, 
    7.135736e-10, 7.169039e-10, 7.179023e-10, 7.22575e-10, 7.206574e-10, 
    7.237095e-10, 7.209675e-10, 7.214533e-10, 7.238088e-10, 7.211157e-10, 
    7.270068e-10, 7.230125e-10, 7.304322e-10, 7.26443e-10, 7.306821e-10, 
    7.299124e-10, 7.311869e-10, 7.323283e-10, 7.337644e-10, 7.364142e-10, 
    7.358006e-10, 7.380167e-10, 7.153846e-10, 7.167416e-10, 7.166222e-10, 
    7.180423e-10, 7.190927e-10, 7.213693e-10, 7.250209e-10, 7.236478e-10, 
    7.261688e-10, 7.266749e-10, 7.228449e-10, 7.251963e-10, 7.176498e-10, 
    7.188689e-10, 7.181431e-10, 7.154916e-10, 7.239641e-10, 7.196157e-10, 
    7.276456e-10, 7.252898e-10, 7.321656e-10, 7.287459e-10, 7.354628e-10, 
    7.383342e-10, 7.410373e-10, 7.441959e-10, 7.174822e-10, 7.165602e-10, 
    7.182113e-10, 7.204955e-10, 7.226153e-10, 7.254334e-10, 7.257219e-10, 
    7.262498e-10, 7.276175e-10, 7.287674e-10, 7.264166e-10, 7.290556e-10, 
    7.191514e-10, 7.243415e-10, 7.162115e-10, 7.186594e-10, 7.203609e-10, 
    7.196146e-10, 7.234909e-10, 7.244044e-10, 7.281171e-10, 7.261979e-10, 
    7.376254e-10, 7.325693e-10, 7.466013e-10, 7.426795e-10, 7.16238e-10, 
    7.174791e-10, 7.217987e-10, 7.197434e-10, 7.256216e-10, 7.270686e-10, 
    7.28245e-10, 7.297487e-10, 7.299111e-10, 7.308021e-10, 7.293421e-10, 
    7.307445e-10, 7.254394e-10, 7.278101e-10, 7.213051e-10, 7.228882e-10, 
    7.221599e-10, 7.21361e-10, 7.238267e-10, 7.264536e-10, 7.265099e-10, 
    7.273522e-10, 7.297256e-10, 7.256455e-10, 7.382777e-10, 7.304757e-10, 
    7.188325e-10, 7.21223e-10, 7.215646e-10, 7.206386e-10, 7.269235e-10, 
    7.246462e-10, 7.307804e-10, 7.291225e-10, 7.31839e-10, 7.304891e-10, 
    7.302905e-10, 7.285568e-10, 7.274774e-10, 7.247505e-10, 7.22532e-10, 
    7.207729e-10, 7.211819e-10, 7.231143e-10, 7.266143e-10, 7.299258e-10, 
    7.292004e-10, 7.316325e-10, 7.251954e-10, 7.278945e-10, 7.268512e-10, 
    7.295715e-10, 7.236113e-10, 7.286862e-10, 7.223141e-10, 7.228728e-10, 
    7.24601e-10, 7.280774e-10, 7.288468e-10, 7.29668e-10, 7.291613e-10, 
    7.267033e-10, 7.263006e-10, 7.24559e-10, 7.240781e-10, 7.227511e-10, 
    7.216525e-10, 7.226562e-10, 7.237103e-10, 7.267043e-10, 7.294025e-10, 
    7.323445e-10, 7.330646e-10, 7.365019e-10, 7.337035e-10, 7.383212e-10, 
    7.34395e-10, 7.411918e-10, 7.289805e-10, 7.342798e-10, 7.246796e-10, 
    7.257139e-10, 7.275843e-10, 7.318749e-10, 7.295587e-10, 7.322676e-10, 
    7.262848e-10, 7.231809e-10, 7.22378e-10, 7.208799e-10, 7.224123e-10, 
    7.222877e-10, 7.237541e-10, 7.232829e-10, 7.268037e-10, 7.249125e-10, 
    7.302854e-10, 7.322463e-10, 7.377844e-10, 7.411796e-10, 7.446363e-10, 
    7.461624e-10, 7.466268e-10, 7.46821e-10 ;

 SOIL2C =
  5.783956, 5.783962, 5.78396, 5.783966, 5.783963, 5.783966, 5.783957, 
    5.783962, 5.783959, 5.783956, 5.783975, 5.783966, 5.783984, 5.783978, 
    5.783993, 5.783983, 5.783995, 5.783993, 5.784, 5.783998, 5.784007, 5.784, 
    5.784011, 5.784005, 5.784006, 5.784, 5.783967, 5.783974, 5.783967, 
    5.783968, 5.783967, 5.783963, 5.78396, 5.783955, 5.783956, 5.78396, 
    5.783968, 5.783966, 5.783973, 5.783973, 5.783981, 5.783977, 5.78399, 
    5.783987, 5.783998, 5.783995, 5.783998, 5.783997, 5.783998, 5.783994, 
    5.783995, 5.783992, 5.783978, 5.783982, 5.783969, 5.783962, 5.783957, 
    5.783954, 5.783954, 5.783955, 5.78396, 5.783965, 5.783968, 5.78397, 
    5.783973, 5.783979, 5.783983, 5.783991, 5.78399, 5.783992, 5.783995, 
    5.783999, 5.783998, 5.784, 5.783992, 5.783998, 5.783989, 5.783991, 
    5.783973, 5.783966, 5.783963, 5.783961, 5.783955, 5.783959, 5.783957, 
    5.783961, 5.783964, 5.783962, 5.78397, 5.783967, 5.783983, 5.783977, 
    5.783995, 5.78399, 5.783996, 5.783993, 5.783998, 5.783993, 5.784, 
    5.784002, 5.784001, 5.784005, 5.783993, 5.783998, 5.783962, 5.783963, 
    5.783964, 5.783959, 5.783959, 5.783955, 5.783959, 5.78396, 5.783964, 
    5.783966, 5.783968, 5.783973, 5.783978, 5.783985, 5.78399, 5.783994, 
    5.783992, 5.783994, 5.783992, 5.78399, 5.784001, 5.783996, 5.784005, 
    5.784004, 5.784, 5.784004, 5.783963, 5.783962, 5.783957, 5.783961, 
    5.783955, 5.783958, 5.78396, 5.783967, 5.783969, 5.78397, 5.783973, 
    5.783977, 5.783984, 5.783989, 5.783995, 5.783995, 5.783995, 5.783996, 
    5.783993, 5.783996, 5.783997, 5.783996, 5.784004, 5.784002, 5.784004, 
    5.784002, 5.783962, 5.783964, 5.783963, 5.783965, 5.783964, 5.78397, 
    5.783972, 5.783981, 5.783977, 5.783983, 5.783978, 5.783978, 5.783983, 
    5.783978, 5.783989, 5.783982, 5.783996, 5.783988, 5.783997, 5.783995, 
    5.783998, 5.783999, 5.784002, 5.784008, 5.784006, 5.78401, 5.783967, 
    5.783969, 5.783969, 5.783972, 5.783974, 5.783978, 5.783986, 5.783983, 
    5.783988, 5.783988, 5.783981, 5.783986, 5.783971, 5.783974, 5.783972, 
    5.783967, 5.783984, 5.783975, 5.78399, 5.783986, 5.783999, 5.783993, 
    5.784006, 5.784011, 5.784016, 5.784022, 5.783971, 5.783969, 5.783972, 
    5.783977, 5.783981, 5.783986, 5.783987, 5.783988, 5.78399, 5.783993, 
    5.783988, 5.783993, 5.783974, 5.783984, 5.783968, 5.783973, 5.783977, 
    5.783975, 5.783983, 5.783984, 5.783991, 5.783988, 5.78401, 5.784, 
    5.784027, 5.784019, 5.783968, 5.783971, 5.783979, 5.783976, 5.783987, 
    5.783989, 5.783992, 5.783995, 5.783995, 5.783997, 5.783994, 5.783997, 
    5.783986, 5.783991, 5.783978, 5.783981, 5.78398, 5.783978, 5.783983, 
    5.783988, 5.783988, 5.78399, 5.783995, 5.783987, 5.784011, 5.783996, 
    5.783974, 5.783978, 5.783979, 5.783977, 5.783989, 5.783985, 5.783997, 
    5.783993, 5.783998, 5.783996, 5.783996, 5.783992, 5.78399, 5.783985, 
    5.783981, 5.783978, 5.783978, 5.783982, 5.783988, 5.783995, 5.783994, 
    5.783998, 5.783986, 5.783991, 5.783989, 5.783994, 5.783983, 5.783993, 
    5.78398, 5.783981, 5.783985, 5.783991, 5.783993, 5.783994, 5.783993, 
    5.783989, 5.783988, 5.783985, 5.783984, 5.783981, 5.783979, 5.783981, 
    5.783983, 5.783989, 5.783994, 5.783999, 5.784001, 5.784008, 5.784002, 
    5.784011, 5.784004, 5.784017, 5.783993, 5.784003, 5.783985, 5.783987, 
    5.78399, 5.783998, 5.783994, 5.783999, 5.783988, 5.783982, 5.78398, 
    5.783978, 5.78398, 5.78398, 5.783983, 5.783982, 5.783989, 5.783985, 
    5.783996, 5.783999, 5.78401, 5.784017, 5.784023, 5.784026, 5.784027, 
    5.784028 ;

 SOIL2C_TO_SOIL1C =
  1.057637e-09, 1.062304e-09, 1.061397e-09, 1.065162e-09, 1.063073e-09, 
    1.065538e-09, 1.058583e-09, 1.062489e-09, 1.059996e-09, 1.058057e-09, 
    1.072468e-09, 1.06533e-09, 1.079884e-09, 1.075331e-09, 1.086769e-09, 
    1.079175e-09, 1.088301e-09, 1.08655e-09, 1.091819e-09, 1.090309e-09, 
    1.097048e-09, 1.092515e-09, 1.100541e-09, 1.095966e-09, 1.096681e-09, 
    1.092366e-09, 1.066766e-09, 1.071579e-09, 1.066481e-09, 1.067167e-09, 
    1.066859e-09, 1.063116e-09, 1.06123e-09, 1.05728e-09, 1.057997e-09, 
    1.060898e-09, 1.067476e-09, 1.065243e-09, 1.070871e-09, 1.070744e-09, 
    1.077009e-09, 1.074184e-09, 1.084715e-09, 1.081722e-09, 1.090372e-09, 
    1.088197e-09, 1.09027e-09, 1.089642e-09, 1.090278e-09, 1.087088e-09, 
    1.088455e-09, 1.085647e-09, 1.074713e-09, 1.077926e-09, 1.068343e-09, 
    1.062581e-09, 1.058754e-09, 1.056039e-09, 1.056423e-09, 1.057155e-09, 
    1.060915e-09, 1.064452e-09, 1.067146e-09, 1.068949e-09, 1.070725e-09, 
    1.076102e-09, 1.078948e-09, 1.085321e-09, 1.084171e-09, 1.086119e-09, 
    1.08798e-09, 1.091106e-09, 1.090591e-09, 1.091968e-09, 1.086068e-09, 
    1.089989e-09, 1.083516e-09, 1.085286e-09, 1.071207e-09, 1.065846e-09, 
    1.063566e-09, 1.061571e-09, 1.056718e-09, 1.060069e-09, 1.058748e-09, 
    1.061892e-09, 1.063889e-09, 1.062901e-09, 1.068998e-09, 1.066628e-09, 
    1.079116e-09, 1.073737e-09, 1.087763e-09, 1.084407e-09, 1.088568e-09, 
    1.086445e-09, 1.090083e-09, 1.086808e-09, 1.092481e-09, 1.093716e-09, 
    1.092872e-09, 1.096114e-09, 1.086627e-09, 1.09027e-09, 1.062874e-09, 
    1.063035e-09, 1.063785e-09, 1.060486e-09, 1.060284e-09, 1.057261e-09, 
    1.059951e-09, 1.061096e-09, 1.064005e-09, 1.065725e-09, 1.067361e-09, 
    1.070957e-09, 1.074973e-09, 1.080589e-09, 1.084624e-09, 1.087329e-09, 
    1.085671e-09, 1.087135e-09, 1.085498e-09, 1.084731e-09, 1.093253e-09, 
    1.088467e-09, 1.095648e-09, 1.09525e-09, 1.092001e-09, 1.095295e-09, 
    1.063148e-09, 1.062221e-09, 1.059002e-09, 1.061521e-09, 1.056931e-09, 
    1.0595e-09, 1.060977e-09, 1.066677e-09, 1.06793e-09, 1.069091e-09, 
    1.071385e-09, 1.074329e-09, 1.079493e-09, 1.083986e-09, 1.088089e-09, 
    1.087788e-09, 1.087894e-09, 1.08881e-09, 1.08654e-09, 1.089183e-09, 
    1.089627e-09, 1.088467e-09, 1.095197e-09, 1.093274e-09, 1.095242e-09, 
    1.09399e-09, 1.062522e-09, 1.064082e-09, 1.063239e-09, 1.064824e-09, 
    1.063707e-09, 1.068673e-09, 1.070162e-09, 1.07713e-09, 1.074271e-09, 
    1.078822e-09, 1.074733e-09, 1.075457e-09, 1.07897e-09, 1.074954e-09, 
    1.083738e-09, 1.077782e-09, 1.088846e-09, 1.082898e-09, 1.089219e-09, 
    1.088071e-09, 1.089971e-09, 1.091673e-09, 1.093815e-09, 1.097766e-09, 
    1.096851e-09, 1.100155e-09, 1.066408e-09, 1.068431e-09, 1.068253e-09, 
    1.070371e-09, 1.071937e-09, 1.075332e-09, 1.080777e-09, 1.07873e-09, 
    1.082489e-09, 1.083243e-09, 1.077532e-09, 1.081039e-09, 1.069786e-09, 
    1.071603e-09, 1.070521e-09, 1.066568e-09, 1.079201e-09, 1.072717e-09, 
    1.084691e-09, 1.081178e-09, 1.091431e-09, 1.086332e-09, 1.096347e-09, 
    1.100629e-09, 1.104659e-09, 1.109369e-09, 1.069536e-09, 1.068161e-09, 
    1.070623e-09, 1.074029e-09, 1.07719e-09, 1.081392e-09, 1.081822e-09, 
    1.08261e-09, 1.084649e-09, 1.086364e-09, 1.082858e-09, 1.086793e-09, 
    1.072025e-09, 1.079764e-09, 1.067641e-09, 1.071291e-09, 1.073828e-09, 
    1.072716e-09, 1.078496e-09, 1.079858e-09, 1.085394e-09, 1.082532e-09, 
    1.099572e-09, 1.092033e-09, 1.112956e-09, 1.107108e-09, 1.06768e-09, 
    1.069531e-09, 1.075972e-09, 1.072908e-09, 1.081673e-09, 1.083831e-09, 
    1.085585e-09, 1.087827e-09, 1.088069e-09, 1.089398e-09, 1.087221e-09, 
    1.089312e-09, 1.081401e-09, 1.084936e-09, 1.075236e-09, 1.077597e-09, 
    1.076511e-09, 1.07532e-09, 1.078996e-09, 1.082914e-09, 1.082997e-09, 
    1.084253e-09, 1.087792e-09, 1.081709e-09, 1.100545e-09, 1.088911e-09, 
    1.071549e-09, 1.075114e-09, 1.075623e-09, 1.074242e-09, 1.083614e-09, 
    1.080218e-09, 1.089365e-09, 1.086893e-09, 1.090944e-09, 1.088931e-09, 
    1.088635e-09, 1.08605e-09, 1.08444e-09, 1.080374e-09, 1.077066e-09, 
    1.074443e-09, 1.075053e-09, 1.077934e-09, 1.083153e-09, 1.088091e-09, 
    1.087009e-09, 1.090636e-09, 1.081037e-09, 1.085062e-09, 1.083506e-09, 
    1.087563e-09, 1.078675e-09, 1.086243e-09, 1.076741e-09, 1.077574e-09, 
    1.080151e-09, 1.085335e-09, 1.086482e-09, 1.087707e-09, 1.086951e-09, 
    1.083286e-09, 1.082685e-09, 1.080088e-09, 1.079371e-09, 1.077393e-09, 
    1.075754e-09, 1.077251e-09, 1.078823e-09, 1.083287e-09, 1.087311e-09, 
    1.091698e-09, 1.092771e-09, 1.097897e-09, 1.093724e-09, 1.100609e-09, 
    1.094755e-09, 1.10489e-09, 1.086682e-09, 1.094583e-09, 1.080268e-09, 
    1.08181e-09, 1.0846e-09, 1.090997e-09, 1.087544e-09, 1.091583e-09, 
    1.082662e-09, 1.078033e-09, 1.076836e-09, 1.074602e-09, 1.076887e-09, 
    1.076702e-09, 1.078888e-09, 1.078186e-09, 1.083436e-09, 1.080615e-09, 
    1.088627e-09, 1.091551e-09, 1.099809e-09, 1.104872e-09, 1.110026e-09, 
    1.112301e-09, 1.112994e-09, 1.113283e-09 ;

 SOIL2C_TO_SOIL3C =
  7.554549e-11, 7.587887e-11, 7.581407e-11, 7.608297e-11, 7.593381e-11, 
    7.610988e-11, 7.561308e-11, 7.589211e-11, 7.571398e-11, 7.55755e-11, 
    7.660483e-11, 7.609497e-11, 7.713456e-11, 7.680935e-11, 7.762637e-11, 
    7.708395e-11, 7.773576e-11, 7.761074e-11, 7.798705e-11, 7.787924e-11, 
    7.836055e-11, 7.803681e-11, 7.86101e-11, 7.828325e-11, 7.833437e-11, 
    7.802613e-11, 7.619759e-11, 7.654134e-11, 7.617722e-11, 7.622624e-11, 
    7.620424e-11, 7.593688e-11, 7.580214e-11, 7.552001e-11, 7.557124e-11, 
    7.577846e-11, 7.624828e-11, 7.60888e-11, 7.649077e-11, 7.648169e-11, 
    7.692921e-11, 7.672743e-11, 7.747968e-11, 7.726587e-11, 7.788375e-11, 
    7.772835e-11, 7.787644e-11, 7.783154e-11, 7.787703e-11, 7.764912e-11, 
    7.774677e-11, 7.754623e-11, 7.676521e-11, 7.699473e-11, 7.631022e-11, 
    7.589863e-11, 7.562531e-11, 7.543136e-11, 7.545878e-11, 7.551105e-11, 
    7.577967e-11, 7.603226e-11, 7.622475e-11, 7.635351e-11, 7.648038e-11, 
    7.68644e-11, 7.70677e-11, 7.75229e-11, 7.744076e-11, 7.757992e-11, 
    7.771289e-11, 7.793612e-11, 7.789937e-11, 7.799772e-11, 7.757626e-11, 
    7.785635e-11, 7.739397e-11, 7.752043e-11, 7.651482e-11, 7.613183e-11, 
    7.596899e-11, 7.582652e-11, 7.547986e-11, 7.571925e-11, 7.562488e-11, 
    7.584941e-11, 7.599208e-11, 7.592152e-11, 7.635703e-11, 7.618771e-11, 
    7.707975e-11, 7.66955e-11, 7.769738e-11, 7.745762e-11, 7.775485e-11, 
    7.760319e-11, 7.786305e-11, 7.762917e-11, 7.803433e-11, 7.812255e-11, 
    7.806226e-11, 7.829386e-11, 7.761621e-11, 7.787643e-11, 7.591954e-11, 
    7.593105e-11, 7.598466e-11, 7.574898e-11, 7.573456e-11, 7.551861e-11, 
    7.571077e-11, 7.57926e-11, 7.600035e-11, 7.612323e-11, 7.624005e-11, 
    7.64969e-11, 7.678376e-11, 7.718493e-11, 7.747317e-11, 7.766638e-11, 
    7.754791e-11, 7.76525e-11, 7.753558e-11, 7.748077e-11, 7.808949e-11, 
    7.774768e-11, 7.826056e-11, 7.823218e-11, 7.800006e-11, 7.823538e-11, 
    7.593913e-11, 7.587291e-11, 7.564298e-11, 7.582292e-11, 7.549509e-11, 
    7.567858e-11, 7.578409e-11, 7.619123e-11, 7.62807e-11, 7.636365e-11, 
    7.652749e-11, 7.673776e-11, 7.710662e-11, 7.742759e-11, 7.772063e-11, 
    7.769916e-11, 7.770672e-11, 7.777217e-11, 7.761002e-11, 7.77988e-11, 
    7.783047e-11, 7.774764e-11, 7.822838e-11, 7.809103e-11, 7.823157e-11, 
    7.814215e-11, 7.589444e-11, 7.600587e-11, 7.594565e-11, 7.605887e-11, 
    7.59791e-11, 7.633381e-11, 7.644017e-11, 7.693785e-11, 7.673361e-11, 
    7.705869e-11, 7.676663e-11, 7.681838e-11, 7.706927e-11, 7.678242e-11, 
    7.740988e-11, 7.698445e-11, 7.777472e-11, 7.734983e-11, 7.780134e-11, 
    7.771936e-11, 7.78551e-11, 7.797667e-11, 7.812963e-11, 7.841185e-11, 
    7.83465e-11, 7.858253e-11, 7.617199e-11, 7.631652e-11, 7.630381e-11, 
    7.645508e-11, 7.656695e-11, 7.680944e-11, 7.719837e-11, 7.705211e-11, 
    7.732063e-11, 7.737454e-11, 7.69666e-11, 7.721705e-11, 7.641326e-11, 
    7.654311e-11, 7.646581e-11, 7.618339e-11, 7.70858e-11, 7.662266e-11, 
    7.747793e-11, 7.722701e-11, 7.795933e-11, 7.759512e-11, 7.831052e-11, 
    7.861634e-11, 7.890424e-11, 7.924063e-11, 7.639542e-11, 7.629721e-11, 
    7.647307e-11, 7.671636e-11, 7.694215e-11, 7.724231e-11, 7.727303e-11, 
    7.732926e-11, 7.747493e-11, 7.75974e-11, 7.734702e-11, 7.762811e-11, 
    7.65732e-11, 7.712601e-11, 7.626007e-11, 7.65208e-11, 7.670203e-11, 
    7.662253e-11, 7.703541e-11, 7.713271e-11, 7.752814e-11, 7.732373e-11, 
    7.854085e-11, 7.800233e-11, 7.949683e-11, 7.907914e-11, 7.62629e-11, 
    7.639508e-11, 7.685517e-11, 7.663626e-11, 7.726236e-11, 7.741647e-11, 
    7.754177e-11, 7.770192e-11, 7.771923e-11, 7.781412e-11, 7.765862e-11, 
    7.780798e-11, 7.724295e-11, 7.749545e-11, 7.680259e-11, 7.697121e-11, 
    7.689364e-11, 7.680855e-11, 7.707118e-11, 7.735097e-11, 7.735696e-11, 
    7.744667e-11, 7.769946e-11, 7.72649e-11, 7.861032e-11, 7.777935e-11, 
    7.653924e-11, 7.679385e-11, 7.683024e-11, 7.673161e-11, 7.740102e-11, 
    7.715845e-11, 7.781181e-11, 7.763522e-11, 7.792456e-11, 7.778078e-11, 
    7.775963e-11, 7.757497e-11, 7.746001e-11, 7.716958e-11, 7.693327e-11, 
    7.674592e-11, 7.678948e-11, 7.69953e-11, 7.736808e-11, 7.772078e-11, 
    7.764352e-11, 7.790257e-11, 7.721696e-11, 7.750443e-11, 7.739331e-11, 
    7.768305e-11, 7.704823e-11, 7.758875e-11, 7.691006e-11, 7.696957e-11, 
    7.715364e-11, 7.752391e-11, 7.760587e-11, 7.769333e-11, 7.763936e-11, 
    7.737756e-11, 7.733467e-11, 7.714917e-11, 7.709795e-11, 7.695661e-11, 
    7.68396e-11, 7.69465e-11, 7.705878e-11, 7.737767e-11, 7.766505e-11, 
    7.797839e-11, 7.805509e-11, 7.842118e-11, 7.812314e-11, 7.861495e-11, 
    7.819678e-11, 7.892069e-11, 7.76201e-11, 7.818451e-11, 7.716203e-11, 
    7.727217e-11, 7.74714e-11, 7.792839e-11, 7.768169e-11, 7.797021e-11, 
    7.733299e-11, 7.700239e-11, 7.691688e-11, 7.67573e-11, 7.692053e-11, 
    7.690725e-11, 7.706344e-11, 7.701325e-11, 7.738826e-11, 7.718682e-11, 
    7.775909e-11, 7.796794e-11, 7.855779e-11, 7.891939e-11, 7.928754e-11, 
    7.945007e-11, 7.949954e-11, 7.952022e-11 ;

 SOIL2C_vr =
  20.00587, 20.00588, 20.00588, 20.00589, 20.00588, 20.00589, 20.00587, 
    20.00588, 20.00587, 20.00587, 20.00592, 20.00589, 20.00594, 20.00593, 
    20.00596, 20.00594, 20.00597, 20.00596, 20.00598, 20.00598, 20.006, 
    20.00599, 20.00601, 20.006, 20.006, 20.00599, 20.0059, 20.00591, 20.0059, 
    20.0059, 20.0059, 20.00588, 20.00588, 20.00586, 20.00587, 20.00588, 
    20.0059, 20.00589, 20.00591, 20.00591, 20.00593, 20.00592, 20.00596, 
    20.00595, 20.00598, 20.00597, 20.00598, 20.00598, 20.00598, 20.00597, 
    20.00597, 20.00596, 20.00592, 20.00593, 20.0059, 20.00588, 20.00587, 
    20.00586, 20.00586, 20.00586, 20.00588, 20.00589, 20.0059, 20.0059, 
    20.00591, 20.00593, 20.00594, 20.00596, 20.00596, 20.00596, 20.00597, 
    20.00598, 20.00598, 20.00598, 20.00596, 20.00598, 20.00595, 20.00596, 
    20.00591, 20.00589, 20.00588, 20.00588, 20.00586, 20.00587, 20.00587, 
    20.00588, 20.00589, 20.00588, 20.0059, 20.0059, 20.00594, 20.00592, 
    20.00597, 20.00596, 20.00597, 20.00596, 20.00598, 20.00597, 20.00599, 
    20.00599, 20.00599, 20.006, 20.00596, 20.00598, 20.00588, 20.00588, 
    20.00589, 20.00587, 20.00587, 20.00586, 20.00587, 20.00588, 20.00589, 
    20.00589, 20.0059, 20.00591, 20.00592, 20.00594, 20.00596, 20.00597, 
    20.00596, 20.00597, 20.00596, 20.00596, 20.00599, 20.00597, 20.006, 
    20.00599, 20.00598, 20.00599, 20.00588, 20.00588, 20.00587, 20.00588, 
    20.00586, 20.00587, 20.00588, 20.0059, 20.0059, 20.00591, 20.00591, 
    20.00592, 20.00594, 20.00595, 20.00597, 20.00597, 20.00597, 20.00597, 
    20.00596, 20.00597, 20.00598, 20.00597, 20.00599, 20.00599, 20.00599, 
    20.00599, 20.00588, 20.00589, 20.00588, 20.00589, 20.00589, 20.0059, 
    20.00591, 20.00593, 20.00592, 20.00594, 20.00592, 20.00593, 20.00594, 
    20.00592, 20.00595, 20.00593, 20.00597, 20.00595, 20.00597, 20.00597, 
    20.00598, 20.00598, 20.00599, 20.006, 20.006, 20.00601, 20.0059, 20.0059, 
    20.0059, 20.00591, 20.00591, 20.00593, 20.00595, 20.00594, 20.00595, 
    20.00595, 20.00593, 20.00595, 20.00591, 20.00591, 20.00591, 20.0059, 
    20.00594, 20.00592, 20.00596, 20.00595, 20.00598, 20.00596, 20.006, 
    20.00601, 20.00603, 20.00604, 20.00591, 20.0059, 20.00591, 20.00592, 
    20.00593, 20.00595, 20.00595, 20.00595, 20.00596, 20.00596, 20.00595, 
    20.00597, 20.00591, 20.00594, 20.0059, 20.00591, 20.00592, 20.00592, 
    20.00594, 20.00594, 20.00596, 20.00595, 20.00601, 20.00598, 20.00606, 
    20.00603, 20.0059, 20.00591, 20.00593, 20.00592, 20.00595, 20.00595, 
    20.00596, 20.00597, 20.00597, 20.00597, 20.00597, 20.00597, 20.00595, 
    20.00596, 20.00593, 20.00593, 20.00593, 20.00593, 20.00594, 20.00595, 
    20.00595, 20.00596, 20.00597, 20.00595, 20.00601, 20.00597, 20.00591, 
    20.00592, 20.00593, 20.00592, 20.00595, 20.00594, 20.00597, 20.00597, 
    20.00598, 20.00597, 20.00597, 20.00596, 20.00596, 20.00594, 20.00593, 
    20.00592, 20.00592, 20.00594, 20.00595, 20.00597, 20.00597, 20.00598, 
    20.00595, 20.00596, 20.00595, 20.00597, 20.00594, 20.00596, 20.00593, 
    20.00593, 20.00594, 20.00596, 20.00596, 20.00597, 20.00597, 20.00595, 
    20.00595, 20.00594, 20.00594, 20.00593, 20.00593, 20.00593, 20.00594, 
    20.00595, 20.00597, 20.00598, 20.00599, 20.006, 20.00599, 20.00601, 
    20.00599, 20.00603, 20.00596, 20.00599, 20.00594, 20.00595, 20.00596, 
    20.00598, 20.00597, 20.00598, 20.00595, 20.00594, 20.00593, 20.00592, 
    20.00593, 20.00593, 20.00594, 20.00594, 20.00595, 20.00594, 20.00597, 
    20.00598, 20.00601, 20.00603, 20.00604, 20.00605, 20.00606, 20.00606,
  20.00534, 20.00536, 20.00535, 20.00537, 20.00536, 20.00537, 20.00534, 
    20.00536, 20.00535, 20.00534, 20.0054, 20.00537, 20.00543, 20.00541, 
    20.00546, 20.00543, 20.00547, 20.00546, 20.00549, 20.00548, 20.00551, 
    20.00549, 20.00552, 20.0055, 20.00551, 20.00549, 20.00538, 20.0054, 
    20.00537, 20.00538, 20.00538, 20.00536, 20.00535, 20.00533, 20.00534, 
    20.00535, 20.00538, 20.00537, 20.00539, 20.00539, 20.00542, 20.00541, 
    20.00546, 20.00544, 20.00548, 20.00547, 20.00548, 20.00548, 20.00548, 
    20.00546, 20.00547, 20.00546, 20.00541, 20.00542, 20.00538, 20.00536, 
    20.00534, 20.00533, 20.00533, 20.00533, 20.00535, 20.00537, 20.00538, 
    20.00539, 20.00539, 20.00542, 20.00543, 20.00546, 20.00545, 20.00546, 
    20.00547, 20.00548, 20.00548, 20.00549, 20.00546, 20.00548, 20.00545, 
    20.00546, 20.0054, 20.00537, 20.00536, 20.00535, 20.00533, 20.00535, 
    20.00534, 20.00536, 20.00536, 20.00536, 20.00539, 20.00538, 20.00543, 
    20.00541, 20.00547, 20.00545, 20.00547, 20.00546, 20.00548, 20.00546, 
    20.00549, 20.00549, 20.00549, 20.0055, 20.00546, 20.00548, 20.00536, 
    20.00536, 20.00536, 20.00535, 20.00535, 20.00533, 20.00535, 20.00535, 
    20.00537, 20.00537, 20.00538, 20.0054, 20.00541, 20.00544, 20.00546, 
    20.00547, 20.00546, 20.00546, 20.00546, 20.00546, 20.00549, 20.00547, 
    20.0055, 20.0055, 20.00549, 20.0055, 20.00536, 20.00536, 20.00534, 
    20.00535, 20.00533, 20.00534, 20.00535, 20.00538, 20.00538, 20.00539, 
    20.0054, 20.00541, 20.00543, 20.00545, 20.00547, 20.00547, 20.00547, 
    20.00547, 20.00546, 20.00547, 20.00548, 20.00547, 20.0055, 20.00549, 
    20.0055, 20.0055, 20.00536, 20.00537, 20.00536, 20.00537, 20.00536, 
    20.00538, 20.00539, 20.00542, 20.00541, 20.00543, 20.00541, 20.00541, 
    20.00543, 20.00541, 20.00545, 20.00542, 20.00547, 20.00545, 20.00547, 
    20.00547, 20.00548, 20.00548, 20.00549, 20.00551, 20.00551, 20.00552, 
    20.00537, 20.00538, 20.00538, 20.00539, 20.0054, 20.00541, 20.00544, 
    20.00543, 20.00545, 20.00545, 20.00542, 20.00544, 20.00539, 20.0054, 
    20.00539, 20.00538, 20.00543, 20.0054, 20.00546, 20.00544, 20.00548, 
    20.00546, 20.0055, 20.00552, 20.00554, 20.00556, 20.00539, 20.00538, 
    20.00539, 20.00541, 20.00542, 20.00544, 20.00544, 20.00545, 20.00546, 
    20.00546, 20.00545, 20.00546, 20.0054, 20.00543, 20.00538, 20.0054, 
    20.00541, 20.0054, 20.00543, 20.00543, 20.00546, 20.00545, 20.00552, 
    20.00549, 20.00558, 20.00555, 20.00538, 20.00539, 20.00542, 20.0054, 
    20.00544, 20.00545, 20.00546, 20.00547, 20.00547, 20.00547, 20.00546, 
    20.00547, 20.00544, 20.00546, 20.00541, 20.00542, 20.00542, 20.00541, 
    20.00543, 20.00545, 20.00545, 20.00545, 20.00547, 20.00544, 20.00552, 
    20.00547, 20.0054, 20.00541, 20.00541, 20.00541, 20.00545, 20.00544, 
    20.00547, 20.00546, 20.00548, 20.00547, 20.00547, 20.00546, 20.00545, 
    20.00544, 20.00542, 20.00541, 20.00541, 20.00542, 20.00545, 20.00547, 
    20.00546, 20.00548, 20.00544, 20.00546, 20.00545, 20.00547, 20.00543, 
    20.00546, 20.00542, 20.00542, 20.00543, 20.00546, 20.00546, 20.00547, 
    20.00546, 20.00545, 20.00545, 20.00543, 20.00543, 20.00542, 20.00541, 
    20.00542, 20.00543, 20.00545, 20.00547, 20.00549, 20.00549, 20.00551, 
    20.00549, 20.00552, 20.0055, 20.00554, 20.00546, 20.0055, 20.00544, 
    20.00544, 20.00545, 20.00548, 20.00547, 20.00548, 20.00545, 20.00543, 
    20.00542, 20.00541, 20.00542, 20.00542, 20.00543, 20.00543, 20.00545, 
    20.00544, 20.00547, 20.00548, 20.00552, 20.00554, 20.00556, 20.00557, 
    20.00558, 20.00558,
  20.00503, 20.00505, 20.00505, 20.00507, 20.00506, 20.00507, 20.00504, 
    20.00505, 20.00504, 20.00503, 20.0051, 20.00507, 20.00514, 20.00512, 
    20.00517, 20.00513, 20.00518, 20.00517, 20.00519, 20.00519, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00522, 20.0052, 20.00507, 20.0051, 
    20.00507, 20.00508, 20.00508, 20.00506, 20.00505, 20.00503, 20.00503, 
    20.00505, 20.00508, 20.00507, 20.00509, 20.00509, 20.00512, 20.00511, 
    20.00516, 20.00515, 20.00519, 20.00518, 20.00519, 20.00518, 20.00519, 
    20.00517, 20.00518, 20.00517, 20.00511, 20.00513, 20.00508, 20.00505, 
    20.00504, 20.00502, 20.00502, 20.00503, 20.00505, 20.00506, 20.00508, 
    20.00508, 20.00509, 20.00512, 20.00513, 20.00516, 20.00516, 20.00517, 
    20.00517, 20.00519, 20.00519, 20.00519, 20.00517, 20.00518, 20.00515, 
    20.00516, 20.0051, 20.00507, 20.00506, 20.00505, 20.00503, 20.00504, 
    20.00504, 20.00505, 20.00506, 20.00506, 20.00508, 20.00507, 20.00513, 
    20.00511, 20.00517, 20.00516, 20.00518, 20.00517, 20.00519, 20.00517, 
    20.0052, 20.0052, 20.0052, 20.00521, 20.00517, 20.00519, 20.00506, 
    20.00506, 20.00506, 20.00504, 20.00504, 20.00503, 20.00504, 20.00505, 
    20.00506, 20.00507, 20.00508, 20.00509, 20.00511, 20.00514, 20.00516, 
    20.00517, 20.00517, 20.00517, 20.00516, 20.00516, 20.0052, 20.00518, 
    20.00521, 20.00521, 20.00519, 20.00521, 20.00506, 20.00505, 20.00504, 
    20.00505, 20.00503, 20.00504, 20.00505, 20.00507, 20.00508, 20.00508, 
    20.0051, 20.00511, 20.00513, 20.00516, 20.00518, 20.00517, 20.00517, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00518, 20.00521, 20.0052, 
    20.00521, 20.0052, 20.00505, 20.00506, 20.00506, 20.00507, 20.00506, 
    20.00508, 20.00509, 20.00512, 20.00511, 20.00513, 20.00511, 20.00512, 
    20.00513, 20.00511, 20.00516, 20.00513, 20.00518, 20.00515, 20.00518, 
    20.00518, 20.00518, 20.00519, 20.0052, 20.00522, 20.00522, 20.00523, 
    20.00507, 20.00508, 20.00508, 20.00509, 20.0051, 20.00512, 20.00514, 
    20.00513, 20.00515, 20.00515, 20.00513, 20.00514, 20.00509, 20.0051, 
    20.00509, 20.00507, 20.00513, 20.0051, 20.00516, 20.00514, 20.00519, 
    20.00517, 20.00521, 20.00524, 20.00525, 20.00528, 20.00509, 20.00508, 
    20.00509, 20.00511, 20.00512, 20.00514, 20.00515, 20.00515, 20.00516, 
    20.00517, 20.00515, 20.00517, 20.0051, 20.00514, 20.00508, 20.0051, 
    20.00511, 20.0051, 20.00513, 20.00514, 20.00516, 20.00515, 20.00523, 
    20.0052, 20.00529, 20.00527, 20.00508, 20.00509, 20.00512, 20.0051, 
    20.00515, 20.00516, 20.00516, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00518, 20.00514, 20.00516, 20.00512, 20.00513, 20.00512, 20.00512, 
    20.00513, 20.00515, 20.00515, 20.00516, 20.00517, 20.00515, 20.00524, 
    20.00518, 20.0051, 20.00511, 20.00512, 20.00511, 20.00516, 20.00514, 
    20.00518, 20.00517, 20.00519, 20.00518, 20.00518, 20.00517, 20.00516, 
    20.00514, 20.00512, 20.00511, 20.00511, 20.00513, 20.00515, 20.00518, 
    20.00517, 20.00519, 20.00514, 20.00516, 20.00515, 20.00517, 20.00513, 
    20.00517, 20.00512, 20.00513, 20.00514, 20.00516, 20.00517, 20.00517, 
    20.00517, 20.00515, 20.00515, 20.00514, 20.00513, 20.00513, 20.00512, 
    20.00513, 20.00513, 20.00515, 20.00517, 20.00519, 20.0052, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00526, 20.00517, 20.00521, 20.00514, 
    20.00515, 20.00516, 20.00519, 20.00517, 20.00519, 20.00515, 20.00513, 
    20.00512, 20.00511, 20.00512, 20.00512, 20.00513, 20.00513, 20.00515, 
    20.00514, 20.00518, 20.00519, 20.00523, 20.00525, 20.00528, 20.00529, 
    20.00529, 20.00529,
  20.00479, 20.00481, 20.00481, 20.00483, 20.00482, 20.00483, 20.0048, 
    20.00481, 20.0048, 20.00479, 20.00486, 20.00483, 20.0049, 20.00488, 
    20.00493, 20.0049, 20.00494, 20.00493, 20.00496, 20.00495, 20.00498, 
    20.00496, 20.005, 20.00498, 20.00498, 20.00496, 20.00484, 20.00486, 
    20.00484, 20.00484, 20.00484, 20.00482, 20.00481, 20.00479, 20.00479, 
    20.00481, 20.00484, 20.00483, 20.00486, 20.00485, 20.00488, 20.00487, 
    20.00492, 20.00491, 20.00495, 20.00494, 20.00495, 20.00495, 20.00495, 
    20.00493, 20.00494, 20.00493, 20.00488, 20.00489, 20.00484, 20.00482, 
    20.0048, 20.00478, 20.00479, 20.00479, 20.00481, 20.00482, 20.00484, 
    20.00485, 20.00485, 20.00488, 20.00489, 20.00493, 20.00492, 20.00493, 
    20.00494, 20.00495, 20.00495, 20.00496, 20.00493, 20.00495, 20.00492, 
    20.00493, 20.00486, 20.00483, 20.00482, 20.00481, 20.00479, 20.0048, 
    20.0048, 20.00481, 20.00482, 20.00482, 20.00485, 20.00484, 20.0049, 
    20.00487, 20.00494, 20.00492, 20.00494, 20.00493, 20.00495, 20.00493, 
    20.00496, 20.00497, 20.00496, 20.00498, 20.00493, 20.00495, 20.00482, 
    20.00482, 20.00482, 20.0048, 20.0048, 20.00479, 20.0048, 20.00481, 
    20.00482, 20.00483, 20.00484, 20.00486, 20.00488, 20.0049, 20.00492, 
    20.00494, 20.00493, 20.00493, 20.00493, 20.00492, 20.00496, 20.00494, 
    20.00498, 20.00497, 20.00496, 20.00497, 20.00482, 20.00481, 20.0048, 
    20.00481, 20.00479, 20.0048, 20.00481, 20.00484, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00492, 20.00494, 20.00494, 20.00494, 
    20.00494, 20.00493, 20.00495, 20.00495, 20.00494, 20.00497, 20.00496, 
    20.00497, 20.00497, 20.00481, 20.00482, 20.00482, 20.00483, 20.00482, 
    20.00484, 20.00485, 20.00489, 20.00487, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00488, 20.00492, 20.00489, 20.00494, 20.00492, 20.00495, 
    20.00494, 20.00495, 20.00496, 20.00497, 20.00499, 20.00498, 20.005, 
    20.00483, 20.00484, 20.00484, 20.00485, 20.00486, 20.00488, 20.0049, 
    20.00489, 20.00491, 20.00492, 20.00489, 20.00491, 20.00485, 20.00486, 
    20.00485, 20.00484, 20.0049, 20.00487, 20.00492, 20.00491, 20.00496, 
    20.00493, 20.00498, 20.005, 20.00502, 20.00504, 20.00485, 20.00484, 
    20.00485, 20.00487, 20.00489, 20.00491, 20.00491, 20.00491, 20.00492, 
    20.00493, 20.00491, 20.00493, 20.00486, 20.0049, 20.00484, 20.00486, 
    20.00487, 20.00487, 20.00489, 20.0049, 20.00493, 20.00491, 20.005, 
    20.00496, 20.00506, 20.00503, 20.00484, 20.00485, 20.00488, 20.00487, 
    20.00491, 20.00492, 20.00493, 20.00494, 20.00494, 20.00495, 20.00494, 
    20.00495, 20.00491, 20.00492, 20.00488, 20.00489, 20.00488, 20.00488, 
    20.0049, 20.00492, 20.00492, 20.00492, 20.00494, 20.00491, 20.005, 
    20.00494, 20.00486, 20.00488, 20.00488, 20.00487, 20.00492, 20.0049, 
    20.00495, 20.00493, 20.00495, 20.00494, 20.00494, 20.00493, 20.00492, 
    20.0049, 20.00489, 20.00487, 20.00488, 20.00489, 20.00492, 20.00494, 
    20.00493, 20.00495, 20.00491, 20.00492, 20.00492, 20.00494, 20.00489, 
    20.00493, 20.00488, 20.00489, 20.0049, 20.00493, 20.00493, 20.00494, 
    20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 20.00489, 20.00488, 
    20.00489, 20.00489, 20.00492, 20.00494, 20.00496, 20.00496, 20.00499, 
    20.00497, 20.005, 20.00497, 20.00502, 20.00493, 20.00497, 20.0049, 
    20.00491, 20.00492, 20.00495, 20.00494, 20.00496, 20.00491, 20.00489, 
    20.00488, 20.00487, 20.00488, 20.00488, 20.00489, 20.00489, 20.00492, 
    20.0049, 20.00494, 20.00496, 20.005, 20.00502, 20.00505, 20.00506, 
    20.00506, 20.00506,
  20.00426, 20.00427, 20.00427, 20.00429, 20.00428, 20.00429, 20.00426, 
    20.00428, 20.00426, 20.00426, 20.00432, 20.00429, 20.00435, 20.00433, 
    20.00438, 20.00435, 20.00438, 20.00438, 20.0044, 20.00439, 20.00442, 
    20.0044, 20.00444, 20.00442, 20.00442, 20.0044, 20.00429, 20.00431, 
    20.00429, 20.0043, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00427, 20.0043, 20.00429, 20.00431, 20.00431, 20.00434, 20.00433, 
    20.00437, 20.00436, 20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 
    20.00438, 20.00439, 20.00437, 20.00433, 20.00434, 20.0043, 20.00428, 
    20.00426, 20.00425, 20.00425, 20.00425, 20.00427, 20.00428, 20.0043, 
    20.0043, 20.00431, 20.00433, 20.00434, 20.00437, 20.00437, 20.00438, 
    20.00438, 20.0044, 20.00439, 20.0044, 20.00438, 20.00439, 20.00437, 
    20.00437, 20.00431, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00426, 20.00427, 20.00428, 20.00428, 20.0043, 20.00429, 20.00435, 
    20.00432, 20.00438, 20.00437, 20.00439, 20.00438, 20.00439, 20.00438, 
    20.0044, 20.00441, 20.00441, 20.00442, 20.00438, 20.00439, 20.00428, 
    20.00428, 20.00428, 20.00427, 20.00427, 20.00425, 20.00426, 20.00427, 
    20.00428, 20.00429, 20.0043, 20.00431, 20.00433, 20.00435, 20.00437, 
    20.00438, 20.00437, 20.00438, 20.00437, 20.00437, 20.00441, 20.00439, 
    20.00442, 20.00442, 20.0044, 20.00442, 20.00428, 20.00427, 20.00426, 
    20.00427, 20.00425, 20.00426, 20.00427, 20.00429, 20.0043, 20.0043, 
    20.00431, 20.00433, 20.00435, 20.00437, 20.00438, 20.00438, 20.00438, 
    20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 20.00442, 20.00441, 
    20.00442, 20.00441, 20.00428, 20.00428, 20.00428, 20.00429, 20.00428, 
    20.0043, 20.00431, 20.00434, 20.00433, 20.00434, 20.00433, 20.00433, 
    20.00434, 20.00433, 20.00437, 20.00434, 20.00439, 20.00436, 20.00439, 
    20.00438, 20.00439, 20.0044, 20.00441, 20.00443, 20.00442, 20.00444, 
    20.00429, 20.0043, 20.0043, 20.00431, 20.00432, 20.00433, 20.00435, 
    20.00434, 20.00436, 20.00436, 20.00434, 20.00435, 20.00431, 20.00431, 
    20.00431, 20.00429, 20.00435, 20.00432, 20.00437, 20.00435, 20.0044, 
    20.00438, 20.00442, 20.00444, 20.00446, 20.00448, 20.0043, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00436, 20.00436, 20.00436, 20.00437, 
    20.00438, 20.00436, 20.00438, 20.00432, 20.00435, 20.0043, 20.00431, 
    20.00432, 20.00432, 20.00434, 20.00435, 20.00437, 20.00436, 20.00443, 
    20.0044, 20.00449, 20.00447, 20.0043, 20.0043, 20.00433, 20.00432, 
    20.00436, 20.00437, 20.00437, 20.00438, 20.00438, 20.00439, 20.00438, 
    20.00439, 20.00436, 20.00437, 20.00433, 20.00434, 20.00434, 20.00433, 
    20.00435, 20.00436, 20.00436, 20.00437, 20.00438, 20.00436, 20.00444, 
    20.00439, 20.00431, 20.00433, 20.00433, 20.00433, 20.00437, 20.00435, 
    20.00439, 20.00438, 20.0044, 20.00439, 20.00439, 20.00438, 20.00437, 
    20.00435, 20.00434, 20.00433, 20.00433, 20.00434, 20.00436, 20.00438, 
    20.00438, 20.0044, 20.00435, 20.00437, 20.00437, 20.00438, 20.00434, 
    20.00438, 20.00434, 20.00434, 20.00435, 20.00437, 20.00438, 20.00438, 
    20.00438, 20.00436, 20.00436, 20.00435, 20.00435, 20.00434, 20.00433, 
    20.00434, 20.00434, 20.00436, 20.00438, 20.0044, 20.0044, 20.00443, 
    20.00441, 20.00444, 20.00441, 20.00446, 20.00438, 20.00441, 20.00435, 
    20.00436, 20.00437, 20.0044, 20.00438, 20.0044, 20.00436, 20.00434, 
    20.00434, 20.00433, 20.00434, 20.00434, 20.00434, 20.00434, 20.00436, 
    20.00435, 20.00439, 20.0044, 20.00443, 20.00446, 20.00448, 20.00449, 
    20.00449, 20.00449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258142, 0.5258147, 0.5258146, 0.525815, 0.5258148, 0.5258151, 0.5258143, 
    0.5258147, 0.5258144, 0.5258142, 0.5258159, 0.5258151, 0.5258167, 
    0.5258162, 0.5258176, 0.5258167, 0.5258178, 0.5258175, 0.5258182, 
    0.525818, 0.5258188, 0.5258182, 0.5258192, 0.5258186, 0.5258187, 
    0.5258182, 0.5258152, 0.5258158, 0.5258152, 0.5258152, 0.5258152, 
    0.5258148, 0.5258146, 0.5258141, 0.5258142, 0.5258145, 0.5258153, 
    0.5258151, 0.5258157, 0.5258157, 0.5258164, 0.5258161, 0.5258173, 
    0.525817, 0.525818, 0.5258178, 0.525818, 0.5258179, 0.525818, 0.5258176, 
    0.5258178, 0.5258175, 0.5258161, 0.5258165, 0.5258154, 0.5258147, 
    0.5258143, 0.525814, 0.525814, 0.5258141, 0.5258145, 0.525815, 0.5258152, 
    0.5258155, 0.5258157, 0.5258163, 0.5258167, 0.5258174, 0.5258173, 
    0.5258175, 0.5258177, 0.525818, 0.525818, 0.5258182, 0.5258175, 
    0.5258179, 0.5258172, 0.5258174, 0.5258157, 0.5258151, 0.5258148, 
    0.5258146, 0.5258141, 0.5258144, 0.5258143, 0.5258147, 0.5258149, 
    0.5258148, 0.5258155, 0.5258152, 0.5258167, 0.525816, 0.5258177, 
    0.5258173, 0.5258178, 0.5258175, 0.5258179, 0.5258176, 0.5258182, 
    0.5258184, 0.5258183, 0.5258186, 0.5258176, 0.525818, 0.5258148, 
    0.5258148, 0.5258149, 0.5258145, 0.5258145, 0.5258141, 0.5258144, 
    0.5258145, 0.5258149, 0.5258151, 0.5258153, 0.5258157, 0.5258162, 
    0.5258169, 0.5258173, 0.5258176, 0.5258175, 0.5258176, 0.5258174, 
    0.5258173, 0.5258183, 0.5258178, 0.5258186, 0.5258186, 0.5258182, 
    0.5258186, 0.5258148, 0.5258147, 0.5258143, 0.5258146, 0.5258141, 
    0.5258144, 0.5258145, 0.5258152, 0.5258154, 0.5258155, 0.5258158, 
    0.5258161, 0.5258167, 0.5258172, 0.5258177, 0.5258177, 0.5258177, 
    0.5258178, 0.5258175, 0.5258179, 0.5258179, 0.5258178, 0.5258185, 
    0.5258183, 0.5258186, 0.5258184, 0.5258147, 0.5258149, 0.5258148, 
    0.525815, 0.5258149, 0.5258154, 0.5258156, 0.5258164, 0.5258161, 
    0.5258166, 0.5258161, 0.5258163, 0.5258167, 0.5258162, 0.5258172, 
    0.5258165, 0.5258178, 0.5258171, 0.5258179, 0.5258177, 0.5258179, 
    0.5258181, 0.5258184, 0.5258188, 0.5258188, 0.5258191, 0.5258152, 
    0.5258154, 0.5258154, 0.5258157, 0.5258158, 0.5258162, 0.5258169, 
    0.5258166, 0.525817, 0.5258172, 0.5258165, 0.5258169, 0.5258156, 
    0.5258158, 0.5258157, 0.5258152, 0.5258167, 0.5258159, 0.5258173, 
    0.5258169, 0.5258181, 0.5258175, 0.5258187, 0.5258192, 0.5258197, 
    0.5258202, 0.5258155, 0.5258154, 0.5258157, 0.5258161, 0.5258164, 
    0.5258169, 0.525817, 0.5258171, 0.5258173, 0.5258175, 0.5258171, 
    0.5258176, 0.5258158, 0.5258167, 0.5258153, 0.5258157, 0.525816, 
    0.5258159, 0.5258166, 0.5258167, 0.5258174, 0.5258171, 0.5258191, 
    0.5258182, 0.5258206, 0.52582, 0.5258153, 0.5258155, 0.5258163, 0.525816, 
    0.525817, 0.5258172, 0.5258175, 0.5258177, 0.5258177, 0.5258179, 
    0.5258176, 0.5258179, 0.5258169, 0.5258173, 0.5258162, 0.5258165, 
    0.5258164, 0.5258162, 0.5258167, 0.5258171, 0.5258171, 0.5258173, 
    0.5258177, 0.525817, 0.5258192, 0.5258178, 0.5258158, 0.5258162, 
    0.5258163, 0.5258161, 0.5258172, 0.5258168, 0.5258179, 0.5258176, 
    0.525818, 0.5258178, 0.5258178, 0.5258175, 0.5258173, 0.5258168, 
    0.5258164, 0.5258161, 0.5258162, 0.5258166, 0.5258172, 0.5258177, 
    0.5258176, 0.525818, 0.5258169, 0.5258174, 0.5258172, 0.5258176, 
    0.5258166, 0.5258175, 0.5258164, 0.5258165, 0.5258168, 0.5258174, 
    0.5258175, 0.5258177, 0.5258176, 0.5258172, 0.5258171, 0.5258168, 
    0.5258167, 0.5258164, 0.5258163, 0.5258164, 0.5258166, 0.5258172, 
    0.5258176, 0.5258182, 0.5258183, 0.5258189, 0.5258184, 0.5258192, 
    0.5258185, 0.5258197, 0.5258176, 0.5258185, 0.5258168, 0.525817, 
    0.5258173, 0.525818, 0.5258176, 0.5258181, 0.5258171, 0.5258166, 
    0.5258164, 0.5258161, 0.5258164, 0.5258164, 0.5258166, 0.5258166, 
    0.5258172, 0.5258169, 0.5258178, 0.5258181, 0.5258191, 0.5258197, 
    0.5258203, 0.5258206, 0.5258206, 0.5258207 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  5.139921e-21, -5.139921e-21, -1.027984e-20, 1.541976e-20, 1.28498e-20, 
    -2.569961e-21, 1.798972e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 2.055969e-20, 1.027984e-20, -1.003089e-36, 2.569961e-20, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 0, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, 2.055969e-20, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, 
    1.003089e-36, -1.541976e-20, -2.569961e-21, 1.798972e-20, 2.569961e-21, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, 1.798972e-20, 1.541976e-20, 
    2.826957e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 1.003089e-36, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, 2.055969e-20, -1.027984e-20, 
    -1.027984e-20, -7.709882e-21, 1.541976e-20, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, 1.798972e-20, 0, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, -1.28498e-20, 1.28498e-20, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.798972e-20, 2.055969e-20, 5.139921e-21, 
    7.709882e-21, 7.709882e-21, -7.709882e-21, -1.28498e-20, -1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -1.027984e-20, -1.798972e-20, 1.541976e-20, 1.28498e-20, 1.28498e-20, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -1.027984e-20, 1.28498e-20, 2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -5.139921e-21, 2.569961e-21, 0, -5.139921e-21, -2.569961e-21, 
    1.541976e-20, -1.28498e-20, -1.003089e-36, -5.139921e-21, 1.798972e-20, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, 0, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, -1.541976e-20, 1.28498e-20, -1.798972e-20, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, 1.003089e-36, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 1.003089e-36, -2.569961e-21, 
    0, -1.027984e-20, -1.28498e-20, -1.28498e-20, 1.003089e-36, 
    -5.139921e-21, -1.003089e-36, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, 1.28498e-20, 1.027984e-20, 
    -1.28498e-20, 0, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -7.709882e-21, -2.312965e-20, 2.569961e-21, -1.541976e-20, 2.312965e-20, 
    -1.003089e-36, -2.569961e-20, 1.027984e-20, -1.027984e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 7.709882e-21, 1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, 1.798972e-20, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -1.003089e-36, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -1.003089e-36, -1.28498e-20, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 1.003089e-36, 7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -3.083953e-20, 5.139921e-21, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -1.28498e-20, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    -1.28498e-20, -7.709882e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -2.569961e-21, 5.139921e-21, 2.312965e-20, -2.312965e-20, 1.541976e-20, 
    -1.541976e-20, -5.139921e-21, -1.541976e-20, -1.28498e-20, -7.709882e-21, 
    1.003089e-36, 1.28498e-20, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, 0, 
    2.569961e-21, -2.569961e-21, -1.798972e-20, 1.28498e-20, 0, 2.055969e-20, 
    7.709882e-21, 2.569961e-20, 1.027984e-20, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.027984e-20, -1.003089e-36, -5.139921e-21, 
    -1.798972e-20, 1.28498e-20, -5.139921e-21, 2.569961e-21, 1.28498e-20, 
    7.709882e-21, -1.027984e-20, 1.027984e-20, 1.28498e-20, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 2.569961e-20, -1.541976e-20, 1.003089e-36, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -1.003089e-36, 0, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, 2.055969e-20, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 1.003089e-36, -1.003089e-36, -1.027984e-20, -1.798972e-20, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, -7.709882e-21, 1.003089e-36, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, 
    0, -5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    1.798972e-20, -5.139921e-21, -7.709882e-21, -7.709882e-21, 1.003089e-36, 
    1.027984e-20, -1.28498e-20, 2.055969e-20, 2.569961e-21, -5.139921e-21, 0, 
    -1.28498e-20, -2.569961e-21, 2.055969e-20, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -2.569961e-21, 1.541976e-20, 0, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21,
  1.027984e-20, 1.003089e-36, 1.003089e-36, -2.569961e-21, -2.569961e-21, 0, 
    1.003089e-36, -1.541976e-20, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    1.027984e-20, 0, 2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -1.003089e-36, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 0, -2.569961e-21, -7.709882e-21, 1.541976e-20, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 0, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -1.541976e-20, 0, -5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 0, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -2.055969e-20, -5.139921e-21, 0, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, 0, 5.139921e-21, 
    -7.709882e-21, 1.027984e-20, 0, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    0, -1.28498e-20, -1.027984e-20, -2.569961e-21, 0, -1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 0, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, -7.709882e-21, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, -1.798972e-20, 
    7.709882e-21, 2.569961e-21, -1.541976e-20, -1.28498e-20, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, 0, 0, 7.709882e-21, 
    -2.569961e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -1.28498e-20, -2.569961e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, 0, 2.569961e-21, -5.139921e-21, 1.28498e-20, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, 1.541976e-20, 0, 1.003089e-36, 
    2.569961e-21, 1.541976e-20, 0, 1.28498e-20, -1.28498e-20, 0, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, 7.709882e-21, 0, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 1.798972e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, -1.28498e-20, 0, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    7.709882e-21, 1.003089e-36, 5.139921e-21, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, 0, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, 0, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, 1.798972e-20, -5.139921e-21, 
    1.28498e-20, 7.709882e-21, -1.28498e-20, 0, 5.139921e-21, 2.569961e-21, 
    -1.541976e-20, -2.569961e-21, 1.28498e-20, -5.139921e-21, 0, 
    1.798972e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -5.139921e-21, 0, -1.28498e-20, 1.28498e-20, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 0, 1.541976e-20, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, -1.027984e-20, 
    0, -5.139921e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, 0, 0, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, -1.28498e-20, 0, -1.027984e-20, 
    -7.709882e-21, 7.709882e-21, 5.139921e-21, 1.798972e-20, 1.003089e-36, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.28498e-20, -1.28498e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -1.798972e-20, 1.003089e-36, 
    -7.709882e-21, -1.027984e-20, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    -7.709882e-21, -2.569961e-21, 1.28498e-20, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, 0, 1.541976e-20, -1.027984e-20, 7.709882e-21, 1.027984e-20, 
    5.139921e-21, 0, 2.055969e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 1.003089e-36, 
    0, -2.569961e-21, 1.027984e-20, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, 0, -7.709882e-21, 1.027984e-20, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 5.139921e-21, 2.569961e-21,
  -5.139921e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    0, 5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    -1.003089e-36, -2.312965e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, 5.139921e-21, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 0, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, -2.055969e-20, -1.003089e-36, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, -1.798972e-20, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, -1.541976e-20, 
    -2.569961e-21, -1.28498e-20, -1.003089e-36, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 1.541976e-20, 0, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 7.709882e-21, -1.798972e-20, 
    0, 2.569961e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 2.055969e-20, -7.709882e-21, -1.28498e-20, -1.003089e-36, 
    -1.28498e-20, 7.709882e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, -1.003089e-36, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, 1.027984e-20, 
    1.541976e-20, -1.027984e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    0, 5.139921e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 0, 
    -5.139921e-21, 0, 7.709882e-21, 7.709882e-21, -2.569961e-21, 
    -1.798972e-20, 0, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -1.28498e-20, -2.569961e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 
    2.569961e-21, -1.027984e-20, 1.027984e-20, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 1.541976e-20, 1.003089e-36, -5.139921e-21, 
    1.541976e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, 0, -1.28498e-20, 
    -1.541976e-20, 1.027984e-20, -1.28498e-20, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, 1.798972e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, -1.541976e-20, 2.569961e-21, 
    -2.569961e-21, 1.003089e-36, 5.139921e-21, -7.709882e-21, -1.28498e-20, 
    -1.541976e-20, -1.027984e-20, -2.569961e-21, 1.28498e-20, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.541976e-20, 
    -2.569961e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, -1.003089e-36, 
    2.569961e-21, 0, -5.139921e-21, 0, -2.569961e-21, 1.541976e-20, 
    2.055969e-20, 2.055969e-20, 1.003089e-36, 7.709882e-21, 1.541976e-20, 
    1.027984e-20, -1.541976e-20, 7.709882e-21, -1.28498e-20, -1.28498e-20, 
    7.709882e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.541976e-20, -2.569961e-21, 2.569961e-21, 
    -1.798972e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, -1.541976e-20, 
    -7.709882e-21, 1.027984e-20, 1.003089e-36, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, -1.28498e-20, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 0, -2.569961e-21, 0, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 0, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, -1.003089e-36, -2.055969e-20, 
    1.027984e-20, -1.003089e-36, 1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, 1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.027984e-20, 
    0, 5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    1.28498e-20, 2.569961e-21, -1.28498e-20, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.003089e-36, 1.541976e-20, -7.709882e-21, 0, 
    -7.709882e-21, 2.312965e-20, 7.709882e-21, 1.798972e-20, 0, 7.709882e-21, 
    0, -2.569961e-21, 0, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -1.003089e-36, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -1.027984e-20, 2.569961e-21, 1.28498e-20, 
    -7.709882e-21, 1.003089e-36, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.28498e-20, 2.569961e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    1.003089e-36, -1.003089e-36, 7.709882e-21, 1.027984e-20, -1.003089e-36,
  -7.709882e-21, 0, -2.569961e-21, 1.798972e-20, 1.003089e-36, 5.139921e-21, 
    -1.003089e-36, -7.709882e-21, -1.003089e-36, -1.28498e-20, 1.28498e-20, 
    5.139921e-21, 0, 2.569961e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 0, 
    5.139921e-21, -1.003089e-36, 1.541976e-20, 1.798972e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -1.541976e-20, 1.541976e-20, 2.569961e-21, 
    1.28498e-20, 1.28498e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -1.798972e-20, 7.709882e-21, 1.28498e-20, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 1.28498e-20, 5.139921e-21, -5.139921e-21, 0, 
    5.139921e-21, 1.541976e-20, -7.709882e-21, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.003089e-36, 5.139921e-21, -1.798972e-20, 
    -1.003089e-36, 1.027984e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -1.798972e-20, -2.569961e-21, -1.541976e-20, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, 1.541976e-20, 
    -1.28498e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 1.003089e-36, 
    -1.541976e-20, -1.28498e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, 1.798972e-20, -2.569961e-21, 0, -2.055969e-20, 
    2.055969e-20, 2.569961e-21, 1.027984e-20, 1.003089e-36, 1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, 1.541976e-20, 1.541976e-20, 
    1.798972e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -1.003089e-36, -2.569961e-21, -2.569961e-21, -7.709882e-21, 1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -1.027984e-20, 1.003089e-36, -5.139921e-21, 
    1.003089e-36, 2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, -1.003089e-36, -7.709882e-21, 1.003089e-36, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, 2.569961e-21, -1.798972e-20, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 1.003089e-36, 1.28498e-20, -2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 2.055969e-20, 2.569961e-21, 
    -5.139921e-21, 1.541976e-20, -1.003089e-36, 1.003089e-36, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, -1.003089e-36, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 1.027984e-20, 
    -1.798972e-20, 2.569961e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    1.027984e-20, 1.798972e-20, 1.027984e-20, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, 7.709882e-21, -1.28498e-20, 1.027984e-20, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    -1.003089e-36, 1.28498e-20, -1.027984e-20, 5.139921e-21, 2.055969e-20, 
    -1.28498e-20, 2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -1.027984e-20, -5.139921e-21, -1.798972e-20, 0, 2.569961e-21, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, 1.798972e-20, 2.569961e-21, -2.569961e-20, -1.541976e-20, 
    0, -2.569961e-21, 7.709882e-21, -1.027984e-20, -1.28498e-20, 
    5.139921e-21, 7.709882e-21, 0, 2.569961e-21, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    7.709882e-21, 2.569961e-21, 1.003089e-36, 7.709882e-21, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, 2.312965e-20, -2.569961e-21, 
    0, -1.28498e-20, 1.28498e-20, -2.569961e-21, 1.28498e-20, 5.139921e-21, 
    7.709882e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, 1.28498e-20, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -1.027984e-20, -1.28498e-20, 
    1.28498e-20, 5.139921e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, 
    1.003089e-36, -5.139921e-21, 1.541976e-20, 1.28498e-20, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, -1.798972e-20, -7.709882e-21, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, -1.003089e-36, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    -2.055969e-20, 1.003089e-36, 5.139921e-21,
  7.709882e-21, -1.798972e-20, 1.28498e-20, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -1.003089e-36, 1.003089e-36, -1.28498e-20, -2.569961e-20, 
    1.28498e-20, -1.541976e-20, 1.28498e-20, -7.709882e-21, -2.569961e-21, 
    -2.826957e-20, 5.139921e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, 
    1.798972e-20, -1.003089e-36, -1.027984e-20, 7.709882e-21, -2.569961e-21, 
    0, -2.569961e-21, 2.569961e-21, 1.027984e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, -1.027984e-20, 1.28498e-20, 
    -5.139921e-21, 1.541976e-20, -2.055969e-20, 1.541976e-20, -1.798972e-20, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -1.28498e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    1.541976e-20, 2.569961e-21, -7.709882e-21, 1.28498e-20, 1.798972e-20, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 
    7.709882e-21, 2.569961e-21, -1.541976e-20, 2.312965e-20, -5.139921e-21, 
    -2.055969e-20, -7.709882e-21, 1.28498e-20, 5.139921e-21, -1.541976e-20, 
    7.709882e-21, -1.28498e-20, -2.055969e-20, -2.569961e-21, -2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 0, -1.798972e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 1.541976e-20, 
    -2.055969e-20, 7.709882e-21, 1.541976e-20, 2.055969e-20, -3.083953e-20, 
    -2.569961e-21, 1.541976e-20, 2.055969e-20, 1.003089e-36, 1.541976e-20, 
    2.569961e-20, 5.139921e-21, 2.569961e-21, -1.003089e-36, 1.003089e-36, 
    -1.541976e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 1.28498e-20, 
    1.28498e-20, -5.139921e-21, 3.009266e-36, -2.569961e-20, 1.003089e-36, 
    1.027984e-20, -2.569961e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 1.541976e-20, -7.709882e-21, -1.28498e-20, 7.709882e-21, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, 2.569961e-21, -7.709882e-21, -1.003089e-36, 5.139921e-21, 
    -5.139921e-21, -1.003089e-36, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -1.28498e-20, 5.139921e-21, -7.709882e-21, 2.312965e-20, -1.003089e-36, 
    -2.569961e-21, -1.28498e-20, 2.569961e-21, -2.312965e-20, -2.569961e-21, 
    7.709882e-21, -1.003089e-36, 5.139921e-21, 1.798972e-20, -1.003089e-36, 
    2.569961e-20, 7.709882e-21, -1.027984e-20, 1.541976e-20, -2.312965e-20, 
    -1.541976e-20, -1.28498e-20, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    2.569961e-21, 0, 5.139921e-21, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -1.798972e-20, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.798972e-20, 1.28498e-20, 1.027984e-20, 
    1.28498e-20, 5.139921e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    1.798972e-20, 1.027984e-20, -2.569961e-21, 1.28498e-20, -2.055969e-20, 
    1.798972e-20, -2.569961e-21, -2.055969e-20, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, -1.541976e-20, -1.027984e-20, 
    1.798972e-20, 2.569961e-21, 1.003089e-36, 1.28498e-20, -2.569961e-21, 
    7.709882e-21, -5.139921e-21, -1.28498e-20, -2.055969e-20, 1.798972e-20, 
    0, 2.569961e-21, -7.709882e-21, 1.003089e-36, -2.055969e-20, 
    1.027984e-20, -7.709882e-21, -1.28498e-20, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 1.541976e-20, 
    1.541976e-20, 1.28498e-20, -2.569961e-21, 0, -5.139921e-21, 1.798972e-20, 
    -2.569961e-21, -1.28498e-20, -2.569961e-21, -1.003089e-36, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    2.569961e-21, 0, 2.569961e-21, 7.709882e-21, -7.709882e-21, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, -7.709882e-21, -5.139921e-21, 1.541976e-20, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, -1.027984e-20, 1.541976e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, 1.027984e-20, 1.28498e-20, 7.709882e-21, 
    7.709882e-21, 5.139921e-21, 1.798972e-20, -2.569961e-21, -1.798972e-20, 
    -1.541976e-20, 1.027984e-20, -1.541976e-20, -1.003089e-36, -2.569961e-21, 
    -1.28498e-20, 1.28498e-20, -7.709882e-21, 5.139921e-21, 1.28498e-20, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 1.003089e-36, -1.798972e-20, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, 1.798972e-20, 
    2.312965e-20, -7.709882e-21, 7.709882e-21, -1.003089e-36, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, 1.798972e-20, 1.027984e-20, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, -5.139921e-21, 
    2.312965e-20, -7.709882e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -2.312965e-20, 1.027984e-20, -1.027984e-20, 1.28498e-20, -7.709882e-21, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, 
    1.003089e-36, 2.569961e-21,
  6.259378e-29, 6.259384e-29, 6.259383e-29, 6.259388e-29, 6.259385e-29, 
    6.259388e-29, 6.259379e-29, 6.259384e-29, 6.259381e-29, 6.259378e-29, 
    6.259398e-29, 6.259388e-29, 6.259407e-29, 6.259401e-29, 6.259417e-29, 
    6.259407e-29, 6.259419e-29, 6.259416e-29, 6.259423e-29, 6.259421e-29, 
    6.25943e-29, 6.259424e-29, 6.259435e-29, 6.259429e-29, 6.25943e-29, 
    6.259424e-29, 6.25939e-29, 6.259396e-29, 6.25939e-29, 6.25939e-29, 
    6.25939e-29, 6.259385e-29, 6.259382e-29, 6.259377e-29, 6.259378e-29, 
    6.259382e-29, 6.259391e-29, 6.259388e-29, 6.259395e-29, 6.259395e-29, 
    6.259404e-29, 6.2594e-29, 6.259414e-29, 6.25941e-29, 6.259422e-29, 
    6.259419e-29, 6.259421e-29, 6.25942e-29, 6.259421e-29, 6.259417e-29, 
    6.259419e-29, 6.259415e-29, 6.259401e-29, 6.259405e-29, 6.259392e-29, 
    6.259384e-29, 6.259379e-29, 6.259376e-29, 6.259376e-29, 6.259377e-29, 
    6.259382e-29, 6.259387e-29, 6.25939e-29, 6.259393e-29, 6.259395e-29, 
    6.259402e-29, 6.259406e-29, 6.259414e-29, 6.259413e-29, 6.259416e-29, 
    6.259418e-29, 6.259422e-29, 6.259422e-29, 6.259423e-29, 6.259416e-29, 
    6.259421e-29, 6.259412e-29, 6.259414e-29, 6.259396e-29, 6.259388e-29, 
    6.259385e-29, 6.259383e-29, 6.259376e-29, 6.259381e-29, 6.259379e-29, 
    6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259393e-29, 6.25939e-29, 
    6.259407e-29, 6.259399e-29, 6.259418e-29, 6.259413e-29, 6.259419e-29, 
    6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259424e-29, 6.259426e-29, 
    6.259425e-29, 6.259429e-29, 6.259416e-29, 6.259421e-29, 6.259385e-29, 
    6.259385e-29, 6.259386e-29, 6.259381e-29, 6.259381e-29, 6.259377e-29, 
    6.259381e-29, 6.259382e-29, 6.259386e-29, 6.259388e-29, 6.259391e-29, 
    6.259396e-29, 6.259401e-29, 6.259408e-29, 6.259414e-29, 6.259417e-29, 
    6.259415e-29, 6.259417e-29, 6.259415e-29, 6.259414e-29, 6.259425e-29, 
    6.259419e-29, 6.259428e-29, 6.259428e-29, 6.259423e-29, 6.259428e-29, 
    6.259385e-29, 6.259384e-29, 6.259379e-29, 6.259383e-29, 6.259377e-29, 
    6.25938e-29, 6.259382e-29, 6.25939e-29, 6.259391e-29, 6.259393e-29, 
    6.259396e-29, 6.2594e-29, 6.259407e-29, 6.259413e-29, 6.259419e-29, 
    6.259418e-29, 6.259418e-29, 6.259419e-29, 6.259416e-29, 6.25942e-29, 
    6.25942e-29, 6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259428e-29, 
    6.259426e-29, 6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259387e-29, 
    6.259386e-29, 6.259393e-29, 6.259394e-29, 6.259404e-29, 6.2594e-29, 
    6.259406e-29, 6.259401e-29, 6.259402e-29, 6.259406e-29, 6.259401e-29, 
    6.259413e-29, 6.259405e-29, 6.259419e-29, 6.259411e-29, 6.25942e-29, 
    6.259419e-29, 6.259421e-29, 6.259423e-29, 6.259426e-29, 6.259431e-29, 
    6.25943e-29, 6.259434e-29, 6.25939e-29, 6.259392e-29, 6.259392e-29, 
    6.259394e-29, 6.259397e-29, 6.259401e-29, 6.259408e-29, 6.259406e-29, 
    6.259411e-29, 6.259412e-29, 6.259404e-29, 6.259409e-29, 6.259394e-29, 
    6.259396e-29, 6.259395e-29, 6.25939e-29, 6.259407e-29, 6.259398e-29, 
    6.259414e-29, 6.259409e-29, 6.259423e-29, 6.259416e-29, 6.259429e-29, 
    6.259435e-29, 6.25944e-29, 6.259447e-29, 6.259393e-29, 6.259391e-29, 
    6.259395e-29, 6.259399e-29, 6.259404e-29, 6.25941e-29, 6.25941e-29, 
    6.259411e-29, 6.259414e-29, 6.259416e-29, 6.259411e-29, 6.259417e-29, 
    6.259397e-29, 6.259407e-29, 6.259391e-29, 6.259396e-29, 6.259399e-29, 
    6.259398e-29, 6.259405e-29, 6.259407e-29, 6.259415e-29, 6.259411e-29, 
    6.259434e-29, 6.259423e-29, 6.259452e-29, 6.259444e-29, 6.259391e-29, 
    6.259393e-29, 6.259402e-29, 6.259398e-29, 6.25941e-29, 6.259413e-29, 
    6.259415e-29, 6.259418e-29, 6.259419e-29, 6.25942e-29, 6.259417e-29, 
    6.25942e-29, 6.25941e-29, 6.259414e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259401e-29, 6.259406e-29, 6.259411e-29, 6.259411e-29, 
    6.259413e-29, 6.259418e-29, 6.25941e-29, 6.259435e-29, 6.259419e-29, 
    6.259396e-29, 6.259401e-29, 6.259402e-29, 6.2594e-29, 6.259413e-29, 
    6.259408e-29, 6.25942e-29, 6.259417e-29, 6.259422e-29, 6.259419e-29, 
    6.259419e-29, 6.259416e-29, 6.259413e-29, 6.259408e-29, 6.259404e-29, 
    6.2594e-29, 6.259401e-29, 6.259405e-29, 6.259412e-29, 6.259419e-29, 
    6.259417e-29, 6.259422e-29, 6.259409e-29, 6.259414e-29, 6.259412e-29, 
    6.259417e-29, 6.259406e-29, 6.259416e-29, 6.259403e-29, 6.259404e-29, 
    6.259408e-29, 6.259414e-29, 6.259416e-29, 6.259418e-29, 6.259417e-29, 
    6.259412e-29, 6.259411e-29, 6.259408e-29, 6.259407e-29, 6.259404e-29, 
    6.259402e-29, 6.259404e-29, 6.259406e-29, 6.259412e-29, 6.259417e-29, 
    6.259423e-29, 6.259425e-29, 6.259431e-29, 6.259426e-29, 6.259435e-29, 
    6.259427e-29, 6.259441e-29, 6.259416e-29, 6.259427e-29, 6.259408e-29, 
    6.25941e-29, 6.259414e-29, 6.259422e-29, 6.259417e-29, 6.259423e-29, 
    6.259411e-29, 6.259405e-29, 6.259404e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259406e-29, 6.259405e-29, 6.259412e-29, 6.259408e-29, 
    6.259419e-29, 6.259423e-29, 6.259434e-29, 6.259441e-29, 6.259447e-29, 
    6.25945e-29, 6.259452e-29, 6.259452e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.13664e-10, 2.146069e-10, 2.144236e-10, 2.151841e-10, 2.147623e-10, 
    2.152603e-10, 2.138552e-10, 2.146443e-10, 2.141406e-10, 2.137489e-10, 
    2.166601e-10, 2.152181e-10, 2.181584e-10, 2.172386e-10, 2.195493e-10, 
    2.180152e-10, 2.198587e-10, 2.195051e-10, 2.205694e-10, 2.202645e-10, 
    2.216258e-10, 2.207102e-10, 2.223316e-10, 2.214072e-10, 2.215518e-10, 
    2.2068e-10, 2.155083e-10, 2.164806e-10, 2.154507e-10, 2.155894e-10, 
    2.155272e-10, 2.14771e-10, 2.143899e-10, 2.13592e-10, 2.137368e-10, 
    2.143229e-10, 2.156517e-10, 2.152007e-10, 2.163375e-10, 2.163118e-10, 
    2.175776e-10, 2.170069e-10, 2.191344e-10, 2.185297e-10, 2.202773e-10, 
    2.198378e-10, 2.202566e-10, 2.201296e-10, 2.202583e-10, 2.196137e-10, 
    2.198898e-10, 2.193227e-10, 2.171137e-10, 2.177629e-10, 2.158269e-10, 
    2.146628e-10, 2.138898e-10, 2.133412e-10, 2.134188e-10, 2.135666e-10, 
    2.143263e-10, 2.150407e-10, 2.155851e-10, 2.159493e-10, 2.163082e-10, 
    2.173943e-10, 2.179692e-10, 2.192567e-10, 2.190244e-10, 2.19418e-10, 
    2.19794e-10, 2.204254e-10, 2.203215e-10, 2.205996e-10, 2.194076e-10, 
    2.201998e-10, 2.188921e-10, 2.192497e-10, 2.164055e-10, 2.153223e-10, 
    2.148618e-10, 2.144589e-10, 2.134784e-10, 2.141555e-10, 2.138885e-10, 
    2.145236e-10, 2.149271e-10, 2.147275e-10, 2.159593e-10, 2.154804e-10, 
    2.180033e-10, 2.169166e-10, 2.197502e-10, 2.190721e-10, 2.199127e-10, 
    2.194838e-10, 2.202187e-10, 2.195573e-10, 2.207032e-10, 2.209527e-10, 
    2.207822e-10, 2.214372e-10, 2.195206e-10, 2.202566e-10, 2.147219e-10, 
    2.147545e-10, 2.149061e-10, 2.142395e-10, 2.141988e-10, 2.13588e-10, 
    2.141315e-10, 2.143629e-10, 2.149505e-10, 2.15298e-10, 2.156284e-10, 
    2.163549e-10, 2.171662e-10, 2.183008e-10, 2.19116e-10, 2.196625e-10, 
    2.193274e-10, 2.196232e-10, 2.192925e-10, 2.191375e-10, 2.208592e-10, 
    2.198924e-10, 2.21343e-10, 2.212627e-10, 2.206062e-10, 2.212718e-10, 
    2.147773e-10, 2.1459e-10, 2.139397e-10, 2.144487e-10, 2.135215e-10, 
    2.140404e-10, 2.143388e-10, 2.154904e-10, 2.157434e-10, 2.15978e-10, 
    2.164414e-10, 2.170361e-10, 2.180793e-10, 2.189871e-10, 2.198159e-10, 
    2.197552e-10, 2.197766e-10, 2.199617e-10, 2.195031e-10, 2.20037e-10, 
    2.201266e-10, 2.198923e-10, 2.21252e-10, 2.208635e-10, 2.21261e-10, 
    2.210081e-10, 2.146509e-10, 2.149661e-10, 2.147958e-10, 2.15116e-10, 
    2.148904e-10, 2.158936e-10, 2.161944e-10, 2.17602e-10, 2.170244e-10, 
    2.179438e-10, 2.171178e-10, 2.172641e-10, 2.179737e-10, 2.171624e-10, 
    2.18937e-10, 2.177338e-10, 2.199689e-10, 2.187672e-10, 2.200442e-10, 
    2.198123e-10, 2.201963e-10, 2.205401e-10, 2.209727e-10, 2.217709e-10, 
    2.21586e-10, 2.222536e-10, 2.154359e-10, 2.158447e-10, 2.158088e-10, 
    2.162366e-10, 2.16553e-10, 2.172388e-10, 2.183388e-10, 2.179252e-10, 
    2.186846e-10, 2.188371e-10, 2.176833e-10, 2.183917e-10, 2.161183e-10, 
    2.164856e-10, 2.162669e-10, 2.154682e-10, 2.180204e-10, 2.167106e-10, 
    2.191295e-10, 2.184198e-10, 2.204911e-10, 2.194609e-10, 2.214843e-10, 
    2.223493e-10, 2.231635e-10, 2.241149e-10, 2.160679e-10, 2.157901e-10, 
    2.162875e-10, 2.169756e-10, 2.176142e-10, 2.184631e-10, 2.1855e-10, 
    2.18709e-10, 2.19121e-10, 2.194674e-10, 2.187593e-10, 2.195542e-10, 
    2.165707e-10, 2.181342e-10, 2.156851e-10, 2.164224e-10, 2.16935e-10, 
    2.167102e-10, 2.178779e-10, 2.181531e-10, 2.192715e-10, 2.186934e-10, 
    2.221357e-10, 2.206127e-10, 2.248395e-10, 2.236582e-10, 2.15693e-10, 
    2.160669e-10, 2.173682e-10, 2.16749e-10, 2.185198e-10, 2.189557e-10, 
    2.193101e-10, 2.19763e-10, 2.198119e-10, 2.200803e-10, 2.196405e-10, 
    2.20063e-10, 2.184649e-10, 2.19179e-10, 2.172195e-10, 2.176964e-10, 
    2.17477e-10, 2.172363e-10, 2.179791e-10, 2.187704e-10, 2.187874e-10, 
    2.190411e-10, 2.19756e-10, 2.18527e-10, 2.223322e-10, 2.19982e-10, 
    2.164746e-10, 2.171947e-10, 2.172977e-10, 2.170187e-10, 2.18912e-10, 
    2.182259e-10, 2.200738e-10, 2.195744e-10, 2.203927e-10, 2.199861e-10, 
    2.199262e-10, 2.19404e-10, 2.190788e-10, 2.182574e-10, 2.175891e-10, 
    2.170591e-10, 2.171824e-10, 2.177645e-10, 2.188188e-10, 2.198163e-10, 
    2.195978e-10, 2.203305e-10, 2.183914e-10, 2.192044e-10, 2.188902e-10, 
    2.197096e-10, 2.179142e-10, 2.194429e-10, 2.175234e-10, 2.176917e-10, 
    2.182123e-10, 2.192596e-10, 2.194913e-10, 2.197387e-10, 2.195861e-10, 
    2.188456e-10, 2.187243e-10, 2.181997e-10, 2.180548e-10, 2.176551e-10, 
    2.173241e-10, 2.176265e-10, 2.17944e-10, 2.188459e-10, 2.196587e-10, 
    2.20545e-10, 2.207619e-10, 2.217973e-10, 2.209543e-10, 2.223453e-10, 
    2.211626e-10, 2.2321e-10, 2.195316e-10, 2.211279e-10, 2.18236e-10, 
    2.185476e-10, 2.19111e-10, 2.204035e-10, 2.197058e-10, 2.205218e-10, 
    2.187196e-10, 2.177845e-10, 2.175427e-10, 2.170914e-10, 2.17553e-10, 
    2.175155e-10, 2.179572e-10, 2.178153e-10, 2.188759e-10, 2.183062e-10, 
    2.199247e-10, 2.205154e-10, 2.221836e-10, 2.232064e-10, 2.242476e-10, 
    2.247073e-10, 2.248472e-10, 2.249057e-10 ;

 SOIL2N_TO_SOIL3N =
  1.526171e-11, 1.532907e-11, 1.531597e-11, 1.53703e-11, 1.534016e-11, 
    1.537573e-11, 1.527537e-11, 1.533174e-11, 1.529575e-11, 1.526778e-11, 
    1.547572e-11, 1.537272e-11, 1.558274e-11, 1.551704e-11, 1.568209e-11, 
    1.557252e-11, 1.570419e-11, 1.567894e-11, 1.575496e-11, 1.573318e-11, 
    1.583042e-11, 1.576501e-11, 1.588083e-11, 1.58148e-11, 1.582513e-11, 
    1.576285e-11, 1.539345e-11, 1.54629e-11, 1.538934e-11, 1.539924e-11, 
    1.53948e-11, 1.534078e-11, 1.531356e-11, 1.525657e-11, 1.526692e-11, 
    1.530878e-11, 1.540369e-11, 1.537147e-11, 1.545268e-11, 1.545085e-11, 
    1.554125e-11, 1.550049e-11, 1.565246e-11, 1.560927e-11, 1.573409e-11, 
    1.57027e-11, 1.573261e-11, 1.572354e-11, 1.573273e-11, 1.568669e-11, 
    1.570642e-11, 1.566591e-11, 1.550812e-11, 1.555449e-11, 1.54162e-11, 
    1.533306e-11, 1.527784e-11, 1.523866e-11, 1.52442e-11, 1.525476e-11, 
    1.530902e-11, 1.536005e-11, 1.539894e-11, 1.542495e-11, 1.545058e-11, 
    1.552816e-11, 1.556923e-11, 1.566119e-11, 1.56446e-11, 1.567271e-11, 
    1.569957e-11, 1.574467e-11, 1.573725e-11, 1.575712e-11, 1.567197e-11, 
    1.572856e-11, 1.563515e-11, 1.566069e-11, 1.545754e-11, 1.538017e-11, 
    1.534727e-11, 1.531849e-11, 1.524846e-11, 1.529682e-11, 1.527775e-11, 
    1.532311e-11, 1.535194e-11, 1.533768e-11, 1.542566e-11, 1.539146e-11, 
    1.557167e-11, 1.549404e-11, 1.569644e-11, 1.564801e-11, 1.570805e-11, 
    1.567741e-11, 1.572991e-11, 1.568266e-11, 1.576451e-11, 1.578233e-11, 
    1.577015e-11, 1.581694e-11, 1.568004e-11, 1.573261e-11, 1.533728e-11, 
    1.533961e-11, 1.535044e-11, 1.530282e-11, 1.529991e-11, 1.525628e-11, 
    1.529511e-11, 1.531164e-11, 1.535361e-11, 1.537843e-11, 1.540203e-11, 
    1.545392e-11, 1.551187e-11, 1.559291e-11, 1.565114e-11, 1.569018e-11, 
    1.566624e-11, 1.568737e-11, 1.566375e-11, 1.565268e-11, 1.577565e-11, 
    1.57066e-11, 1.581021e-11, 1.580448e-11, 1.575759e-11, 1.580513e-11, 
    1.534124e-11, 1.532786e-11, 1.528141e-11, 1.531776e-11, 1.525153e-11, 
    1.52886e-11, 1.530992e-11, 1.539217e-11, 1.541024e-11, 1.5427e-11, 
    1.54601e-11, 1.550258e-11, 1.55771e-11, 1.564194e-11, 1.570114e-11, 
    1.56968e-11, 1.569833e-11, 1.571155e-11, 1.567879e-11, 1.571693e-11, 
    1.572333e-11, 1.570659e-11, 1.580371e-11, 1.577597e-11, 1.580436e-11, 
    1.578629e-11, 1.533221e-11, 1.535472e-11, 1.534256e-11, 1.536543e-11, 
    1.534931e-11, 1.542097e-11, 1.544246e-11, 1.5543e-11, 1.550174e-11, 
    1.556741e-11, 1.550841e-11, 1.551887e-11, 1.556955e-11, 1.55116e-11, 
    1.563836e-11, 1.555242e-11, 1.571206e-11, 1.562623e-11, 1.571744e-11, 
    1.570088e-11, 1.57283e-11, 1.575286e-11, 1.578376e-11, 1.584078e-11, 
    1.582758e-11, 1.587526e-11, 1.538828e-11, 1.541748e-11, 1.541491e-11, 
    1.544547e-11, 1.546807e-11, 1.551706e-11, 1.559563e-11, 1.556608e-11, 
    1.562033e-11, 1.563122e-11, 1.554881e-11, 1.55994e-11, 1.543702e-11, 
    1.546325e-11, 1.544764e-11, 1.539058e-11, 1.557289e-11, 1.547932e-11, 
    1.565211e-11, 1.560142e-11, 1.574936e-11, 1.567578e-11, 1.582031e-11, 
    1.588209e-11, 1.594025e-11, 1.600821e-11, 1.543342e-11, 1.541358e-11, 
    1.544911e-11, 1.549826e-11, 1.554387e-11, 1.560451e-11, 1.561071e-11, 
    1.562207e-11, 1.56515e-11, 1.567624e-11, 1.562566e-11, 1.568244e-11, 
    1.546933e-11, 1.558101e-11, 1.540608e-11, 1.545875e-11, 1.549536e-11, 
    1.54793e-11, 1.556271e-11, 1.558237e-11, 1.566225e-11, 1.562096e-11, 
    1.586684e-11, 1.575805e-11, 1.605996e-11, 1.597558e-11, 1.540664e-11, 
    1.543335e-11, 1.55263e-11, 1.548207e-11, 1.560856e-11, 1.563969e-11, 
    1.5665e-11, 1.569736e-11, 1.570085e-11, 1.572002e-11, 1.568861e-11, 
    1.571878e-11, 1.560464e-11, 1.565565e-11, 1.551568e-11, 1.554974e-11, 
    1.553407e-11, 1.551688e-11, 1.556993e-11, 1.562646e-11, 1.562767e-11, 
    1.564579e-11, 1.569686e-11, 1.560907e-11, 1.588087e-11, 1.5713e-11, 
    1.546247e-11, 1.551391e-11, 1.552126e-11, 1.550133e-11, 1.563657e-11, 
    1.558757e-11, 1.571956e-11, 1.568388e-11, 1.574233e-11, 1.571329e-11, 
    1.570902e-11, 1.567171e-11, 1.564849e-11, 1.558981e-11, 1.554208e-11, 
    1.550422e-11, 1.551303e-11, 1.555461e-11, 1.562992e-11, 1.570117e-11, 
    1.568556e-11, 1.573789e-11, 1.559938e-11, 1.565746e-11, 1.563501e-11, 
    1.569355e-11, 1.55653e-11, 1.567449e-11, 1.553739e-11, 1.554941e-11, 
    1.558659e-11, 1.56614e-11, 1.567795e-11, 1.569562e-11, 1.568472e-11, 
    1.563183e-11, 1.562317e-11, 1.558569e-11, 1.557534e-11, 1.554679e-11, 
    1.552315e-11, 1.554475e-11, 1.556743e-11, 1.563185e-11, 1.568991e-11, 
    1.575321e-11, 1.576871e-11, 1.584266e-11, 1.578245e-11, 1.588181e-11, 
    1.579733e-11, 1.594357e-11, 1.568083e-11, 1.579485e-11, 1.558829e-11, 
    1.561054e-11, 1.565079e-11, 1.574311e-11, 1.569327e-11, 1.575156e-11, 
    1.562283e-11, 1.555604e-11, 1.553876e-11, 1.550652e-11, 1.55395e-11, 
    1.553682e-11, 1.556837e-11, 1.555823e-11, 1.563399e-11, 1.55933e-11, 
    1.570891e-11, 1.57511e-11, 1.587026e-11, 1.594331e-11, 1.601769e-11, 
    1.605052e-11, 1.606051e-11, 1.606469e-11 ;

 SOIL2N_vr =
  1.818715, 1.818716, 1.818716, 1.818717, 1.818717, 1.818717, 1.818715, 
    1.818717, 1.818716, 1.818715, 1.81872, 1.818717, 1.818722, 1.818721, 
    1.818724, 1.818722, 1.818725, 1.818724, 1.818726, 1.818725, 1.818727, 
    1.818726, 1.818728, 1.818727, 1.818727, 1.818726, 1.818718, 1.818719, 
    1.818718, 1.818718, 1.818718, 1.818717, 1.818716, 1.818715, 1.818715, 
    1.818716, 1.818718, 1.818717, 1.818719, 1.818719, 1.818721, 1.81872, 
    1.818723, 1.818722, 1.818725, 1.818725, 1.818725, 1.818725, 1.818725, 
    1.818724, 1.818725, 1.818724, 1.81872, 1.818721, 1.818718, 1.818717, 
    1.818715, 1.818714, 1.818715, 1.818715, 1.818716, 1.818717, 1.818718, 
    1.818719, 1.818719, 1.818721, 1.818722, 1.818724, 1.818723, 1.818724, 
    1.818725, 1.818725, 1.818725, 1.818726, 1.818724, 1.818725, 1.818723, 
    1.818724, 1.818719, 1.818718, 1.818717, 1.818716, 1.818715, 1.818716, 
    1.818715, 1.818716, 1.818717, 1.818717, 1.818719, 1.818718, 1.818722, 
    1.81872, 1.818724, 1.818723, 1.818725, 1.818724, 1.818725, 1.818724, 
    1.818726, 1.818726, 1.818726, 1.818727, 1.818724, 1.818725, 1.818717, 
    1.818717, 1.818717, 1.818716, 1.818716, 1.818715, 1.818716, 1.818716, 
    1.818717, 1.818717, 1.818718, 1.818719, 1.81872, 1.818722, 1.818723, 
    1.818724, 1.818724, 1.818724, 1.818724, 1.818723, 1.818726, 1.818725, 
    1.818727, 1.818727, 1.818726, 1.818727, 1.818717, 1.818716, 1.818715, 
    1.818716, 1.818715, 1.818716, 1.818716, 1.818718, 1.818718, 1.818719, 
    1.818719, 1.81872, 1.818722, 1.818723, 1.818725, 1.818724, 1.818725, 
    1.818725, 1.818724, 1.818725, 1.818725, 1.818725, 1.818727, 1.818726, 
    1.818727, 1.818726, 1.818717, 1.818717, 1.818717, 1.818717, 1.818717, 
    1.818718, 1.818719, 1.818721, 1.81872, 1.818722, 1.81872, 1.818721, 
    1.818722, 1.81872, 1.818723, 1.818721, 1.818725, 1.818723, 1.818725, 
    1.818725, 1.818725, 1.818726, 1.818726, 1.818727, 1.818727, 1.818728, 
    1.818718, 1.818718, 1.818718, 1.818719, 1.81872, 1.818721, 1.818722, 
    1.818722, 1.818723, 1.818723, 1.818721, 1.818722, 1.818719, 1.818719, 
    1.818719, 1.818718, 1.818722, 1.81872, 1.818723, 1.818722, 1.818726, 
    1.818724, 1.818727, 1.818728, 1.81873, 1.818731, 1.818719, 1.818718, 
    1.818719, 1.81872, 1.818721, 1.818722, 1.818723, 1.818723, 1.818723, 
    1.818724, 1.818723, 1.818724, 1.81872, 1.818722, 1.818718, 1.818719, 
    1.81872, 1.81872, 1.818722, 1.818722, 1.818724, 1.818723, 1.818728, 
    1.818726, 1.818732, 1.81873, 1.818718, 1.818719, 1.818721, 1.81872, 
    1.818722, 1.818723, 1.818724, 1.818724, 1.818725, 1.818725, 1.818724, 
    1.818725, 1.818722, 1.818724, 1.81872, 1.818721, 1.818721, 1.818721, 
    1.818722, 1.818723, 1.818723, 1.818723, 1.818724, 1.818722, 1.818728, 
    1.818725, 1.818719, 1.81872, 1.818721, 1.81872, 1.818723, 1.818722, 
    1.818725, 1.818724, 1.818725, 1.818725, 1.818725, 1.818724, 1.818723, 
    1.818722, 1.818721, 1.81872, 1.81872, 1.818721, 1.818723, 1.818725, 
    1.818724, 1.818725, 1.818722, 1.818724, 1.818723, 1.818724, 1.818722, 
    1.818724, 1.818721, 1.818721, 1.818722, 1.818724, 1.818724, 1.818724, 
    1.818724, 1.818723, 1.818723, 1.818722, 1.818722, 1.818721, 1.818721, 
    1.818721, 1.818722, 1.818723, 1.818724, 1.818726, 1.818726, 1.818728, 
    1.818726, 1.818728, 1.818727, 1.81873, 1.818724, 1.818727, 1.818722, 
    1.818723, 1.818723, 1.818725, 1.818724, 1.818726, 1.818723, 1.818721, 
    1.818721, 1.81872, 1.818721, 1.818721, 1.818722, 1.818721, 1.818723, 
    1.818722, 1.818725, 1.818726, 1.818728, 1.81873, 1.818731, 1.818732, 
    1.818732, 1.818732,
  1.818667, 1.818669, 1.818668, 1.81867, 1.818669, 1.81867, 1.818667, 
    1.818669, 1.818668, 1.818667, 1.818673, 1.81867, 1.818676, 1.818674, 
    1.818678, 1.818676, 1.818679, 1.818678, 1.818681, 1.81868, 1.818683, 
    1.818681, 1.818684, 1.818682, 1.818682, 1.818681, 1.818671, 1.818673, 
    1.818671, 1.818671, 1.818671, 1.818669, 1.818668, 1.818667, 1.818667, 
    1.818668, 1.818671, 1.81867, 1.818672, 1.818672, 1.818675, 1.818673, 
    1.818678, 1.818676, 1.81868, 1.818679, 1.81868, 1.81868, 1.81868, 
    1.818679, 1.818679, 1.818678, 1.818674, 1.818675, 1.818671, 1.818669, 
    1.818667, 1.818666, 1.818667, 1.818667, 1.818668, 1.81867, 1.818671, 
    1.818671, 1.818672, 1.818674, 1.818675, 1.818678, 1.818677, 1.818678, 
    1.818679, 1.81868, 1.81868, 1.818681, 1.818678, 1.81868, 1.818677, 
    1.818678, 1.818672, 1.81867, 1.818669, 1.818669, 1.818667, 1.818668, 
    1.818667, 1.818669, 1.818669, 1.818669, 1.818671, 1.818671, 1.818676, 
    1.818673, 1.818679, 1.818678, 1.818679, 1.818678, 1.81868, 1.818678, 
    1.818681, 1.818681, 1.818681, 1.818682, 1.818678, 1.81868, 1.818669, 
    1.818669, 1.818669, 1.818668, 1.818668, 1.818667, 1.818668, 1.818668, 
    1.81867, 1.81867, 1.818671, 1.818672, 1.818674, 1.818676, 1.818678, 
    1.818679, 1.818678, 1.818679, 1.818678, 1.818678, 1.818681, 1.818679, 
    1.818682, 1.818682, 1.818681, 1.818682, 1.818669, 1.818669, 1.818668, 
    1.818669, 1.818667, 1.818668, 1.818668, 1.818671, 1.818671, 1.818672, 
    1.818672, 1.818674, 1.818676, 1.818677, 1.818679, 1.818679, 1.818679, 
    1.818679, 1.818678, 1.818679, 1.81868, 1.818679, 1.818682, 1.818681, 
    1.818682, 1.818681, 1.818669, 1.81867, 1.818669, 1.81867, 1.818669, 
    1.818671, 1.818672, 1.818675, 1.818674, 1.818675, 1.818674, 1.818674, 
    1.818675, 1.818674, 1.818677, 1.818675, 1.818679, 1.818677, 1.818679, 
    1.818679, 1.81868, 1.81868, 1.818681, 1.818683, 1.818682, 1.818684, 
    1.818671, 1.818671, 1.818671, 1.818672, 1.818673, 1.818674, 1.818676, 
    1.818675, 1.818677, 1.818677, 1.818675, 1.818676, 1.818672, 1.818673, 
    1.818672, 1.818671, 1.818676, 1.818673, 1.818678, 1.818676, 1.81868, 
    1.818678, 1.818682, 1.818684, 1.818686, 1.818687, 1.818672, 1.818671, 
    1.818672, 1.818673, 1.818675, 1.818676, 1.818677, 1.818677, 1.818678, 
    1.818678, 1.818677, 1.818678, 1.818673, 1.818676, 1.818671, 1.818672, 
    1.818673, 1.818673, 1.818675, 1.818676, 1.818678, 1.818677, 1.818684, 
    1.818681, 1.818689, 1.818686, 1.818671, 1.818672, 1.818674, 1.818673, 
    1.818676, 1.818677, 1.818678, 1.818679, 1.818679, 1.81868, 1.818679, 
    1.818679, 1.818676, 1.818678, 1.818674, 1.818675, 1.818674, 1.818674, 
    1.818675, 1.818677, 1.818677, 1.818678, 1.818679, 1.818676, 1.818684, 
    1.818679, 1.818673, 1.818674, 1.818674, 1.818674, 1.818677, 1.818676, 
    1.818679, 1.818678, 1.81868, 1.818679, 1.818679, 1.818678, 1.818678, 
    1.818676, 1.818675, 1.818674, 1.818674, 1.818675, 1.818677, 1.818679, 
    1.818679, 1.81868, 1.818676, 1.818678, 1.818677, 1.818679, 1.818675, 
    1.818678, 1.818675, 1.818675, 1.818676, 1.818678, 1.818678, 1.818679, 
    1.818679, 1.818677, 1.818677, 1.818676, 1.818676, 1.818675, 1.818674, 
    1.818675, 1.818675, 1.818677, 1.818679, 1.81868, 1.818681, 1.818683, 
    1.818681, 1.818684, 1.818682, 1.818686, 1.818678, 1.818682, 1.818676, 
    1.818677, 1.818678, 1.81868, 1.818679, 1.81868, 1.818677, 1.818675, 
    1.818675, 1.818674, 1.818675, 1.818675, 1.818675, 1.818675, 1.818677, 
    1.818676, 1.818679, 1.81868, 1.818684, 1.818686, 1.818688, 1.818689, 
    1.818689, 1.818689,
  1.818639, 1.818641, 1.818641, 1.818642, 1.818642, 1.818643, 1.81864, 
    1.818641, 1.81864, 1.818639, 1.818646, 1.818642, 1.818649, 1.818647, 
    1.818652, 1.818648, 1.818652, 1.818652, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818656, 1.818656, 1.818654, 1.818643, 1.818645, 
    1.818643, 1.818643, 1.818643, 1.818642, 1.818641, 1.818639, 1.818639, 
    1.818641, 1.818643, 1.818642, 1.818645, 1.818645, 1.818648, 1.818646, 
    1.818651, 1.81865, 1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 
    1.818652, 1.818653, 1.818651, 1.818647, 1.818648, 1.818644, 1.818641, 
    1.81864, 1.818638, 1.818639, 1.818639, 1.818641, 1.818642, 1.818643, 
    1.818644, 1.818645, 1.818647, 1.818648, 1.818651, 1.818651, 1.818652, 
    1.818652, 1.818654, 1.818653, 1.818654, 1.818651, 1.818653, 1.81865, 
    1.818651, 1.818645, 1.818643, 1.818642, 1.818641, 1.818639, 1.81864, 
    1.81864, 1.818641, 1.818642, 1.818641, 1.818644, 1.818643, 1.818648, 
    1.818646, 1.818652, 1.818651, 1.818653, 1.818652, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818654, 1.818656, 1.818652, 1.818653, 1.818641, 
    1.818642, 1.818642, 1.81864, 1.81864, 1.818639, 1.81864, 1.818641, 
    1.818642, 1.818643, 1.818643, 1.818645, 1.818647, 1.818649, 1.818651, 
    1.818652, 1.818651, 1.818652, 1.818651, 1.818651, 1.818655, 1.818653, 
    1.818656, 1.818655, 1.818654, 1.818655, 1.818642, 1.818641, 1.81864, 
    1.818641, 1.818639, 1.81864, 1.818641, 1.818643, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818649, 1.818651, 1.818652, 1.818652, 1.818652, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 1.818655, 1.818655, 
    1.818655, 1.818655, 1.818641, 1.818642, 1.818642, 1.818642, 1.818642, 
    1.818644, 1.818645, 1.818648, 1.818646, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.818647, 1.81865, 1.818648, 1.818653, 1.81865, 1.818653, 
    1.818652, 1.818653, 1.818654, 1.818655, 1.818657, 1.818656, 1.818658, 
    1.818643, 1.818644, 1.818644, 1.818645, 1.818645, 1.818647, 1.818649, 
    1.818648, 1.81865, 1.81865, 1.818648, 1.818649, 1.818644, 1.818645, 
    1.818645, 1.818643, 1.818648, 1.818646, 1.818651, 1.818649, 1.818654, 
    1.818652, 1.818656, 1.818658, 1.81866, 1.818662, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818648, 1.818649, 1.81865, 1.81865, 1.818651, 
    1.818652, 1.81865, 1.818652, 1.818645, 1.818649, 1.818643, 1.818645, 
    1.818646, 1.818646, 1.818648, 1.818649, 1.818651, 1.81865, 1.818657, 
    1.818654, 1.818663, 1.818661, 1.818644, 1.818644, 1.818647, 1.818646, 
    1.81865, 1.81865, 1.818651, 1.818652, 1.818652, 1.818653, 1.818652, 
    1.818653, 1.818649, 1.818651, 1.818647, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.81865, 1.81865, 1.818651, 1.818652, 1.81865, 1.818658, 
    1.818653, 1.818645, 1.818647, 1.818647, 1.818646, 1.81865, 1.818649, 
    1.818653, 1.818652, 1.818654, 1.818653, 1.818653, 1.818651, 1.818651, 
    1.818649, 1.818648, 1.818646, 1.818647, 1.818648, 1.81865, 1.818652, 
    1.818652, 1.818653, 1.818649, 1.818651, 1.81865, 1.818652, 1.818648, 
    1.818652, 1.818647, 1.818648, 1.818649, 1.818651, 1.818652, 1.818652, 
    1.818652, 1.81865, 1.81865, 1.818649, 1.818649, 1.818648, 1.818647, 
    1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818654, 1.818657, 
    1.818655, 1.818658, 1.818655, 1.81866, 1.818652, 1.818655, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818652, 1.818654, 1.81865, 1.818648, 
    1.818648, 1.818647, 1.818648, 1.818647, 1.818648, 1.818648, 1.81865, 
    1.818649, 1.818653, 1.818654, 1.818657, 1.81866, 1.818662, 1.818663, 
    1.818663, 1.818663,
  1.818617, 1.818619, 1.818619, 1.818621, 1.81862, 1.818621, 1.818618, 
    1.818619, 1.818618, 1.818618, 1.818624, 1.818621, 1.818627, 1.818625, 
    1.81863, 1.818627, 1.818631, 1.81863, 1.818632, 1.818632, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818635, 1.818633, 1.818621, 1.818624, 
    1.818621, 1.818622, 1.818622, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818619, 1.818622, 1.818621, 1.818623, 1.818623, 1.818626, 1.818625, 
    1.818629, 1.818628, 1.818632, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.81863, 1.818631, 1.81863, 1.818625, 1.818626, 1.818622, 1.81862, 
    1.818618, 1.818617, 1.818617, 1.818617, 1.818619, 1.81862, 1.818622, 
    1.818622, 1.818623, 1.818626, 1.818627, 1.81863, 1.818629, 1.81863, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.81863, 1.818632, 1.818629, 
    1.81863, 1.818623, 1.818621, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818618, 1.818619, 1.81862, 1.81862, 1.818622, 1.818621, 1.818627, 
    1.818624, 1.818631, 1.818629, 1.818631, 1.81863, 1.818632, 1.81863, 
    1.818633, 1.818633, 1.818633, 1.818634, 1.81863, 1.818632, 1.81862, 
    1.81862, 1.81862, 1.818619, 1.818619, 1.818617, 1.818618, 1.818619, 
    1.81862, 1.818621, 1.818622, 1.818623, 1.818625, 1.818628, 1.818629, 
    1.818631, 1.81863, 1.81863, 1.81863, 1.818629, 1.818633, 1.818631, 
    1.818634, 1.818634, 1.818633, 1.818634, 1.81862, 1.818619, 1.818618, 
    1.818619, 1.818617, 1.818618, 1.818619, 1.818621, 1.818622, 1.818622, 
    1.818623, 1.818625, 1.818627, 1.818629, 1.818631, 1.818631, 1.818631, 
    1.818631, 1.81863, 1.818631, 1.818632, 1.818631, 1.818634, 1.818633, 
    1.818634, 1.818633, 1.81862, 1.81862, 1.81862, 1.818621, 1.81862, 
    1.818622, 1.818623, 1.818626, 1.818625, 1.818627, 1.818625, 1.818625, 
    1.818627, 1.818625, 1.818629, 1.818626, 1.818631, 1.818629, 1.818631, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.818635, 1.818635, 1.818636, 
    1.818621, 1.818622, 1.818622, 1.818623, 1.818624, 1.818625, 1.818628, 
    1.818627, 1.818628, 1.818629, 1.818626, 1.818628, 1.818623, 1.818624, 
    1.818623, 1.818621, 1.818627, 1.818624, 1.818629, 1.818628, 1.818632, 
    1.81863, 1.818635, 1.818636, 1.818638, 1.81864, 1.818623, 1.818622, 
    1.818623, 1.818625, 1.818626, 1.818628, 1.818628, 1.818628, 1.818629, 
    1.81863, 1.818629, 1.81863, 1.818624, 1.818627, 1.818622, 1.818623, 
    1.818625, 1.818624, 1.818627, 1.818627, 1.81863, 1.818628, 1.818636, 
    1.818633, 1.818642, 1.818639, 1.818622, 1.818623, 1.818625, 1.818624, 
    1.818628, 1.818629, 1.81863, 1.818631, 1.818631, 1.818631, 1.81863, 
    1.818631, 1.818628, 1.81863, 1.818625, 1.818626, 1.818626, 1.818625, 
    1.818627, 1.818629, 1.818629, 1.818629, 1.818631, 1.818628, 1.818636, 
    1.818631, 1.818624, 1.818625, 1.818625, 1.818625, 1.818629, 1.818627, 
    1.818631, 1.81863, 1.818632, 1.818631, 1.818631, 1.81863, 1.818629, 
    1.818627, 1.818626, 1.818625, 1.818625, 1.818626, 1.818629, 1.818631, 
    1.81863, 1.818632, 1.818628, 1.81863, 1.818629, 1.818631, 1.818627, 
    1.81863, 1.818626, 1.818626, 1.818627, 1.81863, 1.81863, 1.818631, 
    1.81863, 1.818629, 1.818628, 1.818627, 1.818627, 1.818626, 1.818625, 
    1.818626, 1.818627, 1.818629, 1.818631, 1.818632, 1.818633, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818638, 1.81863, 1.818634, 1.818627, 
    1.818628, 1.818629, 1.818632, 1.818631, 1.818632, 1.818628, 1.818626, 
    1.818626, 1.818625, 1.818626, 1.818626, 1.818627, 1.818627, 1.818629, 
    1.818628, 1.818631, 1.818632, 1.818636, 1.818638, 1.818641, 1.818642, 
    1.818642, 1.818642,
  1.818569, 1.81857, 1.81857, 1.818572, 1.818571, 1.818572, 1.818569, 
    1.81857, 1.81857, 1.818569, 1.818574, 1.818572, 1.818577, 1.818576, 
    1.81858, 1.818577, 1.818581, 1.81858, 1.818582, 1.818581, 1.818584, 
    1.818582, 1.818585, 1.818583, 1.818584, 1.818582, 1.818572, 1.818574, 
    1.818572, 1.818572, 1.818572, 1.818571, 1.81857, 1.818568, 1.818569, 
    1.81857, 1.818572, 1.818572, 1.818574, 1.818574, 1.818576, 1.818575, 
    1.818579, 1.818578, 1.818581, 1.818581, 1.818581, 1.818581, 1.818581, 
    1.81858, 1.818581, 1.818579, 1.818575, 1.818576, 1.818573, 1.818571, 
    1.818569, 1.818568, 1.818568, 1.818568, 1.81857, 1.818571, 1.818572, 
    1.818573, 1.818574, 1.818576, 1.818577, 1.818579, 1.818579, 1.81858, 
    1.81858, 1.818582, 1.818581, 1.818582, 1.81858, 1.818581, 1.818579, 
    1.818579, 1.818574, 1.818572, 1.818571, 1.81857, 1.818568, 1.81857, 
    1.818569, 1.81857, 1.818571, 1.818571, 1.818573, 1.818572, 1.818577, 
    1.818575, 1.81858, 1.818579, 1.818581, 1.81858, 1.818581, 1.81858, 
    1.818582, 1.818583, 1.818582, 1.818583, 1.81858, 1.818581, 1.818571, 
    1.818571, 1.818571, 1.81857, 1.81857, 1.818568, 1.81857, 1.81857, 
    1.818571, 1.818572, 1.818572, 1.818574, 1.818575, 1.818578, 1.818579, 
    1.81858, 1.818579, 1.81858, 1.818579, 1.818579, 1.818582, 1.818581, 
    1.818583, 1.818583, 1.818582, 1.818583, 1.818571, 1.81857, 1.818569, 
    1.81857, 1.818568, 1.818569, 1.81857, 1.818572, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818577, 1.818579, 1.81858, 1.81858, 1.81858, 
    1.818581, 1.81858, 1.818581, 1.818581, 1.818581, 1.818583, 1.818582, 
    1.818583, 1.818583, 1.81857, 1.818571, 1.818571, 1.818571, 1.818571, 
    1.818573, 1.818573, 1.818576, 1.818575, 1.818577, 1.818575, 1.818576, 
    1.818577, 1.818575, 1.818579, 1.818576, 1.818581, 1.818578, 1.818581, 
    1.81858, 1.818581, 1.818582, 1.818583, 1.818584, 1.818584, 1.818585, 
    1.818572, 1.818573, 1.818573, 1.818574, 1.818574, 1.818576, 1.818578, 
    1.818577, 1.818578, 1.818579, 1.818576, 1.818578, 1.818573, 1.818574, 
    1.818574, 1.818572, 1.818577, 1.818574, 1.818579, 1.818578, 1.818582, 
    1.81858, 1.818584, 1.818585, 1.818587, 1.818589, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818576, 1.818578, 1.818578, 1.818578, 1.818579, 
    1.81858, 1.818578, 1.81858, 1.818574, 1.818577, 1.818573, 1.818574, 
    1.818575, 1.818574, 1.818577, 1.818577, 1.818579, 1.818578, 1.818585, 
    1.818582, 1.81859, 1.818588, 1.818573, 1.818573, 1.818576, 1.818575, 
    1.818578, 1.818579, 1.818579, 1.81858, 1.81858, 1.818581, 1.81858, 
    1.818581, 1.818578, 1.818579, 1.818576, 1.818576, 1.818576, 1.818576, 
    1.818577, 1.818578, 1.818578, 1.818579, 1.81858, 1.818578, 1.818585, 
    1.818581, 1.818574, 1.818575, 1.818576, 1.818575, 1.818579, 1.818577, 
    1.818581, 1.81858, 1.818582, 1.818581, 1.818581, 1.81858, 1.818579, 
    1.818577, 1.818576, 1.818575, 1.818575, 1.818576, 1.818578, 1.81858, 
    1.81858, 1.818581, 1.818578, 1.818579, 1.818579, 1.81858, 1.818577, 
    1.81858, 1.818576, 1.818576, 1.818577, 1.818579, 1.81858, 1.81858, 
    1.81858, 1.818579, 1.818578, 1.818577, 1.818577, 1.818576, 1.818576, 
    1.818576, 1.818577, 1.818579, 1.81858, 1.818582, 1.818582, 1.818584, 
    1.818583, 1.818585, 1.818583, 1.818587, 1.81858, 1.818583, 1.818577, 
    1.818578, 1.818579, 1.818582, 1.81858, 1.818582, 1.818578, 1.818577, 
    1.818576, 1.818575, 1.818576, 1.818576, 1.818577, 1.818577, 1.818579, 
    1.818578, 1.818581, 1.818582, 1.818585, 1.818587, 1.818589, 1.81859, 
    1.81859, 1.81859,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.292667e-09, 1.298372e-09, 1.297263e-09, 1.301864e-09, 1.299312e-09, 
    1.302325e-09, 1.293824e-09, 1.298598e-09, 1.29555e-09, 1.293181e-09, 
    1.310794e-09, 1.302069e-09, 1.319858e-09, 1.314293e-09, 1.328273e-09, 
    1.318992e-09, 1.330145e-09, 1.328006e-09, 1.334445e-09, 1.3326e-09, 
    1.340836e-09, 1.335297e-09, 1.345106e-09, 1.339513e-09, 1.340388e-09, 
    1.335114e-09, 1.303825e-09, 1.309707e-09, 1.303477e-09, 1.304316e-09, 
    1.303939e-09, 1.299364e-09, 1.297059e-09, 1.292231e-09, 1.293108e-09, 
    1.296654e-09, 1.304693e-09, 1.301964e-09, 1.308842e-09, 1.308687e-09, 
    1.316344e-09, 1.312892e-09, 1.325763e-09, 1.322105e-09, 1.332677e-09, 
    1.330018e-09, 1.332553e-09, 1.331784e-09, 1.332563e-09, 1.328663e-09, 
    1.330334e-09, 1.326902e-09, 1.313538e-09, 1.317465e-09, 1.305753e-09, 
    1.29871e-09, 1.294033e-09, 1.290714e-09, 1.291184e-09, 1.292078e-09, 
    1.296674e-09, 1.300996e-09, 1.30429e-09, 1.306493e-09, 1.308664e-09, 
    1.315235e-09, 1.318714e-09, 1.326503e-09, 1.325098e-09, 1.327479e-09, 
    1.329754e-09, 1.333573e-09, 1.332945e-09, 1.334628e-09, 1.327416e-09, 
    1.332209e-09, 1.324297e-09, 1.326461e-09, 1.309253e-09, 1.3027e-09, 
    1.299914e-09, 1.297476e-09, 1.291544e-09, 1.29564e-09, 1.294026e-09, 
    1.297868e-09, 1.300309e-09, 1.299102e-09, 1.306554e-09, 1.303656e-09, 
    1.31892e-09, 1.312345e-09, 1.329489e-09, 1.325386e-09, 1.330472e-09, 
    1.327877e-09, 1.332323e-09, 1.328321e-09, 1.335254e-09, 1.336764e-09, 
    1.335732e-09, 1.339695e-09, 1.3281e-09, 1.332552e-09, 1.299068e-09, 
    1.299265e-09, 1.300182e-09, 1.296149e-09, 1.295902e-09, 1.292207e-09, 
    1.295495e-09, 1.296896e-09, 1.300451e-09, 1.302553e-09, 1.304552e-09, 
    1.308947e-09, 1.313855e-09, 1.32072e-09, 1.325652e-09, 1.328958e-09, 
    1.326931e-09, 1.328721e-09, 1.32672e-09, 1.325782e-09, 1.336198e-09, 
    1.330349e-09, 1.339125e-09, 1.338639e-09, 1.334668e-09, 1.338694e-09, 
    1.299403e-09, 1.29827e-09, 1.294335e-09, 1.297414e-09, 1.291805e-09, 
    1.294945e-09, 1.29675e-09, 1.303717e-09, 1.305248e-09, 1.306667e-09, 
    1.30947e-09, 1.313068e-09, 1.31938e-09, 1.324872e-09, 1.329886e-09, 
    1.329519e-09, 1.329648e-09, 1.330768e-09, 1.327994e-09, 1.331224e-09, 
    1.331766e-09, 1.330348e-09, 1.338574e-09, 1.336224e-09, 1.338629e-09, 
    1.337099e-09, 1.298638e-09, 1.300545e-09, 1.299514e-09, 1.301452e-09, 
    1.300087e-09, 1.306156e-09, 1.307976e-09, 1.316492e-09, 1.312997e-09, 
    1.31856e-09, 1.313562e-09, 1.314448e-09, 1.318741e-09, 1.313833e-09, 
    1.324569e-09, 1.31729e-09, 1.330812e-09, 1.323542e-09, 1.331267e-09, 
    1.329865e-09, 1.332187e-09, 1.334267e-09, 1.336885e-09, 1.341714e-09, 
    1.340596e-09, 1.344634e-09, 1.303388e-09, 1.305861e-09, 1.305643e-09, 
    1.308231e-09, 1.310146e-09, 1.314295e-09, 1.32095e-09, 1.318447e-09, 
    1.323042e-09, 1.323964e-09, 1.316984e-09, 1.32127e-09, 1.307516e-09, 
    1.309738e-09, 1.308415e-09, 1.303582e-09, 1.319024e-09, 1.311099e-09, 
    1.325733e-09, 1.32144e-09, 1.333971e-09, 1.327739e-09, 1.33998e-09, 
    1.345213e-09, 1.350139e-09, 1.355895e-09, 1.307211e-09, 1.30553e-09, 
    1.308539e-09, 1.312702e-09, 1.316566e-09, 1.321702e-09, 1.322227e-09, 
    1.32319e-09, 1.325682e-09, 1.327778e-09, 1.323494e-09, 1.328303e-09, 
    1.310253e-09, 1.319712e-09, 1.304895e-09, 1.309356e-09, 1.312457e-09, 
    1.311097e-09, 1.318161e-09, 1.319826e-09, 1.326593e-09, 1.323095e-09, 
    1.343921e-09, 1.334707e-09, 1.360279e-09, 1.353132e-09, 1.304943e-09, 
    1.307205e-09, 1.315077e-09, 1.311332e-09, 1.322045e-09, 1.324682e-09, 
    1.326826e-09, 1.329566e-09, 1.329862e-09, 1.331486e-09, 1.328825e-09, 
    1.331381e-09, 1.321713e-09, 1.326033e-09, 1.314178e-09, 1.317063e-09, 
    1.315736e-09, 1.31428e-09, 1.318774e-09, 1.323561e-09, 1.323664e-09, 
    1.325199e-09, 1.329524e-09, 1.322088e-09, 1.34511e-09, 1.330891e-09, 
    1.309671e-09, 1.314028e-09, 1.314651e-09, 1.312963e-09, 1.324417e-09, 
    1.320267e-09, 1.331447e-09, 1.328425e-09, 1.333376e-09, 1.330916e-09, 
    1.330554e-09, 1.327394e-09, 1.325427e-09, 1.320457e-09, 1.316414e-09, 
    1.313208e-09, 1.313953e-09, 1.317475e-09, 1.323854e-09, 1.329889e-09, 
    1.328567e-09, 1.332999e-09, 1.321268e-09, 1.326187e-09, 1.324286e-09, 
    1.329243e-09, 1.318381e-09, 1.32763e-09, 1.316017e-09, 1.317035e-09, 
    1.320185e-09, 1.32652e-09, 1.327923e-09, 1.329419e-09, 1.328496e-09, 
    1.324016e-09, 1.323282e-09, 1.320108e-09, 1.319232e-09, 1.316813e-09, 
    1.314811e-09, 1.31664e-09, 1.318561e-09, 1.324018e-09, 1.328935e-09, 
    1.334297e-09, 1.335609e-09, 1.341874e-09, 1.336774e-09, 1.345189e-09, 
    1.338034e-09, 1.350421e-09, 1.328166e-09, 1.337824e-09, 1.320328e-09, 
    1.322213e-09, 1.325622e-09, 1.333441e-09, 1.32922e-09, 1.334157e-09, 
    1.323253e-09, 1.317596e-09, 1.316133e-09, 1.313403e-09, 1.316196e-09, 
    1.315969e-09, 1.318641e-09, 1.317782e-09, 1.324199e-09, 1.320752e-09, 
    1.330544e-09, 1.334118e-09, 1.344211e-09, 1.350398e-09, 1.356698e-09, 
    1.359479e-09, 1.360325e-09, 1.360679e-09 ;

 SOIL2_HR_S3 =
  9.233337e-11, 9.274085e-11, 9.266164e-11, 9.29903e-11, 9.280799e-11, 
    9.302319e-11, 9.241599e-11, 9.275702e-11, 9.253932e-11, 9.237006e-11, 
    9.362812e-11, 9.300496e-11, 9.427558e-11, 9.387809e-11, 9.487668e-11, 
    9.421371e-11, 9.501037e-11, 9.485757e-11, 9.531751e-11, 9.518575e-11, 
    9.577401e-11, 9.537833e-11, 9.607901e-11, 9.567953e-11, 9.574201e-11, 
    9.536527e-11, 9.313039e-11, 9.355053e-11, 9.310549e-11, 9.31654e-11, 
    9.313852e-11, 9.281174e-11, 9.264706e-11, 9.230224e-11, 9.236484e-11, 
    9.261811e-11, 9.319234e-11, 9.299743e-11, 9.348872e-11, 9.347762e-11, 
    9.402459e-11, 9.377796e-11, 9.469738e-11, 9.443606e-11, 9.519124e-11, 
    9.500131e-11, 9.518232e-11, 9.512744e-11, 9.518304e-11, 9.490449e-11, 
    9.502382e-11, 9.477873e-11, 9.382415e-11, 9.410467e-11, 9.326804e-11, 
    9.2765e-11, 9.243094e-11, 9.219388e-11, 9.22274e-11, 9.229128e-11, 
    9.26196e-11, 9.292831e-11, 9.316358e-11, 9.332096e-11, 9.347603e-11, 
    9.394537e-11, 9.419385e-11, 9.475021e-11, 9.464982e-11, 9.48199e-11, 
    9.498242e-11, 9.525525e-11, 9.521035e-11, 9.533055e-11, 9.481543e-11, 
    9.515777e-11, 9.459264e-11, 9.47472e-11, 9.351811e-11, 9.305001e-11, 
    9.2851e-11, 9.267686e-11, 9.225316e-11, 9.254575e-11, 9.243041e-11, 
    9.270484e-11, 9.287921e-11, 9.279297e-11, 9.332526e-11, 9.311831e-11, 
    9.420858e-11, 9.373895e-11, 9.496346e-11, 9.467043e-11, 9.50337e-11, 
    9.484834e-11, 9.516595e-11, 9.48801e-11, 9.537529e-11, 9.548311e-11, 
    9.540943e-11, 9.56925e-11, 9.486426e-11, 9.518231e-11, 9.279055e-11, 
    9.280462e-11, 9.287015e-11, 9.258209e-11, 9.256447e-11, 9.230052e-11, 
    9.253539e-11, 9.26354e-11, 9.288932e-11, 9.303951e-11, 9.318228e-11, 
    9.349621e-11, 9.384682e-11, 9.433713e-11, 9.468942e-11, 9.492557e-11, 
    9.478077e-11, 9.490862e-11, 9.47657e-11, 9.469872e-11, 9.54427e-11, 
    9.502493e-11, 9.565179e-11, 9.56171e-11, 9.533341e-11, 9.562101e-11, 
    9.281449e-11, 9.273356e-11, 9.245253e-11, 9.267245e-11, 9.227178e-11, 
    9.249605e-11, 9.2625e-11, 9.312262e-11, 9.323198e-11, 9.333335e-11, 
    9.35336e-11, 9.379059e-11, 9.424143e-11, 9.463372e-11, 9.499188e-11, 
    9.496564e-11, 9.497488e-11, 9.505488e-11, 9.48567e-11, 9.508742e-11, 
    9.512613e-11, 9.502489e-11, 9.561246e-11, 9.544459e-11, 9.561637e-11, 
    9.550707e-11, 9.275987e-11, 9.289606e-11, 9.282246e-11, 9.296085e-11, 
    9.286335e-11, 9.329688e-11, 9.342687e-11, 9.403515e-11, 9.378553e-11, 
    9.418284e-11, 9.382589e-11, 9.388913e-11, 9.419577e-11, 9.384518e-11, 
    9.461208e-11, 9.409212e-11, 9.505798e-11, 9.453868e-11, 9.509053e-11, 
    9.499033e-11, 9.515624e-11, 9.530482e-11, 9.549177e-11, 9.58367e-11, 
    9.575683e-11, 9.604531e-11, 9.30991e-11, 9.327576e-11, 9.326021e-11, 
    9.344509e-11, 9.358182e-11, 9.38782e-11, 9.435356e-11, 9.417481e-11, 
    9.4503e-11, 9.456887e-11, 9.407029e-11, 9.43764e-11, 9.339399e-11, 
    9.355269e-11, 9.345821e-11, 9.311303e-11, 9.421598e-11, 9.364991e-11, 
    9.469524e-11, 9.438857e-11, 9.528364e-11, 9.483847e-11, 9.571285e-11, 
    9.608664e-11, 9.643852e-11, 9.684967e-11, 9.337218e-11, 9.325215e-11, 
    9.346709e-11, 9.376445e-11, 9.40404e-11, 9.440727e-11, 9.444481e-11, 
    9.451354e-11, 9.469158e-11, 9.484127e-11, 9.453525e-11, 9.48788e-11, 
    9.358947e-11, 9.426512e-11, 9.320675e-11, 9.352542e-11, 9.374693e-11, 
    9.364977e-11, 9.415438e-11, 9.427331e-11, 9.475663e-11, 9.450678e-11, 
    9.599437e-11, 9.533619e-11, 9.716278e-11, 9.665228e-11, 9.32102e-11, 
    9.337178e-11, 9.39341e-11, 9.366654e-11, 9.443177e-11, 9.462013e-11, 
    9.477327e-11, 9.496902e-11, 9.499016e-11, 9.510615e-11, 9.491609e-11, 
    9.509864e-11, 9.440805e-11, 9.471665e-11, 9.386984e-11, 9.407593e-11, 
    9.398112e-11, 9.387712e-11, 9.419811e-11, 9.454007e-11, 9.45474e-11, 
    9.465705e-11, 9.496601e-11, 9.443487e-11, 9.607928e-11, 9.506366e-11, 
    9.354796e-11, 9.385915e-11, 9.390363e-11, 9.378307e-11, 9.460124e-11, 
    9.430478e-11, 9.510332e-11, 9.48875e-11, 9.524113e-11, 9.50654e-11, 
    9.503955e-11, 9.481386e-11, 9.467335e-11, 9.431837e-11, 9.402956e-11, 
    9.380056e-11, 9.385381e-11, 9.410536e-11, 9.456099e-11, 9.499206e-11, 
    9.489763e-11, 9.521425e-11, 9.437628e-11, 9.472764e-11, 9.459183e-11, 
    9.494595e-11, 9.417005e-11, 9.48307e-11, 9.400119e-11, 9.407392e-11, 
    9.42989e-11, 9.475145e-11, 9.485161e-11, 9.495851e-11, 9.489255e-11, 
    9.457257e-11, 9.452015e-11, 9.429343e-11, 9.423082e-11, 9.405809e-11, 
    9.391506e-11, 9.404573e-11, 9.418295e-11, 9.45727e-11, 9.492396e-11, 
    9.530693e-11, 9.540067e-11, 9.584811e-11, 9.548384e-11, 9.608494e-11, 
    9.557385e-11, 9.645862e-11, 9.486902e-11, 9.555885e-11, 9.430914e-11, 
    9.444377e-11, 9.468726e-11, 9.52458e-11, 9.494429e-11, 9.529692e-11, 
    9.45181e-11, 9.411403e-11, 9.400952e-11, 9.381448e-11, 9.401398e-11, 
    9.399775e-11, 9.418865e-11, 9.41273e-11, 9.458565e-11, 9.433945e-11, 
    9.503889e-11, 9.529414e-11, 9.601507e-11, 9.645704e-11, 9.6907e-11, 
    9.710564e-11, 9.71661e-11, 9.719138e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.549107e-11, 2.560354e-11, 2.558168e-11, 2.567239e-11, 2.562208e-11, 
    2.568147e-11, 2.551388e-11, 2.560801e-11, 2.554792e-11, 2.55012e-11, 
    2.584844e-11, 2.567644e-11, 2.602715e-11, 2.591744e-11, 2.619307e-11, 
    2.601008e-11, 2.622997e-11, 2.618779e-11, 2.631474e-11, 2.627837e-11, 
    2.644074e-11, 2.633153e-11, 2.652493e-11, 2.641467e-11, 2.643191e-11, 
    2.632792e-11, 2.571106e-11, 2.582703e-11, 2.570419e-11, 2.572073e-11, 
    2.571331e-11, 2.562311e-11, 2.557766e-11, 2.548248e-11, 2.549976e-11, 
    2.556967e-11, 2.572816e-11, 2.567436e-11, 2.580997e-11, 2.580691e-11, 
    2.595788e-11, 2.588981e-11, 2.614358e-11, 2.607145e-11, 2.627989e-11, 
    2.622747e-11, 2.627743e-11, 2.626228e-11, 2.627763e-11, 2.620074e-11, 
    2.623368e-11, 2.616603e-11, 2.590255e-11, 2.597998e-11, 2.574906e-11, 
    2.561021e-11, 2.5518e-11, 2.545257e-11, 2.546182e-11, 2.547946e-11, 
    2.557008e-11, 2.565529e-11, 2.572022e-11, 2.576366e-11, 2.580646e-11, 
    2.593601e-11, 2.60046e-11, 2.615816e-11, 2.613045e-11, 2.61774e-11, 
    2.622225e-11, 2.629756e-11, 2.628517e-11, 2.631834e-11, 2.617616e-11, 
    2.627065e-11, 2.611467e-11, 2.615733e-11, 2.581808e-11, 2.568888e-11, 
    2.563395e-11, 2.558588e-11, 2.546893e-11, 2.554969e-11, 2.551786e-11, 
    2.55936e-11, 2.564173e-11, 2.561793e-11, 2.576485e-11, 2.570773e-11, 
    2.600866e-11, 2.587904e-11, 2.621702e-11, 2.613614e-11, 2.623641e-11, 
    2.618524e-11, 2.627291e-11, 2.619401e-11, 2.633069e-11, 2.636045e-11, 
    2.634011e-11, 2.641825e-11, 2.618964e-11, 2.627743e-11, 2.561726e-11, 
    2.562114e-11, 2.563923e-11, 2.555972e-11, 2.555486e-11, 2.548201e-11, 
    2.554683e-11, 2.557444e-11, 2.564452e-11, 2.568598e-11, 2.572539e-11, 
    2.581204e-11, 2.590881e-11, 2.604414e-11, 2.614138e-11, 2.620656e-11, 
    2.61666e-11, 2.620188e-11, 2.616244e-11, 2.614395e-11, 2.63493e-11, 
    2.623399e-11, 2.640701e-11, 2.639743e-11, 2.631913e-11, 2.639851e-11, 
    2.562387e-11, 2.560153e-11, 2.552396e-11, 2.558467e-11, 2.547407e-11, 
    2.553597e-11, 2.557157e-11, 2.570892e-11, 2.57391e-11, 2.576708e-11, 
    2.582236e-11, 2.589329e-11, 2.601773e-11, 2.612601e-11, 2.622486e-11, 
    2.621762e-11, 2.622017e-11, 2.624225e-11, 2.618755e-11, 2.625123e-11, 
    2.626192e-11, 2.623398e-11, 2.639615e-11, 2.634982e-11, 2.639723e-11, 
    2.636706e-11, 2.560879e-11, 2.564638e-11, 2.562607e-11, 2.566427e-11, 
    2.563736e-11, 2.575702e-11, 2.57929e-11, 2.596079e-11, 2.589189e-11, 
    2.600156e-11, 2.590303e-11, 2.592049e-11, 2.600513e-11, 2.590836e-11, 
    2.612003e-11, 2.597651e-11, 2.624311e-11, 2.609978e-11, 2.625209e-11, 
    2.622444e-11, 2.627023e-11, 2.631124e-11, 2.636284e-11, 2.645805e-11, 
    2.6436e-11, 2.651562e-11, 2.570243e-11, 2.575119e-11, 2.57469e-11, 
    2.579793e-11, 2.583567e-11, 2.591747e-11, 2.604868e-11, 2.599934e-11, 
    2.608992e-11, 2.610811e-11, 2.597049e-11, 2.605498e-11, 2.578382e-11, 
    2.582762e-11, 2.580155e-11, 2.570627e-11, 2.60107e-11, 2.585446e-11, 
    2.614299e-11, 2.605834e-11, 2.630539e-11, 2.618252e-11, 2.642386e-11, 
    2.652703e-11, 2.662416e-11, 2.673764e-11, 2.57778e-11, 2.574467e-11, 
    2.5804e-11, 2.588607e-11, 2.596224e-11, 2.60635e-11, 2.607387e-11, 
    2.609283e-11, 2.614198e-11, 2.618329e-11, 2.609883e-11, 2.619365e-11, 
    2.583778e-11, 2.602427e-11, 2.573214e-11, 2.58201e-11, 2.588124e-11, 
    2.585442e-11, 2.59937e-11, 2.602653e-11, 2.615993e-11, 2.609097e-11, 
    2.650157e-11, 2.63199e-11, 2.682406e-11, 2.668316e-11, 2.573309e-11, 
    2.577769e-11, 2.59329e-11, 2.585905e-11, 2.607026e-11, 2.612226e-11, 
    2.616453e-11, 2.621855e-11, 2.622439e-11, 2.62564e-11, 2.620394e-11, 
    2.625433e-11, 2.606372e-11, 2.61489e-11, 2.591516e-11, 2.597205e-11, 
    2.594588e-11, 2.591717e-11, 2.600577e-11, 2.610016e-11, 2.610218e-11, 
    2.613245e-11, 2.621772e-11, 2.607112e-11, 2.6525e-11, 2.624467e-11, 
    2.582632e-11, 2.591221e-11, 2.592449e-11, 2.589121e-11, 2.611704e-11, 
    2.603521e-11, 2.625562e-11, 2.619605e-11, 2.629366e-11, 2.624516e-11, 
    2.623802e-11, 2.617573e-11, 2.613695e-11, 2.603896e-11, 2.595925e-11, 
    2.589604e-11, 2.591074e-11, 2.598017e-11, 2.610593e-11, 2.622492e-11, 
    2.619885e-11, 2.628624e-11, 2.605495e-11, 2.615193e-11, 2.611444e-11, 
    2.621219e-11, 2.599803e-11, 2.618038e-11, 2.595142e-11, 2.597149e-11, 
    2.603359e-11, 2.61585e-11, 2.618615e-11, 2.621565e-11, 2.619745e-11, 
    2.610913e-11, 2.609466e-11, 2.603208e-11, 2.60148e-11, 2.596712e-11, 
    2.592765e-11, 2.596371e-11, 2.600159e-11, 2.610917e-11, 2.620612e-11, 
    2.631182e-11, 2.63377e-11, 2.64612e-11, 2.636065e-11, 2.652656e-11, 
    2.638549e-11, 2.662971e-11, 2.619095e-11, 2.638136e-11, 2.603642e-11, 
    2.607358e-11, 2.614079e-11, 2.629495e-11, 2.621173e-11, 2.630906e-11, 
    2.609409e-11, 2.598257e-11, 2.595372e-11, 2.589988e-11, 2.595495e-11, 
    2.595047e-11, 2.600316e-11, 2.598623e-11, 2.611274e-11, 2.604478e-11, 
    2.623784e-11, 2.630829e-11, 2.650728e-11, 2.662927e-11, 2.675346e-11, 
    2.680829e-11, 2.682498e-11, 2.683196e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  1.003089e-36, 2.569961e-21, 5.139921e-21, 1.798972e-20, -5.139921e-21, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, -7.709882e-21, 
    0, 2.569961e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 7.709882e-21, 1.003089e-36, 1.027984e-20, 5.139921e-21, 
    1.541976e-20, -1.28498e-20, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -1.027984e-20, 1.003089e-36, 5.139921e-21, 
    1.003089e-36, 1.027984e-20, 1.28498e-20, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, 1.28498e-20, 2.569961e-21, 
    -1.28498e-20, -2.569961e-21, -1.798972e-20, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, 1.027984e-20, -2.569961e-21, 7.709882e-21, 2.312965e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 1.28498e-20, 1.027984e-20, 
    -2.055969e-20, -7.709882e-21, 1.027984e-20, 7.709882e-21, 7.709882e-21, 
    1.541976e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, -1.28498e-20, -2.569961e-21, 0, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, -1.541976e-20, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, -2.826957e-20, 
    -5.139921e-21, 0, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, 2.569961e-21, 1.28498e-20, -2.312965e-20, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 7.709882e-21, -2.569961e-21, 1.28498e-20, -1.28498e-20, 
    5.139921e-21, 7.709882e-21, 1.798972e-20, 1.541976e-20, -2.569961e-21, 
    2.569961e-21, 2.055969e-20, 1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -2.569961e-21, 7.709882e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, 1.28498e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 2.055969e-20, 2.569961e-21, -1.541976e-20, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    1.798972e-20, -1.003089e-36, -2.055969e-20, 1.541976e-20, 5.139921e-21, 
    -1.798972e-20, -5.139921e-21, 1.541976e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -1.003089e-36, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    -1.541976e-20, 1.541976e-20, -1.798972e-20, -5.139921e-21, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -1.027984e-20, -7.709882e-21, -1.027984e-20, 
    1.027984e-20, -2.569961e-21, 1.28498e-20, -1.28498e-20, -7.709882e-21, 
    1.003089e-36, 1.28498e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -1.027984e-20, 2.569961e-21, 1.798972e-20, -7.709882e-21, 1.541976e-20, 
    -1.003089e-36, -1.28498e-20, 1.798972e-20, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, -1.28498e-20, 1.027984e-20, -5.139921e-21, 1.003089e-36, 
    -2.569961e-21, 2.569961e-21, -1.798972e-20, 7.709882e-21, 7.709882e-21, 
    -1.541976e-20, 1.798972e-20, -7.709882e-21, 5.139921e-21, -1.003089e-36, 
    1.28498e-20, -7.709882e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -1.541976e-20, 1.027984e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 
    0, 7.709882e-21, -1.541976e-20, 1.28498e-20, -7.709882e-21, 
    -5.139921e-21, -2.055969e-20, 7.709882e-21, -2.569961e-21, 1.28498e-20, 
    1.027984e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 1.28498e-20, 
    7.709882e-21, -2.055969e-20, -1.027984e-20, -1.28498e-20, -2.312965e-20, 
    5.139921e-21, -1.003089e-36, -7.709882e-21, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 1.28498e-20, 
    1.027984e-20, 5.139921e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, 1.541976e-20, -1.541976e-20, 2.569961e-21, 
    1.027984e-20, 1.541976e-20, 5.139921e-21, 5.139921e-21, -1.003089e-36, 
    -1.027984e-20, 1.003089e-36, 2.055969e-20, -7.709882e-21, 0, 0, 
    2.569961e-21, -5.139921e-21, 1.003089e-36, 1.28498e-20, 0, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, 7.709882e-21, 1.798972e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 1.003089e-36, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, -2.569961e-21, 0, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 2.055969e-20, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -1.28498e-20, 0, 1.541976e-20, 2.569961e-21,
  2.569961e-21, -1.003089e-36, 7.709882e-21, -1.027984e-20, 7.709882e-21, 
    -1.541976e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 1.003089e-36, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, -2.826957e-20, 1.28498e-20, 0, 
    0, -5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 0, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -1.28498e-20, 7.709882e-21, 1.027984e-20, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, 2.569961e-21, 
    1.027984e-20, -1.541976e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, 1.28498e-20, -7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, 0, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -1.541976e-20, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    0, -7.709882e-21, 5.139921e-21, 0, 0, 5.139921e-21, 1.003089e-36, 
    5.139921e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 0, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, -5.139921e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 1.541976e-20, -7.709882e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 0, 1.027984e-20, 1.28498e-20, -5.139921e-21, 0, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, 0, -2.569961e-21, 0, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, 0, 0, 2.569961e-21, 0, 0, 
    -2.569961e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, 1.541976e-20, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, -1.28498e-20, 
    -2.569961e-21, -1.28498e-20, -7.709882e-21, -1.798972e-20, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, 1.28498e-20, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, -2.569961e-21, -2.569961e-21, 
    0, 2.569961e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, 0, -5.139921e-21, -1.28498e-20, -7.709882e-21, 
    -1.003089e-36, 7.709882e-21, 0, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    2.569961e-21, -1.003089e-36, 5.139921e-21, 0, -2.312965e-20, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 1.027984e-20, 
    -7.709882e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, -1.027984e-20, -1.027984e-20, 0, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 0, -7.709882e-21, 
    -1.28498e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 0, 7.709882e-21, -7.709882e-21, -1.003089e-36, 
    1.541976e-20, -7.709882e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, -1.541976e-20, 
    -2.569961e-21, -2.569961e-21, 1.798972e-20, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    1.003089e-36, 7.709882e-21, 2.569961e-21, -1.027984e-20, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -5.139921e-21, 2.055969e-20, 0, 
    7.709882e-21, -1.798972e-20, 1.027984e-20, 0, 1.541976e-20, 
    -1.541976e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, 0, -1.027984e-20, 0, 0, -2.569961e-21, 0, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 5.139921e-21, 0, 
    -2.569961e-21, -7.709882e-21, -1.003089e-36, 7.709882e-21, -5.139921e-21, 
    -1.28498e-20, -1.541976e-20,
  2.569961e-21, 7.709882e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, -1.027984e-20, -2.312965e-20, -7.709882e-21, 
    -1.541976e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, 7.709882e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, 1.541976e-20, -2.569961e-21, 7.709882e-21, 
    -1.003089e-36, 0, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 0, -5.139921e-21, -2.312965e-20, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -2.055969e-20, 5.139921e-21, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, 1.541976e-20, 0, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.798972e-20, -1.003089e-36, 2.569961e-21, 
    5.139921e-21, -1.798972e-20, -7.709882e-21, -1.003089e-36, -7.709882e-21, 
    1.28498e-20, 1.28498e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 7.709882e-21, -7.709882e-21, 1.28498e-20, 
    1.027984e-20, 1.541976e-20, 1.003089e-36, 1.798972e-20, 1.027984e-20, 
    -1.003089e-36, 2.055969e-20, -7.709882e-21, -7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 7.709882e-21, 1.798972e-20, 1.541976e-20, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -2.312965e-20, -2.569961e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 
    7.709882e-21, 1.28498e-20, -2.569961e-21, 1.027984e-20, 7.709882e-21, 0, 
    -7.709882e-21, 1.003089e-36, -7.709882e-21, -7.709882e-21, 0, 
    2.312965e-20, 2.569961e-21, 1.003089e-36, -7.709882e-21, 1.003089e-36, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, -1.28498e-20, 
    -7.709882e-21, -1.027984e-20, -5.139921e-21, -1.28498e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -1.798972e-20, 1.027984e-20, 2.569961e-21, 0, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -1.798972e-20, 7.709882e-21, 0, 5.139921e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    -1.28498e-20, 0, 7.709882e-21, 0, 1.027984e-20, 0, -1.027984e-20, 
    -2.569961e-21, 0, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 7.709882e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -7.709882e-21, 1.027984e-20, -1.28498e-20, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, 0, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, -7.709882e-21, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, 1.027984e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -1.027984e-20, -1.28498e-20, -1.027984e-20, 1.28498e-20, -1.541976e-20, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.003089e-36, -2.569961e-21, 
    0, 1.28498e-20, -2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 1.541976e-20, -1.798972e-20, 
    -7.709882e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 0, 
    -1.027984e-20, 2.569961e-21, 0, 0, 1.541976e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.003089e-36, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 2.569961e-21, 2.055969e-20, 1.28498e-20, 
    1.003089e-36, -1.003089e-36, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 0, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.798972e-20, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    1.541976e-20, -1.027984e-20, 7.709882e-21, 7.709882e-21, -1.28498e-20, 
    5.139921e-21, 5.139921e-21, 1.28498e-20, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, -7.709882e-21, -1.027984e-20, 0, -5.139921e-21, 
    -7.709882e-21, 1.798972e-20, 0, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 
    1.003089e-36, -1.28498e-20, -1.003089e-36, -1.027984e-20, 0, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 0, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21,
  -1.003089e-36, -5.139921e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, -1.798972e-20, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.003089e-36, 5.139921e-21, 1.28498e-20, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 
    -1.027984e-20, 2.569961e-21, -5.139921e-21, 1.003089e-36, -7.709882e-21, 
    5.139921e-21, 1.027984e-20, -7.709882e-21, 1.798972e-20, 2.826957e-20, 
    -1.027984e-20, 2.569961e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 2.569961e-21, -5.139921e-21, -1.003089e-36, 
    2.569961e-21, -1.28498e-20, 0, 0, -1.28498e-20, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, 1.027984e-20, -1.003089e-36, 
    -2.055969e-20, -2.569961e-21, 1.003089e-36, 1.28498e-20, -7.709882e-21, 
    -5.139921e-21, 1.28498e-20, 1.541976e-20, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, 1.027984e-20, -1.28498e-20, 5.139921e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, 1.003089e-36, 7.709882e-21, -2.569961e-21, 0, 7.709882e-21, 
    2.569961e-21, 1.798972e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, -2.312965e-20, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, -1.541976e-20, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 1.541976e-20, 7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 2.055969e-20, -1.027984e-20, -1.027984e-20, -2.569961e-21, 
    -1.28498e-20, 5.139921e-21, -1.28498e-20, -5.139921e-21, -1.28498e-20, 
    7.709882e-21, -1.28498e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, -1.003089e-36, -2.312965e-20, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 
    1.28498e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, 1.798972e-20, 
    7.709882e-21, 1.003089e-36, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 7.709882e-21, -1.798972e-20, 2.569961e-21, 
    -1.28498e-20, 1.28498e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-21, 2.569961e-20, 
    -7.709882e-21, 1.027984e-20, 0, 1.027984e-20, -1.003089e-36, 
    7.709882e-21, -5.139921e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -1.798972e-20, 1.28498e-20, 0, 
    -5.139921e-21, 7.709882e-21, -1.003089e-36, -5.139921e-21, 0, 
    -7.709882e-21, 1.027984e-20, -1.28498e-20, -7.709882e-21, -1.027984e-20, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, 2.055969e-20, -1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -1.541976e-20, -1.28498e-20, -5.139921e-21, -3.083953e-20, 
    -5.139921e-21, 7.709882e-21, 7.709882e-21, -2.569961e-21, 2.055969e-20, 
    1.003089e-36, 1.541976e-20, 1.28498e-20, 0, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, 1.28498e-20, -5.139921e-21, 1.003089e-36, 
    1.027984e-20, 1.541976e-20, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    2.055969e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    1.003089e-36, 1.027984e-20, 7.709882e-21, 0, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 1.798972e-20, -2.569961e-21, 1.541976e-20, 
    1.003089e-36, 2.055969e-20, -2.569961e-21, -1.027984e-20, 0, 
    2.569961e-21, 7.709882e-21, -1.003089e-36, -1.541976e-20, 7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -7.709882e-21, 1.003089e-36, -2.569961e-21, 
    -5.139921e-21, 0, -1.28498e-20, -7.709882e-21, 7.709882e-21, 
    2.569961e-21, -1.28498e-20, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.027984e-20, 0, 1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 1.28498e-20, 
    -2.055969e-20, 5.139921e-21, 7.709882e-21, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, 2.055969e-20, 7.709882e-21, 7.709882e-21, 2.569961e-21, 
    -1.003089e-36, -1.027984e-20, 7.709882e-21, -1.003089e-36, 7.709882e-21, 
    -7.709882e-21, 1.027984e-20, 0, 1.003089e-36, 1.027984e-20, 1.798972e-20, 
    -1.027984e-20, 1.798972e-20, -2.569961e-21, 1.027984e-20, 2.055969e-20, 
    2.055969e-20, -2.055969e-20, 0, 1.541976e-20, -1.027984e-20, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -1.28498e-20,
  0, 2.569961e-21, -1.28498e-20, 7.709882e-21, -1.003089e-36, 1.798972e-20, 
    7.709882e-21, 1.541976e-20, 2.055969e-20, 7.709882e-21, 1.027984e-20, 
    2.055969e-20, -1.027984e-20, 0, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, -1.28498e-20, -2.055969e-20, 
    -7.709882e-21, 3.340949e-20, -1.541976e-20, 7.709882e-21, -1.541976e-20, 
    1.003089e-36, 1.28498e-20, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, 0, 2.569961e-20, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 1.798972e-20, 2.569961e-21, 1.003089e-36, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -5.015443e-37, -1.798972e-20, 
    -7.709882e-21, 2.569961e-21, 1.28498e-20, 2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -2.312965e-20, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, 0, -5.139921e-21, -1.798972e-20, 
    5.139921e-21, -5.139921e-21, -3.340949e-20, -5.139921e-21, -5.015443e-37, 
    1.027984e-20, 2.569961e-21, -1.798972e-20, -1.541976e-20, -7.709882e-21, 
    2.055969e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, -2.569961e-20, -1.28498e-20, 
    1.027984e-20, -7.709882e-21, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -7.709882e-21, -3.083953e-20, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, 
    -1.798972e-20, 7.709882e-21, 1.798972e-20, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, -1.003089e-36, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, 1.798972e-20, -2.826957e-20, 
    -2.826957e-20, -1.003089e-36, 5.139921e-21, -7.709882e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, -1.798972e-20, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, -1.027984e-20, 1.28498e-20, -2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -3.083953e-20, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 1.003089e-36, 5.139921e-21, -1.798972e-20, 
    5.139921e-21, 1.798972e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 1.003089e-36, -2.569961e-21, 7.709882e-21, 7.709882e-21, 
    1.798972e-20, 1.798972e-20, -7.709882e-21, 5.139921e-21, 1.798972e-20, 
    5.139921e-21, 0, -7.709882e-21, -1.003089e-36, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 0, -7.709882e-21, 1.003089e-36, 7.709882e-21, 
    1.003089e-36, 0, 1.798972e-20, -2.055969e-20, -7.709882e-21, 
    1.003089e-36, -1.798972e-20, 2.569961e-21, 2.055969e-20, 1.28498e-20, 
    -5.139921e-21, 5.139921e-21, -2.312965e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 2.569961e-21, 1.003089e-36, 2.055969e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 2.312965e-20, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, -1.798972e-20, -5.139921e-21, -2.569961e-21, 0, 
    -5.139921e-21, -1.798972e-20, 5.139921e-21, 2.569961e-21, -1.003089e-36, 
    -1.541976e-20, 1.027984e-20, -2.569961e-21, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, 2.055969e-20, 2.569961e-21, 
    1.541976e-20, -1.28498e-20, -2.312965e-20, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -2.312965e-20, -2.569961e-21, 
    -7.709882e-21, 1.541976e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, -1.003089e-36, 1.027984e-20, 
    1.003089e-36, -1.798972e-20, 2.312965e-20, -2.569961e-21, 0, 
    -1.003089e-36, 1.541976e-20, 1.003089e-36, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -1.003089e-36, -1.003089e-36, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, -2.569961e-21, 
    -2.569961e-20, 7.709882e-21, 1.541976e-20, -1.541976e-20, 7.709882e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, 2.312965e-20, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, 1.003089e-36, 7.709882e-21, 1.28498e-20, 
    1.28498e-20, -1.541976e-20, -7.709882e-21, 2.055969e-20, -1.798972e-20, 
    7.709882e-21, -2.569961e-21, -2.055969e-20, 7.709882e-21, -5.139921e-21, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, 1.798972e-20, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.798972e-20, 1.003089e-36, -2.569961e-21, 
    -5.139921e-21, -1.027984e-20, 7.709882e-21, 1.541976e-20, 1.003089e-36, 
    1.027984e-20, 5.139921e-21, 2.569961e-21, 0, 1.28498e-20, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -2.569961e-21, 1.541976e-20, -5.139921e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, -2.055969e-20,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.149711e-12, 5.172433e-12, 5.168016e-12, 5.186343e-12, 5.176177e-12, 
    5.188177e-12, 5.154318e-12, 5.173334e-12, 5.161195e-12, 5.151757e-12, 
    5.221908e-12, 5.18716e-12, 5.258011e-12, 5.235847e-12, 5.291529e-12, 
    5.254562e-12, 5.298983e-12, 5.290463e-12, 5.31611e-12, 5.308763e-12, 
    5.341564e-12, 5.319501e-12, 5.358571e-12, 5.336296e-12, 5.33978e-12, 
    5.318773e-12, 5.194154e-12, 5.217582e-12, 5.192766e-12, 5.196107e-12, 
    5.194608e-12, 5.176386e-12, 5.167203e-12, 5.147976e-12, 5.151466e-12, 
    5.165589e-12, 5.197609e-12, 5.18674e-12, 5.214135e-12, 5.213516e-12, 
    5.244016e-12, 5.230264e-12, 5.281531e-12, 5.26696e-12, 5.309069e-12, 
    5.298478e-12, 5.308571e-12, 5.305511e-12, 5.308611e-12, 5.293079e-12, 
    5.299734e-12, 5.286067e-12, 5.232839e-12, 5.248481e-12, 5.20183e-12, 
    5.173779e-12, 5.155152e-12, 5.141934e-12, 5.143802e-12, 5.147365e-12, 
    5.165672e-12, 5.182886e-12, 5.196005e-12, 5.20478e-12, 5.213427e-12, 
    5.239598e-12, 5.253454e-12, 5.284477e-12, 5.278879e-12, 5.288363e-12, 
    5.297425e-12, 5.312638e-12, 5.310134e-12, 5.316836e-12, 5.288114e-12, 
    5.307202e-12, 5.27569e-12, 5.284309e-12, 5.215774e-12, 5.189672e-12, 
    5.178575e-12, 5.168865e-12, 5.145239e-12, 5.161554e-12, 5.155122e-12, 
    5.170425e-12, 5.180148e-12, 5.175339e-12, 5.20502e-12, 5.193481e-12, 
    5.254275e-12, 5.228088e-12, 5.296368e-12, 5.280028e-12, 5.300285e-12, 
    5.289948e-12, 5.307659e-12, 5.291719e-12, 5.319331e-12, 5.325344e-12, 
    5.321235e-12, 5.337019e-12, 5.290836e-12, 5.308571e-12, 5.175204e-12, 
    5.175989e-12, 5.179643e-12, 5.163581e-12, 5.162598e-12, 5.14788e-12, 
    5.160976e-12, 5.166553e-12, 5.180712e-12, 5.189087e-12, 5.197048e-12, 
    5.214553e-12, 5.234103e-12, 5.261443e-12, 5.281087e-12, 5.294255e-12, 
    5.286181e-12, 5.293309e-12, 5.28534e-12, 5.281606e-12, 5.32309e-12, 
    5.299795e-12, 5.334749e-12, 5.332815e-12, 5.316996e-12, 5.333033e-12, 
    5.176539e-12, 5.172026e-12, 5.156356e-12, 5.168619e-12, 5.146277e-12, 
    5.158783e-12, 5.165973e-12, 5.193721e-12, 5.199819e-12, 5.205472e-12, 
    5.216638e-12, 5.230968e-12, 5.256107e-12, 5.277981e-12, 5.297952e-12, 
    5.296489e-12, 5.297004e-12, 5.301465e-12, 5.290414e-12, 5.30328e-12, 
    5.305438e-12, 5.299793e-12, 5.332556e-12, 5.323196e-12, 5.332774e-12, 
    5.32668e-12, 5.173494e-12, 5.181088e-12, 5.176984e-12, 5.184701e-12, 
    5.179264e-12, 5.203438e-12, 5.210686e-12, 5.244605e-12, 5.230685e-12, 
    5.25284e-12, 5.232936e-12, 5.236462e-12, 5.253561e-12, 5.234012e-12, 
    5.276774e-12, 5.247781e-12, 5.301638e-12, 5.272682e-12, 5.303453e-12, 
    5.297866e-12, 5.307117e-12, 5.315402e-12, 5.325826e-12, 5.34506e-12, 
    5.340606e-12, 5.356692e-12, 5.19241e-12, 5.20226e-12, 5.201394e-12, 
    5.211703e-12, 5.219327e-12, 5.235853e-12, 5.26236e-12, 5.252392e-12, 
    5.270692e-12, 5.274365e-12, 5.246564e-12, 5.263632e-12, 5.208853e-12, 
    5.217702e-12, 5.212434e-12, 5.193187e-12, 5.254688e-12, 5.223124e-12, 
    5.281412e-12, 5.264311e-12, 5.31422e-12, 5.289398e-12, 5.338154e-12, 
    5.358997e-12, 5.378617e-12, 5.401543e-12, 5.207637e-12, 5.200943e-12, 
    5.212929e-12, 5.22951e-12, 5.244897e-12, 5.265354e-12, 5.267448e-12, 
    5.27128e-12, 5.281207e-12, 5.289554e-12, 5.272491e-12, 5.291647e-12, 
    5.219753e-12, 5.257428e-12, 5.198412e-12, 5.216181e-12, 5.228533e-12, 
    5.223115e-12, 5.251253e-12, 5.257885e-12, 5.284834e-12, 5.270903e-12, 
    5.353851e-12, 5.317151e-12, 5.419002e-12, 5.390537e-12, 5.198605e-12, 
    5.207614e-12, 5.238969e-12, 5.22405e-12, 5.26672e-12, 5.277224e-12, 
    5.285763e-12, 5.296678e-12, 5.297857e-12, 5.304324e-12, 5.293726e-12, 
    5.303905e-12, 5.265397e-12, 5.282606e-12, 5.235386e-12, 5.246878e-12, 
    5.241592e-12, 5.235793e-12, 5.253691e-12, 5.272759e-12, 5.273168e-12, 
    5.279282e-12, 5.29651e-12, 5.266893e-12, 5.358586e-12, 5.301955e-12, 
    5.217438e-12, 5.23479e-12, 5.237271e-12, 5.230549e-12, 5.27617e-12, 
    5.259639e-12, 5.304166e-12, 5.292132e-12, 5.31185e-12, 5.302052e-12, 
    5.30061e-12, 5.288026e-12, 5.280191e-12, 5.260397e-12, 5.244293e-12, 
    5.231524e-12, 5.234493e-12, 5.24852e-12, 5.273926e-12, 5.297963e-12, 
    5.292697e-12, 5.310352e-12, 5.263626e-12, 5.283218e-12, 5.275645e-12, 
    5.295391e-12, 5.252127e-12, 5.288965e-12, 5.242711e-12, 5.246766e-12, 
    5.259311e-12, 5.284546e-12, 5.290131e-12, 5.296092e-12, 5.292414e-12, 
    5.274571e-12, 5.271649e-12, 5.259006e-12, 5.255515e-12, 5.245884e-12, 
    5.237909e-12, 5.245194e-12, 5.252846e-12, 5.274579e-12, 5.294165e-12, 
    5.31552e-12, 5.320746e-12, 5.345696e-12, 5.325384e-12, 5.358902e-12, 
    5.330403e-12, 5.379738e-12, 5.291102e-12, 5.329567e-12, 5.259882e-12, 
    5.267389e-12, 5.280967e-12, 5.312111e-12, 5.295298e-12, 5.314962e-12, 
    5.271534e-12, 5.249003e-12, 5.243175e-12, 5.2323e-12, 5.243424e-12, 
    5.242519e-12, 5.253164e-12, 5.249743e-12, 5.275301e-12, 5.261572e-12, 
    5.300574e-12, 5.314807e-12, 5.355006e-12, 5.37965e-12, 5.40474e-12, 
    5.415816e-12, 5.419188e-12, 5.420597e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.115576e-11, 3.129322e-11, 3.12665e-11, 3.137737e-11, 3.131587e-11, 
    3.138847e-11, 3.118363e-11, 3.129867e-11, 3.122523e-11, 3.116813e-11, 
    3.159254e-11, 3.138232e-11, 3.181097e-11, 3.167687e-11, 3.201375e-11, 
    3.179009e-11, 3.205885e-11, 3.20073e-11, 3.216246e-11, 3.211801e-11, 
    3.231647e-11, 3.218298e-11, 3.241936e-11, 3.228459e-11, 3.230567e-11, 
    3.217858e-11, 3.142463e-11, 3.156637e-11, 3.141623e-11, 3.143644e-11, 
    3.142738e-11, 3.131714e-11, 3.126158e-11, 3.114525e-11, 3.116637e-11, 
    3.125181e-11, 3.144553e-11, 3.137978e-11, 3.154552e-11, 3.154177e-11, 
    3.17263e-11, 3.164309e-11, 3.195326e-11, 3.18651e-11, 3.211987e-11, 
    3.20558e-11, 3.211686e-11, 3.209834e-11, 3.21171e-11, 3.202313e-11, 
    3.206339e-11, 3.19807e-11, 3.165868e-11, 3.175331e-11, 3.147107e-11, 
    3.130136e-11, 3.118867e-11, 3.11087e-11, 3.112001e-11, 3.114155e-11, 
    3.125232e-11, 3.135646e-11, 3.143583e-11, 3.148892e-11, 3.154123e-11, 
    3.169957e-11, 3.17834e-11, 3.197109e-11, 3.193722e-11, 3.199459e-11, 
    3.204942e-11, 3.214146e-11, 3.212631e-11, 3.216686e-11, 3.199309e-11, 
    3.210857e-11, 3.191793e-11, 3.197007e-11, 3.155543e-11, 3.139752e-11, 
    3.133038e-11, 3.127163e-11, 3.11287e-11, 3.12274e-11, 3.118849e-11, 
    3.128107e-11, 3.13399e-11, 3.13108e-11, 3.149037e-11, 3.142056e-11, 
    3.178836e-11, 3.162993e-11, 3.204302e-11, 3.194417e-11, 3.206672e-11, 
    3.200419e-11, 3.211133e-11, 3.20149e-11, 3.218196e-11, 3.221833e-11, 
    3.219347e-11, 3.228897e-11, 3.200956e-11, 3.211685e-11, 3.130999e-11, 
    3.131473e-11, 3.133684e-11, 3.123966e-11, 3.123372e-11, 3.114467e-11, 
    3.122391e-11, 3.125765e-11, 3.134331e-11, 3.139397e-11, 3.144214e-11, 
    3.154805e-11, 3.166632e-11, 3.183173e-11, 3.195058e-11, 3.203024e-11, 
    3.19814e-11, 3.202452e-11, 3.197631e-11, 3.195371e-11, 3.22047e-11, 
    3.206376e-11, 3.227523e-11, 3.226353e-11, 3.216782e-11, 3.226485e-11, 
    3.131806e-11, 3.129076e-11, 3.119596e-11, 3.127015e-11, 3.113498e-11, 
    3.121063e-11, 3.125414e-11, 3.142201e-11, 3.14589e-11, 3.14931e-11, 
    3.156066e-11, 3.164735e-11, 3.179945e-11, 3.193179e-11, 3.205261e-11, 
    3.204376e-11, 3.204688e-11, 3.207386e-11, 3.200701e-11, 3.208484e-11, 
    3.20979e-11, 3.206375e-11, 3.226196e-11, 3.220534e-11, 3.226328e-11, 
    3.222641e-11, 3.129964e-11, 3.134558e-11, 3.132075e-11, 3.136744e-11, 
    3.133455e-11, 3.14808e-11, 3.152465e-11, 3.172986e-11, 3.164564e-11, 
    3.177968e-11, 3.165926e-11, 3.16806e-11, 3.178404e-11, 3.166577e-11, 
    3.192448e-11, 3.174907e-11, 3.207491e-11, 3.189973e-11, 3.208589e-11, 
    3.205209e-11, 3.210806e-11, 3.215818e-11, 3.222125e-11, 3.233761e-11, 
    3.231067e-11, 3.240799e-11, 3.141408e-11, 3.147367e-11, 3.146843e-11, 
    3.15308e-11, 3.157693e-11, 3.167691e-11, 3.183728e-11, 3.177697e-11, 
    3.188769e-11, 3.190991e-11, 3.174171e-11, 3.184498e-11, 3.151356e-11, 
    3.15671e-11, 3.153523e-11, 3.141878e-11, 3.179086e-11, 3.15999e-11, 
    3.195254e-11, 3.184908e-11, 3.215104e-11, 3.200086e-11, 3.229583e-11, 
    3.242193e-11, 3.254063e-11, 3.267933e-11, 3.15062e-11, 3.146571e-11, 
    3.153822e-11, 3.163854e-11, 3.173163e-11, 3.185539e-11, 3.186806e-11, 
    3.189124e-11, 3.195131e-11, 3.20018e-11, 3.189857e-11, 3.201446e-11, 
    3.157951e-11, 3.180744e-11, 3.145039e-11, 3.15579e-11, 3.163262e-11, 
    3.159985e-11, 3.177008e-11, 3.18102e-11, 3.197325e-11, 3.188896e-11, 
    3.23908e-11, 3.216876e-11, 3.278497e-11, 3.261275e-11, 3.145156e-11, 
    3.150607e-11, 3.169577e-11, 3.160551e-11, 3.186366e-11, 3.19272e-11, 
    3.197886e-11, 3.20449e-11, 3.205203e-11, 3.209116e-11, 3.202704e-11, 
    3.208863e-11, 3.185566e-11, 3.195976e-11, 3.167409e-11, 3.174361e-11, 
    3.171163e-11, 3.167655e-11, 3.178483e-11, 3.190019e-11, 3.190266e-11, 
    3.193966e-11, 3.204388e-11, 3.18647e-11, 3.241945e-11, 3.207682e-11, 
    3.15655e-11, 3.167048e-11, 3.168549e-11, 3.164482e-11, 3.192083e-11, 
    3.182082e-11, 3.209021e-11, 3.20174e-11, 3.21367e-11, 3.207741e-11, 
    3.206869e-11, 3.199256e-11, 3.194515e-11, 3.18254e-11, 3.172797e-11, 
    3.165072e-11, 3.166868e-11, 3.175354e-11, 3.190725e-11, 3.205267e-11, 
    3.202082e-11, 3.212763e-11, 3.184494e-11, 3.196347e-11, 3.191765e-11, 
    3.203712e-11, 3.177537e-11, 3.199824e-11, 3.17184e-11, 3.174293e-11, 
    3.181883e-11, 3.19715e-11, 3.200529e-11, 3.204136e-11, 3.20191e-11, 
    3.191115e-11, 3.189347e-11, 3.181699e-11, 3.179587e-11, 3.17376e-11, 
    3.168935e-11, 3.173343e-11, 3.177972e-11, 3.19112e-11, 3.20297e-11, 
    3.215889e-11, 3.219052e-11, 3.234146e-11, 3.221858e-11, 3.242135e-11, 
    3.224894e-11, 3.254742e-11, 3.201116e-11, 3.224388e-11, 3.182229e-11, 
    3.186771e-11, 3.194985e-11, 3.213827e-11, 3.203656e-11, 3.215552e-11, 
    3.189278e-11, 3.175647e-11, 3.172121e-11, 3.165541e-11, 3.172271e-11, 
    3.171724e-11, 3.178164e-11, 3.176094e-11, 3.191557e-11, 3.183251e-11, 
    3.206847e-11, 3.215458e-11, 3.239779e-11, 3.254688e-11, 3.269867e-11, 
    3.276569e-11, 3.278609e-11, 3.279461e-11 ;

 SOILC =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 SOILC_HR =
  6.190983e-08, 6.218286e-08, 6.212978e-08, 6.234999e-08, 6.222784e-08, 
    6.237203e-08, 6.196519e-08, 6.219368e-08, 6.204782e-08, 6.193441e-08, 
    6.277735e-08, 6.235982e-08, 6.321117e-08, 6.294484e-08, 6.361391e-08, 
    6.316971e-08, 6.370349e-08, 6.360111e-08, 6.390928e-08, 6.382099e-08, 
    6.421514e-08, 6.395003e-08, 6.44195e-08, 6.415184e-08, 6.41937e-08, 
    6.394128e-08, 6.244386e-08, 6.272536e-08, 6.242718e-08, 6.246731e-08, 
    6.244931e-08, 6.223036e-08, 6.212002e-08, 6.188898e-08, 6.193092e-08, 
    6.210062e-08, 6.248537e-08, 6.235477e-08, 6.268395e-08, 6.267651e-08, 
    6.3043e-08, 6.287775e-08, 6.349378e-08, 6.331869e-08, 6.382468e-08, 
    6.369742e-08, 6.38187e-08, 6.378193e-08, 6.381918e-08, 6.363254e-08, 
    6.371251e-08, 6.354828e-08, 6.29087e-08, 6.309665e-08, 6.253609e-08, 
    6.219904e-08, 6.197521e-08, 6.181637e-08, 6.183883e-08, 6.188163e-08, 
    6.210161e-08, 6.230846e-08, 6.246609e-08, 6.257154e-08, 6.267544e-08, 
    6.298992e-08, 6.315641e-08, 6.352918e-08, 6.346192e-08, 6.357588e-08, 
    6.368477e-08, 6.386757e-08, 6.383748e-08, 6.391802e-08, 6.357288e-08, 
    6.380225e-08, 6.34236e-08, 6.352716e-08, 6.270364e-08, 6.239001e-08, 
    6.225666e-08, 6.213998e-08, 6.185609e-08, 6.205214e-08, 6.197485e-08, 
    6.215873e-08, 6.227556e-08, 6.221778e-08, 6.257442e-08, 6.243577e-08, 
    6.316627e-08, 6.28516e-08, 6.367206e-08, 6.347572e-08, 6.371913e-08, 
    6.359492e-08, 6.380773e-08, 6.361621e-08, 6.394799e-08, 6.402023e-08, 
    6.397087e-08, 6.416053e-08, 6.360559e-08, 6.38187e-08, 6.221616e-08, 
    6.222558e-08, 6.226949e-08, 6.207648e-08, 6.206467e-08, 6.188782e-08, 
    6.204519e-08, 6.21122e-08, 6.228234e-08, 6.238297e-08, 6.247863e-08, 
    6.268897e-08, 6.292388e-08, 6.325241e-08, 6.348845e-08, 6.364667e-08, 
    6.354966e-08, 6.363531e-08, 6.353956e-08, 6.349468e-08, 6.399316e-08, 
    6.371325e-08, 6.413325e-08, 6.411001e-08, 6.391993e-08, 6.411263e-08, 
    6.22322e-08, 6.217797e-08, 6.198967e-08, 6.213703e-08, 6.186856e-08, 
    6.201883e-08, 6.210523e-08, 6.243865e-08, 6.251192e-08, 6.257985e-08, 
    6.271402e-08, 6.288621e-08, 6.318828e-08, 6.345113e-08, 6.36911e-08, 
    6.367352e-08, 6.367971e-08, 6.373331e-08, 6.360052e-08, 6.375511e-08, 
    6.378105e-08, 6.371322e-08, 6.41069e-08, 6.399443e-08, 6.410952e-08, 
    6.403629e-08, 6.21956e-08, 6.228685e-08, 6.223754e-08, 6.233027e-08, 
    6.226494e-08, 6.255542e-08, 6.264251e-08, 6.305007e-08, 6.288282e-08, 
    6.314902e-08, 6.290986e-08, 6.295224e-08, 6.315769e-08, 6.292279e-08, 
    6.343662e-08, 6.308824e-08, 6.373539e-08, 6.338745e-08, 6.37572e-08, 
    6.369006e-08, 6.380122e-08, 6.390078e-08, 6.402603e-08, 6.425714e-08, 
    6.420363e-08, 6.439692e-08, 6.24229e-08, 6.254125e-08, 6.253084e-08, 
    6.265472e-08, 6.274633e-08, 6.294491e-08, 6.326341e-08, 6.314364e-08, 
    6.336354e-08, 6.340768e-08, 6.307361e-08, 6.327871e-08, 6.262048e-08, 
    6.272681e-08, 6.266351e-08, 6.243223e-08, 6.317123e-08, 6.279195e-08, 
    6.349235e-08, 6.328687e-08, 6.388658e-08, 6.358832e-08, 6.417417e-08, 
    6.442461e-08, 6.466037e-08, 6.493585e-08, 6.260586e-08, 6.252544e-08, 
    6.266945e-08, 6.286869e-08, 6.305359e-08, 6.32994e-08, 6.332456e-08, 
    6.33706e-08, 6.348989e-08, 6.359019e-08, 6.338515e-08, 6.361533e-08, 
    6.275145e-08, 6.320415e-08, 6.249503e-08, 6.270854e-08, 6.285696e-08, 
    6.279186e-08, 6.312996e-08, 6.320965e-08, 6.353348e-08, 6.336608e-08, 
    6.436279e-08, 6.39218e-08, 6.514564e-08, 6.480359e-08, 6.249734e-08, 
    6.260559e-08, 6.298236e-08, 6.28031e-08, 6.331581e-08, 6.344202e-08, 
    6.354463e-08, 6.367578e-08, 6.368995e-08, 6.376766e-08, 6.364031e-08, 
    6.376263e-08, 6.329992e-08, 6.35067e-08, 6.293931e-08, 6.307739e-08, 
    6.301387e-08, 6.294419e-08, 6.315926e-08, 6.338838e-08, 6.339329e-08, 
    6.346676e-08, 6.367377e-08, 6.331789e-08, 6.441968e-08, 6.373919e-08, 
    6.272364e-08, 6.293214e-08, 6.296194e-08, 6.288117e-08, 6.342937e-08, 
    6.323073e-08, 6.376577e-08, 6.362117e-08, 6.38581e-08, 6.374036e-08, 
    6.372304e-08, 6.357183e-08, 6.347768e-08, 6.323983e-08, 6.304632e-08, 
    6.289289e-08, 6.292857e-08, 6.309711e-08, 6.34024e-08, 6.369122e-08, 
    6.362795e-08, 6.384009e-08, 6.327863e-08, 6.351405e-08, 6.342306e-08, 
    6.366032e-08, 6.314046e-08, 6.358311e-08, 6.302731e-08, 6.307604e-08, 
    6.322679e-08, 6.353001e-08, 6.359712e-08, 6.366874e-08, 6.362455e-08, 
    6.341015e-08, 6.337503e-08, 6.322313e-08, 6.318118e-08, 6.306544e-08, 
    6.296961e-08, 6.305716e-08, 6.31491e-08, 6.341025e-08, 6.364559e-08, 
    6.390219e-08, 6.3965e-08, 6.426479e-08, 6.402072e-08, 6.442347e-08, 
    6.408103e-08, 6.467384e-08, 6.360878e-08, 6.407099e-08, 6.323365e-08, 
    6.332385e-08, 6.3487e-08, 6.386124e-08, 6.365921e-08, 6.389548e-08, 
    6.337365e-08, 6.310292e-08, 6.303289e-08, 6.290222e-08, 6.303588e-08, 
    6.302501e-08, 6.315292e-08, 6.311182e-08, 6.341892e-08, 6.325396e-08, 
    6.37226e-08, 6.389362e-08, 6.437666e-08, 6.467278e-08, 6.497426e-08, 
    6.510736e-08, 6.514787e-08, 6.516481e-08 ;

 SOILC_LOSS =
  6.190983e-08, 6.218286e-08, 6.212978e-08, 6.234999e-08, 6.222784e-08, 
    6.237203e-08, 6.196519e-08, 6.219368e-08, 6.204782e-08, 6.193441e-08, 
    6.277735e-08, 6.235982e-08, 6.321117e-08, 6.294484e-08, 6.361391e-08, 
    6.316971e-08, 6.370349e-08, 6.360111e-08, 6.390928e-08, 6.382099e-08, 
    6.421514e-08, 6.395003e-08, 6.44195e-08, 6.415184e-08, 6.41937e-08, 
    6.394128e-08, 6.244386e-08, 6.272536e-08, 6.242718e-08, 6.246731e-08, 
    6.244931e-08, 6.223036e-08, 6.212002e-08, 6.188898e-08, 6.193092e-08, 
    6.210062e-08, 6.248537e-08, 6.235477e-08, 6.268395e-08, 6.267651e-08, 
    6.3043e-08, 6.287775e-08, 6.349378e-08, 6.331869e-08, 6.382468e-08, 
    6.369742e-08, 6.38187e-08, 6.378193e-08, 6.381918e-08, 6.363254e-08, 
    6.371251e-08, 6.354828e-08, 6.29087e-08, 6.309665e-08, 6.253609e-08, 
    6.219904e-08, 6.197521e-08, 6.181637e-08, 6.183883e-08, 6.188163e-08, 
    6.210161e-08, 6.230846e-08, 6.246609e-08, 6.257154e-08, 6.267544e-08, 
    6.298992e-08, 6.315641e-08, 6.352918e-08, 6.346192e-08, 6.357588e-08, 
    6.368477e-08, 6.386757e-08, 6.383748e-08, 6.391802e-08, 6.357288e-08, 
    6.380225e-08, 6.34236e-08, 6.352716e-08, 6.270364e-08, 6.239001e-08, 
    6.225666e-08, 6.213998e-08, 6.185609e-08, 6.205214e-08, 6.197485e-08, 
    6.215873e-08, 6.227556e-08, 6.221778e-08, 6.257442e-08, 6.243577e-08, 
    6.316627e-08, 6.28516e-08, 6.367206e-08, 6.347572e-08, 6.371913e-08, 
    6.359492e-08, 6.380773e-08, 6.361621e-08, 6.394799e-08, 6.402023e-08, 
    6.397087e-08, 6.416053e-08, 6.360559e-08, 6.38187e-08, 6.221616e-08, 
    6.222558e-08, 6.226949e-08, 6.207648e-08, 6.206467e-08, 6.188782e-08, 
    6.204519e-08, 6.21122e-08, 6.228234e-08, 6.238297e-08, 6.247863e-08, 
    6.268897e-08, 6.292388e-08, 6.325241e-08, 6.348845e-08, 6.364667e-08, 
    6.354966e-08, 6.363531e-08, 6.353956e-08, 6.349468e-08, 6.399316e-08, 
    6.371325e-08, 6.413325e-08, 6.411001e-08, 6.391993e-08, 6.411263e-08, 
    6.22322e-08, 6.217797e-08, 6.198967e-08, 6.213703e-08, 6.186856e-08, 
    6.201883e-08, 6.210523e-08, 6.243865e-08, 6.251192e-08, 6.257985e-08, 
    6.271402e-08, 6.288621e-08, 6.318828e-08, 6.345113e-08, 6.36911e-08, 
    6.367352e-08, 6.367971e-08, 6.373331e-08, 6.360052e-08, 6.375511e-08, 
    6.378105e-08, 6.371322e-08, 6.41069e-08, 6.399443e-08, 6.410952e-08, 
    6.403629e-08, 6.21956e-08, 6.228685e-08, 6.223754e-08, 6.233027e-08, 
    6.226494e-08, 6.255542e-08, 6.264251e-08, 6.305007e-08, 6.288282e-08, 
    6.314902e-08, 6.290986e-08, 6.295224e-08, 6.315769e-08, 6.292279e-08, 
    6.343662e-08, 6.308824e-08, 6.373539e-08, 6.338745e-08, 6.37572e-08, 
    6.369006e-08, 6.380122e-08, 6.390078e-08, 6.402603e-08, 6.425714e-08, 
    6.420363e-08, 6.439692e-08, 6.24229e-08, 6.254125e-08, 6.253084e-08, 
    6.265472e-08, 6.274633e-08, 6.294491e-08, 6.326341e-08, 6.314364e-08, 
    6.336354e-08, 6.340768e-08, 6.307361e-08, 6.327871e-08, 6.262048e-08, 
    6.272681e-08, 6.266351e-08, 6.243223e-08, 6.317123e-08, 6.279195e-08, 
    6.349235e-08, 6.328687e-08, 6.388658e-08, 6.358832e-08, 6.417417e-08, 
    6.442461e-08, 6.466037e-08, 6.493585e-08, 6.260586e-08, 6.252544e-08, 
    6.266945e-08, 6.286869e-08, 6.305359e-08, 6.32994e-08, 6.332456e-08, 
    6.33706e-08, 6.348989e-08, 6.359019e-08, 6.338515e-08, 6.361533e-08, 
    6.275145e-08, 6.320415e-08, 6.249503e-08, 6.270854e-08, 6.285696e-08, 
    6.279186e-08, 6.312996e-08, 6.320965e-08, 6.353348e-08, 6.336608e-08, 
    6.436279e-08, 6.39218e-08, 6.514564e-08, 6.480359e-08, 6.249734e-08, 
    6.260559e-08, 6.298236e-08, 6.28031e-08, 6.331581e-08, 6.344202e-08, 
    6.354463e-08, 6.367578e-08, 6.368995e-08, 6.376766e-08, 6.364031e-08, 
    6.376263e-08, 6.329992e-08, 6.35067e-08, 6.293931e-08, 6.307739e-08, 
    6.301387e-08, 6.294419e-08, 6.315926e-08, 6.338838e-08, 6.339329e-08, 
    6.346676e-08, 6.367377e-08, 6.331789e-08, 6.441968e-08, 6.373919e-08, 
    6.272364e-08, 6.293214e-08, 6.296194e-08, 6.288117e-08, 6.342937e-08, 
    6.323073e-08, 6.376577e-08, 6.362117e-08, 6.38581e-08, 6.374036e-08, 
    6.372304e-08, 6.357183e-08, 6.347768e-08, 6.323983e-08, 6.304632e-08, 
    6.289289e-08, 6.292857e-08, 6.309711e-08, 6.34024e-08, 6.369122e-08, 
    6.362795e-08, 6.384009e-08, 6.327863e-08, 6.351405e-08, 6.342306e-08, 
    6.366032e-08, 6.314046e-08, 6.358311e-08, 6.302731e-08, 6.307604e-08, 
    6.322679e-08, 6.353001e-08, 6.359712e-08, 6.366874e-08, 6.362455e-08, 
    6.341015e-08, 6.337503e-08, 6.322313e-08, 6.318118e-08, 6.306544e-08, 
    6.296961e-08, 6.305716e-08, 6.31491e-08, 6.341025e-08, 6.364559e-08, 
    6.390219e-08, 6.3965e-08, 6.426479e-08, 6.402072e-08, 6.442347e-08, 
    6.408103e-08, 6.467384e-08, 6.360878e-08, 6.407099e-08, 6.323365e-08, 
    6.332385e-08, 6.3487e-08, 6.386124e-08, 6.365921e-08, 6.389548e-08, 
    6.337365e-08, 6.310292e-08, 6.303289e-08, 6.290222e-08, 6.303588e-08, 
    6.302501e-08, 6.315292e-08, 6.311182e-08, 6.341892e-08, 6.325396e-08, 
    6.37226e-08, 6.389362e-08, 6.437666e-08, 6.467278e-08, 6.497426e-08, 
    6.510736e-08, 6.514787e-08, 6.516481e-08 ;

 SOILICE =
  94.68816, 95.13689, 95.04955, 95.41229, 95.21095, 95.44865, 94.77901, 
    95.15474, 94.91476, 94.72849, 96.11891, 95.4285, 96.8395, 96.39663, 
    97.51165, 96.77051, 97.66153, 97.4902, 98.00642, 97.85835, 98.52058, 
    98.07481, 98.86496, 98.41399, 98.48446, 98.06012, 95.56716, 96.03278, 
    95.53962, 95.60591, 95.57616, 95.21511, 95.03352, 94.65391, 94.72275, 
    95.00159, 95.63573, 95.42014, 95.96407, 95.95177, 96.55968, 96.28527, 
    97.31081, 97.0186, 97.86452, 97.65134, 97.85451, 97.79287, 97.85531, 
    97.54277, 97.6766, 97.40187, 96.33663, 96.6489, 95.71952, 95.16358, 
    94.79547, 94.53485, 94.57167, 94.64188, 95.00322, 95.34379, 95.60387, 
    95.77811, 95.95, 96.47157, 96.74834, 97.36996, 97.25758, 97.44801, 
    97.63015, 97.93645, 97.88599, 98.0211, 97.44298, 97.82695, 97.1936, 
    97.36656, 95.99682, 95.47827, 95.25848, 95.06633, 94.59998, 94.92188, 
    94.79489, 95.09716, 95.28956, 95.19437, 95.78288, 95.55379, 96.76476, 
    96.24192, 97.60889, 97.28064, 97.68768, 97.47984, 97.83614, 97.51543, 
    98.0714, 98.19274, 98.10981, 98.4286, 97.49767, 97.85452, 95.1917, 
    95.20722, 95.27955, 94.96189, 94.94248, 94.65202, 94.91044, 95.02063, 
    95.30072, 95.46666, 95.62458, 95.9724, 96.36185, 96.90817, 97.3019, 
    97.5664, 97.40415, 97.54739, 97.38728, 97.31229, 98.14727, 97.67785, 
    98.38271, 98.34361, 98.02431, 98.34801, 95.21812, 95.12882, 94.81923, 
    95.06145, 94.62043, 94.86713, 95.00919, 95.55859, 95.67957, 95.79186, 
    96.01387, 96.2993, 96.80137, 97.23959, 97.64075, 97.61132, 97.62168, 
    97.71143, 97.4892, 97.74795, 97.79143, 97.67779, 98.33838, 98.14936, 
    98.34278, 98.21968, 95.15784, 95.30817, 95.22691, 95.37974, 95.27206, 
    95.75149, 95.89554, 96.57149, 96.29369, 96.73604, 96.33855, 96.40891, 
    96.75052, 96.36, 97.2154, 96.63495, 97.71493, 97.13336, 97.75144, 
    97.63901, 97.8252, 97.99216, 98.20246, 98.59126, 98.50114, 98.82684, 
    95.53255, 95.72807, 95.71084, 95.9157, 96.0674, 96.39673, 96.92649, 
    96.72705, 97.09339, 97.16705, 96.61057, 96.952, 95.85906, 96.0351, 
    95.93025, 95.54797, 96.773, 96.14303, 97.30841, 96.96557, 97.96835, 
    97.46883, 98.45155, 98.87362, 99.27184, 99.73857, 95.83488, 95.7019, 
    95.94008, 96.27028, 96.57729, 96.98646, 97.02838, 97.10518, 97.3043, 
    97.47192, 97.12949, 97.51397, 96.07598, 96.8278, 95.65166, 96.00484, 
    96.25079, 96.14284, 96.70427, 96.83691, 97.37714, 97.09763, 98.76936, 
    98.02747, 100.0948, 99.51434, 95.65547, 95.83442, 96.45895, 96.16146, 
    97.01381, 97.22437, 97.39575, 97.61514, 97.63882, 97.76898, 97.55576, 
    97.76055, 96.98733, 97.33237, 96.38741, 96.61686, 96.51126, 96.39552, 
    96.75302, 97.13487, 97.14303, 97.26569, 97.6119, 97.01727, 98.8654, 
    97.72142, 96.0298, 96.3756, 96.42503, 96.29094, 97.20325, 96.87203, 
    97.76581, 97.52372, 97.92057, 97.72324, 97.69423, 97.44121, 97.28391, 
    96.88721, 96.56522, 96.31038, 96.36959, 96.64967, 97.15826, 97.64098, 
    97.53511, 97.89037, 96.95184, 97.34468, 97.19273, 97.58925, 96.72176, 
    97.46022, 96.5336, 96.61461, 96.86547, 97.37138, 97.48351, 97.60336, 
    97.52939, 97.17119, 97.11258, 96.85936, 96.78954, 96.59697, 96.43774, 
    96.58321, 96.73615, 97.17133, 97.56461, 97.99454, 98.09994, 98.60422, 
    98.19361, 98.8718, 98.29507, 99.29477, 97.50309, 98.2781, 96.87688, 
    97.02721, 97.29951, 97.92588, 97.58739, 97.98332, 97.11028, 96.65935, 
    96.54288, 96.32586, 96.54784, 96.52978, 96.74248, 96.6741, 97.18581, 
    96.91071, 97.6935, 97.98019, 98.79268, 99.29288, 99.80368, 100.0297, 
    100.0986, 100.1274,
  94.56142, 95.02821, 94.93734, 95.31439, 95.10522, 95.35104, 94.65591, 
    95.04681, 94.79713, 94.60334, 96.02686, 95.33073, 96.75284, 96.30653, 
    97.42994, 96.68336, 97.58088, 97.40825, 97.92813, 97.77901, 98.44598, 
    97.99699, 98.79263, 98.3386, 98.40958, 97.98222, 95.47047, 95.94005, 
    95.44272, 95.50957, 95.47955, 95.10957, 94.92075, 94.52575, 94.59737, 
    94.88748, 95.53965, 95.32225, 95.87054, 95.85813, 96.47083, 96.19428, 
    97.22755, 96.93317, 97.78524, 97.57054, 97.77516, 97.71307, 97.77597, 
    97.46121, 97.596, 97.31927, 96.24606, 96.56075, 95.62409, 95.05607, 
    94.67305, 94.40189, 94.44019, 94.51326, 94.88918, 95.24337, 95.50746, 
    95.68311, 95.85635, 96.38218, 96.66099, 97.28719, 97.17392, 97.3658, 
    97.54919, 97.85769, 97.80686, 97.94294, 97.36067, 97.74744, 97.10945, 
    97.28371, 95.90381, 95.38085, 95.15476, 94.95482, 94.46966, 94.80456, 
    94.67246, 94.98685, 95.18698, 95.08795, 95.68791, 95.45699, 96.67753, 
    96.15063, 97.52779, 97.19716, 97.60713, 97.39779, 97.75668, 97.43364, 
    97.99358, 98.11581, 98.03228, 98.35325, 97.41576, 97.77519, 95.08519, 
    95.10134, 95.17656, 94.84619, 94.82599, 94.5238, 94.79263, 94.90728, 
    95.19856, 95.36915, 95.52836, 95.87897, 96.27151, 96.82198, 97.21857, 
    97.48498, 97.32155, 97.46583, 97.30456, 97.22901, 98.07002, 97.59727, 
    98.30704, 98.26768, 97.94619, 98.27211, 95.11267, 95.01978, 94.69775, 
    94.94971, 94.49092, 94.7476, 94.8954, 95.46188, 95.58378, 95.69699, 
    95.92075, 96.20843, 96.71437, 97.15584, 97.55986, 97.53022, 97.54066, 
    97.63107, 97.40724, 97.66785, 97.71165, 97.59718, 98.26241, 98.07207, 
    98.26685, 98.14288, 95.04996, 95.20632, 95.12182, 95.28078, 95.16879, 
    95.65636, 95.80157, 96.48279, 96.20277, 96.64856, 96.24798, 96.3189, 
    96.66326, 96.26958, 97.13152, 96.54677, 97.63459, 97.04894, 97.67136, 
    97.55811, 97.74564, 97.9138, 98.12555, 98.51707, 98.42632, 98.75422, 
    95.43557, 95.63271, 95.61529, 95.8218, 95.97472, 96.30659, 96.84041, 
    96.63944, 97.00851, 97.08273, 96.52206, 96.86613, 95.76475, 95.94223, 
    95.83649, 95.45115, 96.68581, 96.051, 97.22514, 96.87976, 97.88982, 
    97.38677, 98.37639, 98.80143, 99.20216, 99.67202, 95.74035, 95.60628, 
    95.84636, 96.17924, 96.48856, 96.90082, 96.94302, 97.02042, 97.22097, 
    97.38982, 97.04495, 97.43217, 95.98354, 96.741, 95.55568, 95.91175, 
    96.15958, 96.05075, 96.61647, 96.75012, 97.2944, 97.01278, 98.69648, 
    97.94943, 100.0304, 99.44633, 95.55948, 95.73985, 96.36935, 96.06951, 
    96.92834, 97.14048, 97.31309, 97.5341, 97.55794, 97.68904, 97.47427, 
    97.68053, 96.9017, 97.24927, 96.2972, 96.52843, 96.42199, 96.30537, 
    96.6656, 97.05039, 97.05852, 97.18212, 97.53111, 96.93183, 98.79333, 
    97.64138, 95.93679, 96.28539, 96.33512, 96.19997, 97.1192, 96.78554, 
    97.68583, 97.44199, 97.84167, 97.64295, 97.61374, 97.35889, 97.20045, 
    96.80083, 96.4764, 96.21956, 96.27924, 96.5615, 97.07394, 97.56014, 
    97.45352, 97.81126, 96.86592, 97.2617, 97.10864, 97.50801, 96.63412, 
    97.37829, 96.4445, 96.52614, 96.77892, 97.28864, 97.40149, 97.52224, 
    97.4477, 97.08694, 97.02788, 96.77274, 96.70242, 96.50835, 96.3479, 
    96.49451, 96.64865, 97.08705, 97.48322, 97.91621, 98.02231, 98.53026, 
    98.11678, 98.79979, 98.21914, 99.22546, 97.42137, 98.20189, 96.7904, 
    96.94184, 97.21624, 97.84715, 97.50613, 97.90496, 97.02555, 96.5713, 
    96.45386, 96.23518, 96.45886, 96.44065, 96.65497, 96.58606, 97.10163, 
    96.82448, 97.61304, 97.90179, 98.71986, 99.22343, 99.73743, 99.9649, 
    100.0342, 100.0632,
  129.9302, 130.6424, 130.5037, 131.0702, 130.7599, 131.1261, 130.0743, 
    130.6708, 130.2898, 129.9941, 132.1563, 131.0951, 133.2638, 132.5828, 
    134.2974, 133.1577, 134.5279, 134.2643, 135.0584, 134.8306, 135.8499, 
    135.1637, 136.3799, 135.6857, 135.7942, 135.1411, 131.3081, 132.0239, 
    131.2658, 131.3677, 131.3219, 130.7666, 130.4784, 129.8758, 129.985, 
    130.4277, 131.4135, 131.0822, 131.918, 131.899, 132.8335, 132.4116, 
    133.9884, 133.539, 134.8401, 134.5122, 134.8247, 134.7299, 134.826, 
    134.3452, 134.551, 134.1284, 132.4906, 132.9707, 131.5422, 130.6849, 
    130.1005, 129.6868, 129.7453, 129.8567, 130.4303, 130.9649, 131.3645, 
    131.6322, 131.8963, 132.6982, 133.1236, 134.0794, 133.9065, 134.1995, 
    134.4796, 134.9508, 134.8732, 135.0811, 134.1917, 134.7824, 133.8081, 
    134.0741, 131.9686, 131.1715, 130.834, 130.5304, 129.7902, 130.3011, 
    130.0996, 130.5793, 130.8816, 130.7336, 131.6395, 131.2876, 133.1488, 
    132.3451, 134.4469, 133.942, 134.5681, 134.2483, 134.7965, 134.3031, 
    135.1584, 135.3452, 135.2176, 135.7081, 134.2758, 134.8248, 130.7294, 
    130.754, 130.8662, 130.3647, 130.3338, 129.8728, 130.2829, 130.4579, 
    130.8987, 131.1537, 131.3963, 131.9308, 132.5294, 133.3693, 133.9747, 
    134.3815, 134.1319, 134.3522, 134.106, 133.9906, 135.2752, 134.553, 
    135.6375, 135.5773, 135.086, 135.5841, 130.7713, 130.6295, 130.1382, 
    130.5226, 129.8226, 130.2142, 130.4397, 131.295, 131.4808, 131.6534, 
    131.9945, 132.4332, 133.2051, 133.8789, 134.4958, 134.4506, 134.4665, 
    134.6046, 134.2628, 134.6608, 134.7277, 134.5529, 135.5693, 135.2784, 
    135.576, 135.3866, 130.6756, 130.9102, 130.7853, 131.0202, 130.8548, 
    131.5914, 131.8128, 132.8517, 132.4246, 133.1046, 132.4935, 132.6017, 
    133.1271, 132.5265, 133.8418, 132.9493, 134.61, 133.7157, 134.6662, 
    134.4932, 134.7796, 135.0365, 135.3601, 135.9586, 135.8198, 136.3212, 
    131.2549, 131.5554, 131.5288, 131.8436, 132.0768, 132.5829, 133.3974, 
    133.0907, 133.654, 133.7673, 132.9116, 133.4367, 131.7567, 132.0273, 
    131.866, 131.2786, 133.1615, 132.1931, 133.9847, 133.4575, 134.9999, 
    134.2315, 135.7435, 136.3933, 137.0063, 137.7253, 131.7195, 131.5151, 
    131.8811, 132.3887, 132.8605, 133.4896, 133.554, 133.6722, 133.9783, 
    134.2362, 133.7096, 134.3008, 132.0902, 133.2457, 131.438, 131.9808, 
    132.3587, 132.1927, 133.0557, 133.2596, 134.0905, 133.6605, 136.2328, 
    135.091, 138.274, 137.3799, 131.4438, 131.7187, 132.6787, 132.2213, 
    133.5316, 133.8555, 134.119, 134.4565, 134.4929, 134.6932, 134.3651, 
    134.6802, 133.491, 134.0215, 132.5686, 132.9214, 132.759, 132.5811, 
    133.1307, 133.7179, 133.7303, 133.919, 134.4519, 133.537, 136.3809, 
    134.6203, 132.019, 132.5506, 132.6265, 132.4203, 133.823, 133.3137, 
    134.6882, 134.3158, 134.9263, 134.6228, 134.5781, 134.1889, 133.947, 
    133.337, 132.842, 132.4502, 132.5412, 132.9718, 133.7538, 134.4963, 
    134.3334, 134.8799, 133.4364, 134.0405, 133.8068, 134.4167, 133.0826, 
    134.2185, 132.7933, 132.9179, 133.3036, 134.0816, 134.254, 134.4384, 
    134.3246, 133.7737, 133.6835, 133.2942, 133.1868, 132.8907, 132.646, 
    132.8696, 133.1048, 133.7739, 134.3788, 135.0402, 135.2023, 135.9787, 
    135.3467, 136.3908, 135.5031, 137.0419, 134.2843, 135.4767, 133.3211, 
    133.5522, 133.9711, 134.9347, 134.4138, 135.023, 133.68, 132.9868, 
    132.8076, 132.474, 132.8152, 132.7874, 133.1144, 133.0093, 133.7961, 
    133.3731, 134.5771, 135.0182, 136.2686, 137.0388, 137.8254, 138.1737, 
    138.2798, 138.3241,
  195.7734, 196.8862, 196.6695, 197.5698, 197.0699, 197.66, 195.9986, 
    196.9306, 196.3352, 195.8733, 199.3256, 197.61, 201.1182, 200.0159, 
    202.7931, 200.9465, 203.1668, 202.7394, 204.0273, 203.6577, 205.281, 
    204.198, 206.1129, 205.0235, 205.1937, 204.1614, 197.9542, 199.1115, 
    197.8858, 198.0505, 197.9766, 197.0803, 196.6299, 195.6884, 195.8591, 
    196.5506, 198.1246, 197.5892, 198.9402, 198.9096, 200.4215, 199.7388, 
    202.2922, 201.5641, 203.6732, 203.1413, 203.6482, 203.4944, 203.6502, 
    202.8706, 203.2043, 202.5192, 199.8666, 200.6436, 198.3327, 196.9526, 
    196.0394, 195.3933, 195.4846, 195.6586, 196.5546, 197.3996, 198.0453, 
    198.4781, 198.9052, 200.2025, 200.8912, 202.4398, 202.1595, 202.6343, 
    203.0884, 203.8527, 203.7267, 204.064, 202.6217, 203.5795, 202.0001, 
    202.4312, 199.0221, 197.7335, 197.1881, 196.7112, 195.5548, 196.3529, 
    196.038, 196.7876, 197.265, 197.0288, 198.49, 197.921, 200.9321, 
    199.6311, 203.0354, 202.217, 203.2319, 202.7136, 203.6024, 202.8023, 
    204.1896, 204.4894, 204.2855, 205.0586, 202.758, 203.6483, 197.0222, 
    197.0607, 197.2402, 196.4521, 196.404, 195.6837, 196.3244, 196.5978, 
    197.2927, 197.7047, 198.0968, 198.961, 199.9294, 201.2891, 202.27, 
    202.9294, 202.5249, 202.882, 202.4828, 202.2959, 204.3791, 203.2075, 
    204.9478, 204.8534, 204.0721, 204.8641, 197.0877, 196.8661, 196.0983, 
    196.699, 195.6054, 196.2171, 196.5695, 197.933, 198.2334, 198.5123, 
    199.064, 199.7737, 201.0232, 202.1148, 203.1149, 203.0414, 203.0673, 
    203.2912, 202.737, 203.3823, 203.4908, 203.2073, 204.8408, 204.3842, 
    204.8514, 204.5543, 196.9381, 197.3112, 197.1095, 197.4889, 197.2216, 
    198.4122, 198.7701, 200.451, 199.7598, 200.8606, 199.8714, 200.0464, 
    200.8968, 199.9247, 202.0546, 200.609, 203.2999, 201.8503, 203.391, 
    203.1105, 203.575, 203.9918, 204.5127, 205.4515, 205.2338, 206.0206, 
    197.8682, 198.3539, 198.311, 198.82, 199.1971, 200.0161, 201.3347, 
    200.8381, 201.7504, 201.9339, 200.5481, 201.3983, 198.6794, 199.117, 
    198.8562, 197.9066, 200.9526, 199.3853, 202.2863, 201.432, 203.9323, 
    202.6862, 205.1141, 206.1339, 207.0966, 208.2265, 198.6192, 198.2888, 
    198.8806, 199.7017, 200.4653, 201.4841, 201.5884, 201.7798, 202.276, 
    202.6938, 201.8405, 202.7987, 199.2188, 201.089, 198.1641, 199.0418, 
    199.6532, 199.3847, 200.7813, 201.1116, 202.4576, 201.7609, 205.882, 
    204.08, 209.0895, 207.6836, 198.1735, 198.618, 200.1709, 199.431, 
    201.5521, 202.0768, 202.5039, 203.051, 203.1101, 203.4348, 202.9029, 
    203.4137, 201.4862, 202.346, 199.9929, 200.5638, 200.301, 200.013, 
    200.9027, 201.8539, 201.8741, 202.1798, 203.0434, 201.5608, 206.1144, 
    203.3166, 199.1036, 199.9637, 200.0865, 199.7529, 202.0242, 201.1991, 
    203.4268, 202.823, 203.813, 203.3206, 203.2483, 202.6173, 202.2252, 
    201.2369, 200.4353, 199.8012, 199.9485, 200.6455, 201.9121, 203.1155, 
    202.8515, 203.7377, 201.3978, 202.3767, 201.998, 202.9865, 200.8249, 
    202.6651, 200.3566, 200.5582, 201.1827, 202.4433, 202.7227, 203.0217, 
    202.8371, 201.9443, 201.7982, 201.1675, 200.9937, 200.5143, 200.1181, 
    200.4801, 200.8608, 201.9446, 202.925, 203.9977, 204.2608, 205.4831, 
    204.4917, 206.1299, 204.7369, 207.1525, 202.7718, 204.6956, 201.2111, 
    201.5855, 202.2642, 203.8265, 202.9818, 203.9698, 201.7925, 200.6697, 
    200.3797, 199.8398, 200.392, 200.3471, 200.8765, 200.7062, 201.9807, 
    201.2954, 203.2465, 203.962, 205.9382, 207.1477, 208.384, 208.9317, 
    209.0986, 209.1684,
  319.7102, 321.5075, 321.1573, 322.6125, 321.8044, 322.7585, 320.0737, 
    321.5792, 320.6173, 319.8715, 325.4546, 322.6776, 328.3621, 326.5736, 
    331.0837, 328.0833, 331.6917, 330.9965, 333.0863, 332.4908, 335.1092, 
    333.355, 336.4668, 334.6893, 334.9669, 333.2973, 323.2344, 325.1077, 
    323.1238, 323.3902, 323.2706, 321.8212, 321.0933, 319.5731, 319.8485, 
    320.9652, 323.5101, 322.6439, 324.8305, 324.781, 327.2316, 326.1245, 
    330.2693, 329.0862, 332.5159, 331.6502, 332.4753, 332.2249, 332.4785, 
    331.2097, 331.7528, 330.6384, 326.3316, 327.5919, 323.8468, 321.6148, 
    320.1396, 319.0969, 319.2441, 319.525, 320.9718, 322.3374, 323.3819, 
    324.0823, 324.7739, 326.8762, 327.9937, 330.5092, 330.0536, 330.8255, 
    331.5642, 332.8083, 332.6031, 333.144, 330.805, 332.3634, 329.7945, 
    330.4953, 324.9629, 322.8773, 321.9954, 321.2246, 319.3574, 320.6458, 
    320.1374, 321.3481, 322.1198, 321.7379, 324.1015, 323.1807, 328.06, 
    325.9498, 331.478, 330.1471, 331.7977, 330.9544, 332.4007, 331.0988, 
    333.3417, 333.8188, 333.4927, 334.7467, 331.0268, 332.4753, 321.7273, 
    321.7895, 322.0797, 320.8062, 320.7284, 319.5656, 320.6, 321.0415, 
    322.1646, 322.8307, 323.4651, 324.8641, 326.4334, 328.6396, 330.2332, 
    331.3055, 330.6476, 331.2284, 330.5792, 330.2753, 333.64, 331.7579, 
    334.5661, 334.4122, 333.1567, 334.4295, 321.8332, 321.4751, 320.2347, 
    321.205, 319.4391, 320.4266, 320.9957, 323.2001, 323.6861, 324.1377, 
    325.0311, 326.1811, 328.2079, 329.9809, 331.6072, 331.4878, 331.5298, 
    331.8942, 330.9925, 332.0424, 332.2191, 331.7576, 334.3916, 333.6481, 
    334.4089, 333.9246, 321.5914, 322.1945, 321.8685, 322.4818, 322.0497, 
    323.9755, 324.555, 327.2794, 326.1584, 327.9439, 326.3393, 326.6232, 
    328.0026, 326.4258, 329.883, 327.5357, 331.9084, 329.551, 332.0566, 
    331.6002, 332.3562, 333.0304, 333.8569, 335.3875, 335.0324, 336.3163, 
    323.0953, 323.8812, 323.8118, 324.6359, 325.2466, 326.5739, 328.7137, 
    327.9074, 329.3888, 329.687, 327.4369, 328.8169, 324.4081, 325.1167, 
    324.6945, 323.1573, 328.0933, 325.5514, 330.2596, 328.8717, 332.9368, 
    330.9099, 334.8372, 336.5012, 338.074, 339.9221, 324.3107, 323.7759, 
    324.734, 326.0642, 327.3026, 328.9562, 329.1257, 329.4366, 330.2429, 
    330.9223, 329.5351, 331.0929, 325.2816, 328.3147, 323.574, 324.9949, 
    325.9856, 325.5505, 327.8154, 328.3514, 330.5382, 329.4059, 336.0898, 
    333.1692, 341.3355, 339.0337, 323.5893, 324.3088, 326.8251, 325.6255, 
    329.0668, 329.9192, 330.6135, 331.5034, 331.5995, 332.1279, 331.2624, 
    332.0936, 328.9597, 330.3567, 326.5363, 327.4624, 327.036, 326.5691, 
    328.0124, 329.5569, 329.5898, 330.0866, 331.4908, 329.0808, 336.4691, 
    331.9353, 325.0952, 326.4889, 326.6881, 326.1473, 329.8336, 328.4934, 
    332.115, 331.1324, 332.7437, 331.9421, 331.8243, 330.7978, 330.1603, 
    328.5548, 327.2539, 326.2257, 326.4645, 327.5949, 329.6516, 331.6083, 
    331.1787, 332.6209, 328.8161, 330.4066, 329.7911, 331.3983, 327.8861, 
    330.8754, 327.1262, 327.4532, 328.4669, 330.515, 330.9693, 331.4556, 
    331.1554, 329.7039, 329.4666, 328.4422, 328.16, 327.382, 326.7393, 
    327.3265, 327.9443, 329.7044, 331.2984, 333.0397, 333.4538, 335.4389, 
    333.8224, 336.4944, 334.2219, 338.1651, 331.0491, 334.1548, 328.513, 
    329.121, 330.2237, 332.7655, 331.3907, 332.9958, 329.4572, 327.6341, 
    327.1637, 326.2881, 327.1837, 327.1108, 327.9697, 327.6935, 329.763, 
    328.6498, 331.8214, 332.9834, 336.1816, 338.1574, 340.18, 341.0769, 
    341.3503, 341.4647,
  524.6362, 527.9112, 527.2731, 529.9263, 528.4524, 530.1926, 525.3007, 
    528.0417, 526.2898, 524.9329, 535.1221, 530.045, 540.4579, 537.1735, 
    545.4712, 539.9454, 546.5938, 545.3104, 549.1837, 548.0705, 553.063, 
    549.6983, 555.673, 552.257, 552.7897, 549.5878, 531.0616, 534.4869, 
    530.8596, 531.3462, 531.1277, 528.4829, 527.1564, 524.3782, 524.8911, 
    526.9232, 531.5651, 529.9836, 533.9798, 533.8891, 538.3809, 536.3499, 
    543.9693, 541.7901, 548.1169, 546.5172, 548.0417, 547.5788, 548.0477, 
    545.7039, 546.7066, 544.6497, 536.7297, 539.0425, 532.1805, 528.1065, 
    525.4206, 523.4825, 523.7594, 524.2877, 526.9351, 529.4243, 531.331, 
    532.6111, 533.8761, 537.7286, 539.7807, 544.4114, 543.5718, 544.9949, 
    546.3583, 548.6575, 548.2782, 549.2941, 544.9571, 547.8348, 543.0943, 
    544.3858, 534.2219, 530.4097, 528.8004, 527.3958, 523.9724, 526.3417, 
    525.4164, 527.6207, 529.0274, 528.3311, 532.6462, 530.9636, 539.9026, 
    536.0297, 546.1991, 543.744, 546.7896, 545.2328, 547.9037, 545.4991, 
    549.6728, 550.587, 549.9621, 552.3671, 545.3663, 548.0418, 528.3116, 
    528.4252, 528.9542, 526.6336, 526.492, 524.364, 526.2582, 527.0621, 
    529.109, 530.3245, 531.4831, 534.0413, 536.9163, 540.9684, 543.9027, 
    545.8807, 544.6667, 545.7384, 544.5406, 543.9802, 550.2443, 546.7161, 
    552.0204, 551.7252, 549.3184, 551.7584, 528.5048, 527.8521, 525.5936, 
    527.36, 524.1262, 525.9426, 526.9787, 530.9989, 531.8869, 532.7123, 
    534.3468, 536.4537, 540.1744, 543.4376, 546.4377, 546.2172, 546.2949, 
    546.9678, 545.303, 547.2417, 547.5681, 546.7155, 551.6857, 550.2599, 
    551.7189, 550.79, 528.0641, 529.1636, 528.5692, 529.6877, 528.8994, 
    532.4156, 533.4754, 538.4686, 536.4122, 539.6893, 536.7438, 537.2643, 
    539.7971, 536.9024, 543.2573, 538.9393, 546.994, 542.6456, 547.2679, 
    546.4247, 547.8215, 549.0765, 550.6602, 553.5977, 552.9157, 555.3835, 
    530.8077, 532.2434, 532.1166, 533.6236, 534.7415, 537.1741, 541.1046, 
    539.6224, 542.3472, 542.8963, 538.7581, 541.2944, 533.2067, 534.5035, 
    533.7308, 530.9209, 539.9638, 535.2996, 543.9514, 541.3953, 548.8974, 
    545.1506, 552.5407, 555.739, 558.7693, 562.2427, 533.0287, 532.0509, 
    533.803, 536.2394, 538.5114, 541.5508, 541.8629, 542.4351, 543.9206, 
    545.1736, 542.6165, 545.4882, 534.8053, 540.3709, 531.682, 534.2806, 
    536.0953, 535.298, 539.4532, 540.4384, 544.465, 542.3787, 554.9477, 
    549.3423, 564.8874, 560.5832, 531.7098, 533.0253, 537.6348, 535.4355, 
    541.7543, 543.324, 544.6039, 546.2459, 546.4234, 547.3995, 545.8011, 
    547.3362, 541.5573, 544.1303, 537.1052, 538.8048, 538.022, 537.1652, 
    539.8152, 542.6566, 542.7172, 543.6324, 546.2225, 541.7802, 555.6771, 
    547.0435, 534.4642, 537.0181, 537.3836, 536.3918, 543.1664, 540.6996, 
    547.3757, 545.5612, 548.538, 547.0563, 546.8387, 544.9438, 543.7684, 
    540.8124, 538.4219, 536.5354, 536.9733, 539.0482, 542.8309, 546.4396, 
    545.6467, 548.3111, 541.2931, 544.2224, 543.088, 546.0519, 539.5831, 
    545.0868, 538.1875, 538.788, 540.6508, 544.4221, 545.2603, 546.1577, 
    545.6036, 542.9274, 542.4903, 540.6053, 540.0865, 538.6572, 537.4776, 
    538.5553, 539.6901, 542.9283, 545.8675, 549.0944, 549.8876, 553.6963, 
    550.5939, 555.7258, 551.3597, 558.9449, 545.4073, 551.2312, 540.7356, 
    541.8542, 543.8851, 548.5783, 546.038, 549.0102, 542.4731, 539.1201, 
    538.2563, 536.65, 538.2931, 538.1592, 539.7369, 539.2292, 543.0363, 
    540.9871, 546.8334, 548.9865, 555.1243, 558.9301, 562.7249, 564.4031, 
    564.9152, 565.1295,
  947.2838, 954.1564, 952.8134, 958.4071, 955.2968, 958.97, 948.6698, 
    954.4313, 950.7461, 947.8985, 969.2881, 958.6579, 980.3278, 973.5209, 
    990.7889, 979.2632, 993.1436, 990.4521, 998.5929, 996.2478, 1006.801, 
    999.6788, 1012.354, 1005.091, 1006.221, 999.4456, 960.808, 967.9803, 
    960.3805, 961.4104, 960.9479, 955.3611, 952.5677, 946.7616, 947.811, 
    952.0774, 961.8741, 958.5283, 966.9371, 966.7508, 976.019, 971.8199, 
    987.6457, 983.0991, 996.3455, 992.9828, 996.1871, 995.2134, 996.1998, 
    991.2768, 993.3805, 989.0688, 972.604, 977.39, 963.1784, 954.5679, 
    948.9214, 944.9503, 945.5099, 946.5786, 952.1024, 957.347, 961.3782, 
    964.0917, 966.724, 974.6688, 978.9212, 988.5703, 986.8151, 989.7913, 
    992.6494, 997.4839, 996.685, 998.826, 989.7121, 995.7519, 985.8182, 
    988.5167, 967.4349, 959.4288, 956.0305, 953.0714, 945.9407, 950.8552, 
    948.9126, 953.545, 956.5095, 955.0411, 964.1661, 960.6005, 979.1743, 
    971.1592, 992.3152, 987.1749, 993.5547, 990.2895, 995.897, 990.8476, 
    999.6248, 1001.556, 1000.236, 1005.325, 990.5692, 996.1874, 955.0002, 
    955.2394, 956.3549, 951.4685, 951.1709, 946.733, 950.6798, 952.3695, 
    956.6816, 959.2488, 961.7003, 967.0635, 972.9896, 981.3889, 987.5066, 
    991.6475, 989.1043, 991.349, 988.8405, 987.6686, 1000.832, 993.4003, 
    1004.59, 1003.964, 998.8771, 1004.035, 955.4073, 954.032, 949.2843, 
    952.9962, 946.2518, 950.017, 952.194, 960.6752, 962.5559, 964.3064, 
    967.6921, 972.0341, 979.7388, 986.535, 992.816, 992.3533, 992.5162, 
    993.9291, 990.4365, 994.5046, 995.1907, 993.3991, 1003.88, 1000.865, 
    1003.951, 1001.985, 954.4786, 956.7967, 955.5429, 957.9031, 956.2394, 
    963.6769, 965.9005, 976.2006, 971.9484, 978.7314, 972.6332, 973.7089, 
    978.9553, 972.9609, 986.1584, 977.1758, 993.9841, 984.882, 994.5598, 
    992.7888, 995.7239, 998.367, 1001.71, 1007.937, 1006.488, 1011.737, 
    960.2706, 963.3117, 963.0428, 966.205, 968.5043, 973.5223, 981.6723, 
    978.5926, 984.2598, 985.405, 976.8002, 982.0672, 965.3486, 968.0146, 
    966.4254, 960.5102, 979.3013, 969.6539, 987.6084, 982.2771, 997.9894, 
    990.1174, 1005.693, 1012.495, 1018.976, 1026.654, 964.9781, 962.9036, 
    966.5739, 971.5917, 976.2893, 982.6008, 983.2506, 984.4431, 987.5439, 
    990.1655, 984.8212, 990.8246, 968.6357, 980.1469, 962.1218, 967.5558, 
    971.2944, 969.6506, 978.2416, 980.2872, 988.6823, 984.3255, 1010.809, 
    998.9277, 1032.464, 1022.954, 962.1808, 964.9707, 974.4749, 969.9338, 
    983.0247, 986.2976, 988.973, 992.4135, 992.7859, 994.8365, 991.4805, 
    994.7033, 982.6144, 987.9824, 973.3798, 976.8972, 975.276, 973.5038, 
    978.9928, 984.905, 985.0313, 986.9418, 992.3644, 983.0783, 1012.363, 
    994.088, 967.9335, 973.1997, 973.9553, 971.9063, 985.9686, 980.83, 
    994.7863, 990.9777, 997.2322, 994.1151, 993.658, 989.6844, 987.2258, 
    981.0646, 976.104, 972.2029, 973.1074, 977.4016, 985.2687, 992.82, 
    991.1567, 996.7543, 982.0645, 988.1749, 985.8051, 992.0066, 978.5112, 
    989.9837, 975.6186, 976.8624, 980.7285, 988.5925, 990.347, 992.2284, 
    991.0665, 985.4697, 984.5581, 980.634, 979.556, 976.5913, 974.1497, 
    976.3802, 978.7331, 985.4718, 991.6196, 998.4048, 1000.078, 1008.146, 
    1001.57, 1012.467, 1003.19, 1019.352, 990.6551, 1002.918, 980.9048, 
    983.2325, 987.4698, 997.3171, 991.9772, 998.2272, 984.5223, 977.5508, 
    975.761, 972.4394, 975.8372, 975.5599, 978.8302, 977.777, 985.697, 
    981.4279, 993.6467, 998.1773, 1011.185, 1019.321, 1027.731, 1031.413, 
    1032.524, 1032.99,
  1829.892, 1849.354, 1845.526, 1861.551, 1852.614, 1863.175, 1833.792, 
    1850.139, 1839.658, 1831.62, 1893.773, 1862.274, 1928.095, 1906.815, 
    1960.692, 1924.742, 1968.122, 1959.633, 1985.508, 1977.993, 2012.213, 
    1989.004, 2030.649, 2006.597, 2010.305, 1988.253, 1868.495, 1889.772, 
    1867.256, 1870.244, 1868.901, 1852.798, 1844.827, 1828.426, 1831.374, 
    1843.433, 1871.592, 1861.9, 1886.59, 1886.023, 1914.58, 1901.557, 
    1950.849, 1936.76, 1978.305, 1967.613, 1977.799, 1974.694, 1977.84, 
    1962.227, 1968.872, 1955.294, 1903.978, 1918.864, 1875.391, 1850.529, 
    1834.501, 1823.355, 1824.92, 1827.913, 1843.505, 1858.498, 1870.151, 
    1878.059, 1885.941, 1910.377, 1923.666, 1953.735, 1948.262, 1957.558, 
    1966.559, 1981.948, 1979.39, 1986.257, 1957.31, 1976.41, 1945.165, 
    1953.568, 1888.107, 1864.501, 1854.716, 1846.261, 1826.125, 1839.966, 
    1834.476, 1847.61, 1856.09, 1851.883, 1878.276, 1867.893, 1924.462, 
    1899.52, 1965.503, 1949.381, 1969.424, 1959.122, 1976.873, 1960.876, 
    1988.83, 1995.075, 1990.802, 2007.362, 1960.001, 1977.8, 1851.765, 
    1852.45, 1855.647, 1841.705, 1840.861, 1828.346, 1839.47, 1844.264, 
    1856.585, 1863.981, 1871.086, 1886.975, 1905.17, 1931.448, 1950.415, 
    1963.396, 1955.406, 1962.455, 1954.58, 1950.92, 1992.729, 1968.935, 
    2004.955, 2002.911, 1986.422, 2003.141, 1852.931, 1848.999, 1835.525, 
    1846.047, 1826.997, 1837.595, 1843.765, 1868.11, 1873.576, 1878.687, 
    1888.892, 1902.217, 1926.239, 1947.39, 1967.086, 1965.623, 1966.137, 
    1970.612, 1959.584, 1972.439, 1974.622, 1968.931, 2002.638, 1992.836, 
    2002.868, 1996.467, 1850.274, 1856.915, 1853.319, 1860.098, 1855.316, 
    1876.847, 1883.437, 1915.147, 1901.953, 1923.07, 1904.068, 1907.397, 
    1923.773, 1905.081, 1946.221, 1918.194, 1970.786, 1942.264, 1972.615, 
    1966.999, 1976.321, 1984.782, 1995.576, 2015.958, 2011.184, 2028.585, 
    1866.937, 1875.78, 1874.995, 1884.362, 1891.373, 1906.819, 1932.345, 
    1922.634, 1940.34, 1943.883, 1917.019, 1933.587, 1881.762, 1889.876, 
    1885.032, 1867.631, 1924.862, 1894.894, 1950.732, 1934.232, 1983.569, 
    1958.582, 2008.57, 2031.12, 2053.035, 2079.241, 1880.653, 1874.59, 
    1885.484, 1900.853, 1915.424, 1935.227, 1937.227, 1940.906, 1950.531, 
    1958.733, 1942.076, 1960.804, 1891.775, 1927.525, 1872.312, 1888.476, 
    1899.937, 1894.884, 1921.533, 1927.967, 1954.085, 1940.543, 2025.486, 
    1986.585, 2099.51, 2066.706, 1872.484, 1880.632, 1909.774, 1895.753, 
    1936.531, 1946.653, 1954.994, 1965.813, 1966.99, 1973.494, 1962.869, 
    1973.071, 1935.268, 1951.899, 1906.378, 1917.322, 1912.265, 1906.762, 
    1923.891, 1942.335, 1942.726, 1948.656, 1965.658, 1936.696, 2030.678, 
    1971.116, 1889.629, 1905.82, 1908.162, 1901.823, 1945.631, 1929.681, 
    1973.335, 1961.286, 1981.141, 1971.202, 1969.752, 1957.223, 1949.54, 
    1930.422, 1914.845, 1902.738, 1905.534, 1918.9, 1943.461, 1967.098, 
    1961.849, 1979.612, 1933.578, 1952.5, 1945.124, 1964.528, 1922.379, 
    1958.162, 1913.332, 1917.214, 1929.36, 1953.804, 1959.303, 1965.228, 
    1961.565, 1944.084, 1941.262, 1929.062, 1925.663, 1916.366, 1908.765, 
    1915.707, 1923.075, 1944.09, 1963.308, 1984.903, 1990.294, 2016.65, 
    1995.122, 2031.026, 2000.387, 2054.322, 1960.271, 1999.501, 1929.917, 
    1937.171, 1950.3, 1981.413, 1964.435, 1984.333, 1941.151, 1919.367, 
    1913.776, 1903.469, 1914.013, 1913.15, 1923.38, 1920.076, 1944.789, 
    1931.571, 1969.716, 1984.172, 2026.741, 2054.214, 2082.901, 2095.762, 
    2099.725, 2101.389,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.482451, 4.50081, 4.497236, 4.512078, 4.50384, 4.513565, 4.486168, 
    4.50154, 4.491722, 4.484101, 4.540988, 4.512741, 4.570472, 4.552351, 
    4.597974, 4.567649, 4.604106, 4.597096, 4.618218, 4.61216, 4.639256, 
    4.621017, 4.653348, 4.634895, 4.637779, 4.620416, 4.518414, 4.537464, 
    4.517287, 4.52, 4.518782, 4.50401, 4.49658, 4.48105, 4.483866, 4.495274, 
    4.52122, 4.512399, 4.534654, 4.53415, 4.559023, 4.547795, 4.589756, 
    4.5778, 4.612413, 4.60369, 4.612003, 4.609481, 4.612036, 4.599247, 
    4.604723, 4.593482, 4.549897, 4.562674, 4.524648, 4.501902, 4.486841, 
    4.476179, 4.477685, 4.480557, 4.495341, 4.509275, 4.519916, 4.527045, 
    4.534078, 4.555418, 4.566742, 4.592177, 4.587578, 4.59537, 4.602823, 
    4.615355, 4.613291, 4.618819, 4.595164, 4.610875, 4.58496, 4.592038, 
    4.535993, 4.514777, 4.505785, 4.497923, 4.478843, 4.492013, 4.486818, 
    4.499184, 4.507056, 4.503161, 4.52724, 4.517867, 4.567414, 4.546021, 
    4.601953, 4.588522, 4.605176, 4.596673, 4.611251, 4.598129, 4.620878, 
    4.625842, 4.622449, 4.635493, 4.597402, 4.612003, 4.503053, 4.503687, 
    4.506647, 4.49365, 4.492856, 4.480973, 4.491545, 4.496053, 4.507513, 
    4.514302, 4.520763, 4.534994, 4.550929, 4.573282, 4.589392, 4.600214, 
    4.593575, 4.599436, 4.592885, 4.589817, 4.623981, 4.604774, 4.633615, 
    4.632016, 4.618951, 4.632196, 4.504134, 4.50048, 4.487813, 4.497724, 
    4.47968, 4.489773, 4.495585, 4.518063, 4.523013, 4.527607, 4.536691, 
    4.548369, 4.568912, 4.586842, 4.603256, 4.602052, 4.602476, 4.606149, 
    4.597056, 4.607643, 4.609422, 4.604772, 4.631802, 4.624067, 4.631982, 
    4.626945, 4.501667, 4.507817, 4.504493, 4.510746, 4.506341, 4.525956, 
    4.531849, 4.559506, 4.54814, 4.566239, 4.549975, 4.552854, 4.566831, 
    4.550853, 4.585853, 4.562102, 4.606292, 4.582496, 4.607786, 4.603185, 
    4.610804, 4.617635, 4.62624, 4.642148, 4.638461, 4.651788, 4.516998, 
    4.524998, 4.524292, 4.532674, 4.538881, 4.552356, 4.574031, 4.565871, 
    4.58086, 4.583874, 4.561105, 4.575075, 4.530357, 4.53756, 4.53327, 
    4.517629, 4.567751, 4.541975, 4.589658, 4.57563, 4.616661, 4.596221, 
    4.636432, 4.653702, 4.669997, 4.689095, 4.529367, 4.523927, 4.533672, 
    4.547182, 4.559743, 4.576485, 4.5782, 4.581343, 4.58949, 4.596349, 
    4.582337, 4.598069, 4.539232, 4.569993, 4.521872, 4.536322, 4.546384, 
    4.541968, 4.564939, 4.570366, 4.59247, 4.581034, 4.649436, 4.61908, 
    4.703672, 4.67992, 4.522027, 4.529349, 4.554902, 4.54273, 4.577604, 
    4.586219, 4.593232, 4.602208, 4.603178, 4.608503, 4.599779, 4.608158, 
    4.576521, 4.590639, 4.551975, 4.561363, 4.557042, 4.552306, 4.566934, 
    4.582558, 4.582891, 4.58791, 4.602076, 4.577746, 4.653366, 4.606557, 
    4.537343, 4.551491, 4.553514, 4.548028, 4.585355, 4.571804, 4.608373, 
    4.598468, 4.614706, 4.606632, 4.605445, 4.595092, 4.588655, 4.572424, 
    4.559249, 4.548823, 4.551246, 4.562705, 4.583514, 4.603266, 4.598934, 
    4.613471, 4.575068, 4.591142, 4.584925, 4.60115, 4.565655, 4.595869, 
    4.557956, 4.561271, 4.571535, 4.592234, 4.596823, 4.601727, 4.5987, 
    4.584044, 4.581645, 4.571285, 4.568428, 4.560549, 4.554034, 4.559986, 
    4.566244, 4.584049, 4.600141, 4.617733, 4.622046, 4.642679, 4.625878, 
    4.653627, 4.630029, 4.670934, 4.597624, 4.629334, 4.572002, 4.578153, 
    4.589294, 4.614923, 4.601073, 4.617273, 4.581552, 4.563101, 4.558336, 
    4.549456, 4.558539, 4.557799, 4.566503, 4.563704, 4.584641, 4.573386, 
    4.605415, 4.617145, 4.650391, 4.670858, 4.691759, 4.701008, 4.703825, 
    4.705004,
  5.614617, 5.637631, 5.633152, 5.651754, 5.641429, 5.653619, 5.619277, 
    5.638547, 5.626239, 5.616685, 5.687986, 5.652586, 5.724919, 5.702219, 
    5.759362, 5.721383, 5.767041, 5.758262, 5.784709, 5.777124, 5.81105, 
    5.788213, 5.828689, 5.80559, 5.8092, 5.787461, 5.659695, 5.683571, 
    5.658283, 5.661682, 5.660156, 5.641643, 5.632331, 5.61286, 5.616391, 
    5.630693, 5.663211, 5.652156, 5.680044, 5.679413, 5.710576, 5.69651, 
    5.74907, 5.734096, 5.77744, 5.766518, 5.776927, 5.773769, 5.776968, 
    5.760956, 5.767813, 5.753736, 5.699143, 5.715149, 5.667507, 5.639002, 
    5.620121, 5.606753, 5.608641, 5.612243, 5.630776, 5.648241, 5.661576, 
    5.67051, 5.679322, 5.706062, 5.720246, 5.752102, 5.746342, 5.756101, 
    5.765432, 5.781126, 5.77854, 5.785462, 5.755842, 5.775516, 5.743063, 
    5.751927, 5.681727, 5.655137, 5.643868, 5.634013, 5.610094, 5.626604, 
    5.620091, 5.635593, 5.64546, 5.640578, 5.670754, 5.659009, 5.721088, 
    5.694289, 5.764343, 5.747524, 5.76838, 5.75773, 5.775987, 5.759554, 
    5.788039, 5.794256, 5.790007, 5.806337, 5.758645, 5.776928, 5.640442, 
    5.641238, 5.644947, 5.628657, 5.627661, 5.612763, 5.626018, 5.631669, 
    5.646032, 5.654541, 5.662639, 5.680471, 5.700437, 5.728437, 5.748613, 
    5.762166, 5.753852, 5.761192, 5.752988, 5.749145, 5.791926, 5.767877, 
    5.803986, 5.801983, 5.785627, 5.802209, 5.641797, 5.637217, 5.621339, 
    5.633762, 5.611142, 5.623796, 5.631083, 5.659256, 5.665458, 5.671216, 
    5.682597, 5.697229, 5.722963, 5.745421, 5.765975, 5.764467, 5.764998, 
    5.769597, 5.758211, 5.771468, 5.773696, 5.767873, 5.801715, 5.792033, 
    5.801941, 5.795635, 5.638705, 5.646414, 5.642248, 5.650084, 5.644563, 
    5.669147, 5.676532, 5.711182, 5.696941, 5.719615, 5.699241, 5.702848, 
    5.720359, 5.70034, 5.744182, 5.714436, 5.769776, 5.739979, 5.771647, 
    5.765886, 5.775426, 5.78398, 5.794753, 5.81467, 5.810053, 5.826736, 
    5.65792, 5.667945, 5.667061, 5.677564, 5.685342, 5.702223, 5.729376, 
    5.719154, 5.737928, 5.741703, 5.713183, 5.730683, 5.674661, 5.683687, 
    5.678311, 5.658711, 5.72151, 5.68922, 5.748947, 5.731378, 5.78276, 
    5.757167, 5.807513, 5.829134, 5.849526, 5.873429, 5.673421, 5.666603, 
    5.678814, 5.695743, 5.711478, 5.732449, 5.734597, 5.738533, 5.748735, 
    5.757325, 5.739779, 5.75948, 5.685785, 5.724319, 5.664028, 5.682136, 
    5.694743, 5.689209, 5.717986, 5.724784, 5.752469, 5.738145, 5.823793, 
    5.78579, 5.89167, 5.861947, 5.664222, 5.673397, 5.705413, 5.690164, 
    5.73385, 5.74464, 5.753422, 5.764663, 5.765877, 5.772546, 5.761621, 
    5.772113, 5.732493, 5.750175, 5.701746, 5.713507, 5.708094, 5.702161, 
    5.720485, 5.740056, 5.740472, 5.746758, 5.764503, 5.734027, 5.828716, 
    5.770113, 5.683414, 5.701141, 5.703674, 5.6968, 5.743558, 5.726584, 
    5.772383, 5.759979, 5.780312, 5.770202, 5.768716, 5.755751, 5.747691, 
    5.727363, 5.71086, 5.697796, 5.700832, 5.715188, 5.741253, 5.765988, 
    5.760563, 5.778765, 5.730674, 5.750806, 5.74302, 5.763337, 5.718883, 
    5.75673, 5.709239, 5.713391, 5.726248, 5.752175, 5.757918, 5.76406, 
    5.760269, 5.741916, 5.738912, 5.725935, 5.722357, 5.712486, 5.704325, 
    5.711782, 5.719621, 5.741923, 5.762074, 5.784102, 5.789501, 5.815336, 
    5.794302, 5.829044, 5.799502, 5.850704, 5.758925, 5.798631, 5.726833, 
    5.734537, 5.748492, 5.780586, 5.763241, 5.783528, 5.738794, 5.715685, 
    5.709714, 5.69859, 5.709969, 5.709043, 5.719944, 5.716439, 5.742664, 
    5.728567, 5.768679, 5.783367, 5.824986, 5.850606, 5.876761, 5.888336, 
    5.891861, 5.893336,
  8.093345, 8.127498, 8.120849, 8.148464, 8.133135, 8.151232, 8.100258, 
    8.128858, 8.11059, 8.096413, 8.202277, 8.149697, 8.257166, 8.223423, 
    8.30839, 8.25191, 8.319815, 8.306752, 8.346107, 8.334817, 8.385321, 
    8.35132, 8.41159, 8.37719, 8.382565, 8.350202, 8.160254, 8.195717, 
    8.158157, 8.163205, 8.160939, 8.133452, 8.119631, 8.090736, 8.095975, 
    8.1172, 8.165476, 8.14906, 8.190476, 8.189539, 8.235845, 8.214941, 
    8.293079, 8.27081, 8.335288, 8.319036, 8.334524, 8.329824, 8.334585, 
    8.31076, 8.320962, 8.300019, 8.218853, 8.242642, 8.171855, 8.129533, 
    8.101511, 8.081676, 8.084478, 8.089822, 8.117324, 8.143247, 8.163048, 
    8.176315, 8.189404, 8.229136, 8.250219, 8.297589, 8.289021, 8.303538, 
    8.31742, 8.340772, 8.336925, 8.347226, 8.303152, 8.332424, 8.284145, 
    8.297328, 8.192978, 8.153485, 8.136757, 8.122127, 8.086633, 8.111132, 
    8.101467, 8.124473, 8.139119, 8.131872, 8.176679, 8.159236, 8.251471, 
    8.21164, 8.3158, 8.290779, 8.321805, 8.305962, 8.333124, 8.308675, 
    8.351062, 8.360315, 8.353992, 8.378302, 8.307322, 8.334525, 8.131669, 
    8.132851, 8.138356, 8.114178, 8.1127, 8.090593, 8.110261, 8.118649, 
    8.139968, 8.152601, 8.164625, 8.191112, 8.220776, 8.262397, 8.292399, 
    8.31256, 8.300193, 8.31111, 8.298906, 8.293191, 8.356848, 8.321057, 
    8.374802, 8.371819, 8.347472, 8.372156, 8.13368, 8.126883, 8.103318, 
    8.121755, 8.088189, 8.106965, 8.117778, 8.159602, 8.168812, 8.177363, 
    8.194269, 8.216009, 8.254259, 8.287652, 8.318228, 8.315984, 8.316773, 
    8.323617, 8.306676, 8.326401, 8.329716, 8.321052, 8.371421, 8.357006, 
    8.371757, 8.362369, 8.129091, 8.140535, 8.13435, 8.145985, 8.137788, 
    8.174291, 8.185261, 8.236746, 8.215582, 8.249282, 8.218999, 8.22436, 
    8.250388, 8.220633, 8.28581, 8.241582, 8.323883, 8.27956, 8.326667, 
    8.318095, 8.33229, 8.34502, 8.361055, 8.39071, 8.383835, 8.40868, 
    8.157618, 8.172506, 8.171192, 8.186793, 8.198347, 8.223431, 8.263792, 
    8.248595, 8.276508, 8.282123, 8.239719, 8.265736, 8.182481, 8.195889, 
    8.187902, 8.158793, 8.252098, 8.204109, 8.292896, 8.266768, 8.343204, 
    8.305124, 8.380053, 8.412252, 8.442634, 8.47826, 8.180639, 8.170512, 
    8.188649, 8.2138, 8.237185, 8.268361, 8.271555, 8.277408, 8.292582, 
    8.305358, 8.279262, 8.308563, 8.199006, 8.256273, 8.166688, 8.193585, 
    8.212316, 8.204092, 8.246859, 8.256966, 8.298136, 8.276832, 8.404299, 
    8.347714, 8.505456, 8.461143, 8.166977, 8.180603, 8.228171, 8.20551, 
    8.270444, 8.286491, 8.299552, 8.316277, 8.318082, 8.328004, 8.311749, 
    8.327361, 8.268428, 8.294723, 8.22272, 8.2402, 8.232155, 8.223338, 
    8.250573, 8.279673, 8.280292, 8.28964, 8.316038, 8.270708, 8.411631, 
    8.324386, 8.195482, 8.221823, 8.225586, 8.215372, 8.284882, 8.259642, 
    8.327762, 8.309307, 8.339561, 8.324516, 8.322305, 8.303018, 8.291028, 
    8.260798, 8.236266, 8.216852, 8.221363, 8.242701, 8.281454, 8.318247, 
    8.310177, 8.337258, 8.265722, 8.295661, 8.284081, 8.314302, 8.248192, 
    8.304474, 8.233856, 8.240028, 8.259142, 8.297698, 8.306241, 8.315378, 
    8.309738, 8.282439, 8.277972, 8.258676, 8.253356, 8.238684, 8.226554, 
    8.237637, 8.24929, 8.28245, 8.312425, 8.345202, 8.353237, 8.391703, 
    8.360385, 8.41212, 8.368128, 8.44439, 8.307739, 8.366829, 8.260011, 
    8.271465, 8.29222, 8.33997, 8.31416, 8.344348, 8.277797, 8.243439, 
    8.234563, 8.218032, 8.234941, 8.233565, 8.24977, 8.244559, 8.283552, 
    8.262589, 8.32225, 8.344109, 8.406075, 8.444242, 8.483227, 8.500484, 
    8.505741, 8.50794,
  12.6655, 12.72096, 12.71016, 12.75503, 12.73012, 12.75953, 12.67672, 
    12.72317, 12.6935, 12.67048, 12.84254, 12.75704, 12.9319, 12.87696, 
    13.01538, 12.92334, 13.03401, 13.01271, 13.07691, 13.05849, 13.14093, 
    13.08542, 13.18384, 13.12765, 13.13643, 13.08359, 12.7742, 12.83187, 
    12.77079, 12.779, 12.77531, 12.73064, 12.70819, 12.66126, 12.66977, 
    12.70424, 12.78269, 12.756, 12.82334, 12.82182, 12.89718, 12.86315, 
    12.99042, 12.95413, 13.05925, 13.03274, 13.05801, 13.05034, 13.05811, 
    13.01925, 13.03588, 13.00173, 12.86952, 12.90825, 12.79306, 12.72427, 
    12.67876, 12.64656, 12.6511, 12.65978, 12.70444, 12.74655, 12.77874, 
    12.80031, 12.8216, 12.88626, 12.92058, 12.99777, 12.98381, 13.00747, 
    13.03011, 13.0682, 13.06192, 13.07873, 13.00684, 13.05458, 12.97586, 
    12.99735, 12.82741, 12.7632, 12.73601, 12.71224, 12.6546, 12.69438, 
    12.67869, 12.71605, 12.73985, 12.72807, 12.8009, 12.77254, 12.92262, 
    12.85778, 13.02746, 12.98667, 13.03726, 13.01142, 13.05572, 13.01585, 
    13.08499, 13.1001, 13.08978, 13.12946, 13.01364, 13.05801, 12.72774, 
    12.72966, 12.73861, 12.69933, 12.69693, 12.66103, 12.69296, 12.70659, 
    12.74123, 12.76176, 12.7813, 12.82438, 12.87265, 12.94042, 12.98931, 
    13.02218, 13.00202, 13.01982, 12.99992, 12.9906, 13.09444, 13.03604, 
    13.12375, 13.11888, 13.07913, 13.11943, 12.73101, 12.71996, 12.68169, 
    12.71163, 12.65713, 12.68761, 12.70517, 12.77314, 12.78811, 12.80202, 
    12.82951, 12.86489, 12.92716, 12.98157, 13.03142, 13.02777, 13.02905, 
    13.04021, 13.01259, 13.04475, 13.05016, 13.03603, 13.11823, 13.0947, 
    13.11878, 13.10345, 12.72355, 12.74215, 12.7321, 12.751, 12.73768, 
    12.79702, 12.81486, 12.89864, 12.86419, 12.91906, 12.86975, 12.87848, 
    12.92086, 12.87241, 12.97857, 12.90652, 13.04065, 12.96838, 13.04519, 
    13.03121, 13.05436, 13.07513, 13.10131, 13.14973, 13.1385, 13.17909, 
    12.76991, 12.79412, 12.79198, 12.81735, 12.83615, 12.87697, 12.94269, 
    12.91794, 12.96341, 12.97256, 12.90349, 12.94586, 12.81034, 12.83215, 
    12.81916, 12.77182, 12.92365, 12.84552, 12.99012, 12.94754, 13.07217, 
    13.01006, 13.13233, 13.18493, 13.23459, 13.29288, 12.80734, 12.79088, 
    12.82037, 12.86129, 12.89936, 12.95014, 12.95534, 12.96488, 12.98961, 
    13.01044, 12.9679, 13.01566, 12.83722, 12.93044, 12.78466, 12.8284, 
    12.85888, 12.8455, 12.91511, 12.93157, 12.99866, 12.96394, 13.17193, 
    13.07953, 13.3374, 13.26487, 12.78513, 12.80728, 12.88468, 12.8478, 
    12.95353, 12.97968, 13.00097, 13.02824, 13.03119, 13.04737, 13.02086, 
    13.04632, 12.95024, 12.9931, 12.87581, 12.90427, 12.89117, 12.87682, 
    12.92116, 12.96857, 12.96958, 12.98481, 13.02785, 12.95396, 13.18391, 
    13.04147, 12.83149, 12.87435, 12.88048, 12.86385, 12.97706, 12.93593, 
    13.04698, 13.01688, 13.06623, 13.04168, 13.03807, 13.00662, 12.98708, 
    12.93782, 12.89786, 12.86626, 12.8736, 12.90834, 12.97147, 13.03146, 
    13.01829, 13.06247, 12.94584, 12.99463, 12.97575, 13.02502, 12.91728, 
    13.009, 12.89394, 12.90399, 12.93512, 12.99795, 13.01188, 13.02678, 
    13.01758, 12.97308, 12.9658, 12.93436, 12.92569, 12.9018, 12.88205, 
    12.90009, 12.91907, 12.97309, 13.02196, 13.07543, 13.08854, 13.15135, 
    13.10021, 13.18471, 13.11285, 13.23747, 13.01432, 13.11073, 12.93653, 
    12.95519, 12.98902, 13.06689, 13.02479, 13.07404, 12.96551, 12.90954, 
    12.89509, 12.86818, 12.89571, 12.89347, 12.91985, 12.91137, 12.97489, 
    12.94073, 13.03799, 13.07365, 13.17483, 13.23722, 13.301, 13.32926, 
    13.33786, 13.34147,
  20.5999, 20.69597, 20.67725, 20.75503, 20.71184, 20.76283, 20.61933, 
    20.6998, 20.64838, 20.60852, 20.90694, 20.75851, 21.06235, 20.96676, 
    21.20782, 21.04745, 21.24033, 21.20317, 21.31521, 21.28304, 21.42711, 
    21.33008, 21.50221, 21.40389, 21.41924, 21.32689, 20.78827, 20.8884, 
    20.78236, 20.7966, 20.79021, 20.71273, 20.67382, 20.59257, 20.60729, 
    20.66698, 20.80301, 20.75671, 20.87359, 20.87094, 21.00193, 20.94275, 
    21.1643, 21.10106, 21.28439, 21.23811, 21.28221, 21.26883, 21.28238, 
    21.21457, 21.24359, 21.18402, 20.95382, 21.02118, 20.82101, 20.7017, 
    20.62285, 20.56712, 20.57499, 20.59, 20.66733, 20.74033, 20.79615, 
    20.8336, 20.87056, 20.98293, 21.04266, 21.17712, 21.15277, 21.19403, 
    21.23351, 21.30001, 21.28905, 21.3184, 21.19293, 21.27623, 21.13892, 
    21.17638, 20.88066, 20.76919, 20.72204, 20.68085, 20.58104, 20.64991, 
    20.62273, 20.68745, 20.7287, 20.70828, 20.83462, 20.7854, 21.04621, 
    20.93341, 21.2289, 21.15777, 21.24599, 21.20092, 21.27822, 21.20864, 
    21.32934, 21.35573, 21.33769, 21.40706, 21.20479, 21.28222, 20.70771, 
    20.71104, 20.72655, 20.65848, 20.65432, 20.59217, 20.64746, 20.67106, 
    20.73109, 20.7667, 20.8006, 20.87538, 20.95926, 21.07719, 21.16237, 
    21.21969, 21.18452, 21.21556, 21.18086, 21.16462, 21.34584, 21.24387, 
    21.39707, 21.38856, 21.3191, 21.38952, 20.71338, 20.69423, 20.62794, 
    20.6798, 20.58541, 20.63819, 20.66861, 20.78644, 20.81242, 20.83655, 
    20.88431, 20.94578, 21.05411, 21.14888, 21.23581, 21.22943, 21.23168, 
    21.25115, 21.20295, 21.25908, 21.26852, 21.24385, 21.38742, 21.34629, 
    21.38838, 21.36159, 20.70045, 20.73269, 20.71526, 20.74804, 20.72495, 
    20.82788, 20.85885, 21.00448, 20.94457, 21.04, 20.95424, 20.9694, 
    21.04313, 20.95886, 21.14365, 21.01818, 21.25191, 21.1259, 21.25983, 
    21.23544, 21.27585, 21.31212, 21.35784, 21.44251, 21.42287, 21.49389, 
    20.78084, 20.82284, 20.81914, 20.86318, 20.89583, 20.96678, 21.08115, 
    21.03805, 21.11724, 21.13317, 21.0129, 21.08666, 20.851, 20.88888, 
    20.86632, 20.78415, 21.04798, 20.91212, 21.16378, 21.08959, 21.30694, 
    21.19854, 21.41207, 21.50411, 21.59112, 21.69336, 20.8458, 20.81721, 
    20.86843, 20.93953, 21.00572, 21.09411, 21.10317, 21.11979, 21.16289, 
    21.19921, 21.12505, 21.20832, 20.89769, 21.05982, 20.80643, 20.88237, 
    20.93533, 20.91207, 21.03313, 21.06178, 21.17867, 21.11815, 21.48136, 
    21.3198, 21.77154, 21.64421, 20.80724, 20.8457, 20.9802, 20.91608, 
    21.10002, 21.14558, 21.1827, 21.23026, 21.2354, 21.26364, 21.21738, 
    21.26181, 21.0943, 21.16897, 20.96477, 21.01427, 20.99148, 20.96651, 
    21.04366, 21.12622, 21.12798, 21.15453, 21.22958, 21.10077, 21.50233, 
    21.25334, 20.88773, 20.96223, 20.97288, 20.94397, 21.14101, 21.06938, 
    21.26295, 21.21043, 21.29656, 21.25371, 21.24742, 21.19255, 21.15847, 
    21.07266, 21.00312, 20.94816, 20.96092, 21.02135, 21.13128, 21.23587, 
    21.21291, 21.29, 21.08662, 21.17164, 21.13874, 21.22465, 21.03691, 
    21.19669, 20.99629, 21.01378, 21.06796, 21.17743, 21.20172, 21.22771, 
    21.21166, 21.13408, 21.12139, 21.06664, 21.05155, 21.00997, 20.97562, 
    21.007, 21.04002, 21.1341, 21.2193, 21.31264, 21.33554, 21.44535, 
    21.35593, 21.50373, 21.37802, 21.59616, 21.20597, 21.37431, 21.07042, 
    21.10292, 21.16186, 21.29772, 21.22424, 21.3102, 21.12089, 21.02344, 
    20.9983, 20.9515, 20.99937, 20.99547, 21.04138, 21.02662, 21.13724, 
    21.07773, 21.24726, 21.30952, 21.48644, 21.59573, 21.70762, 21.75724, 
    21.77237, 21.77869,
  34.64178, 34.82255, 34.7873, 34.9339, 34.85246, 34.94861, 34.67831, 
    34.82977, 34.73297, 34.65799, 35.22099, 34.94045, 35.51581, 35.33433, 
    35.79281, 35.48749, 35.85484, 35.78393, 35.99794, 35.93643, 36.21229, 
    36.02638, 36.3565, 36.16775, 36.19719, 36.02027, 34.99663, 35.18589, 
    34.98547, 35.01235, 35.00028, 34.85415, 34.78085, 34.62801, 34.65568, 
    34.76797, 35.02445, 34.93707, 35.15787, 35.15286, 35.40105, 35.28883, 
    35.70983, 35.58942, 35.939, 35.85061, 35.93484, 35.90927, 35.93517, 
    35.80567, 35.86107, 35.74742, 35.30981, 35.4376, 35.05845, 34.83335, 
    34.68494, 34.5802, 34.59498, 34.62318, 34.76862, 34.90616, 35.01151, 
    35.08224, 35.15214, 35.365, 35.47839, 35.73426, 35.68786, 35.76649, 
    35.84183, 35.96887, 35.94791, 36.00405, 35.7644, 35.92341, 35.66148, 
    35.73284, 35.17124, 34.96061, 34.87169, 34.79408, 34.60635, 34.73584, 
    34.68471, 34.80651, 34.88423, 34.84576, 35.08418, 34.99121, 35.48513, 
    35.27113, 35.83303, 35.69738, 35.86566, 35.77964, 35.92722, 35.79436, 
    36.02497, 36.07548, 36.04095, 36.17384, 35.78701, 35.93485, 34.84468, 
    34.85095, 34.88018, 34.75196, 34.74414, 34.62725, 34.73122, 34.77564, 
    34.88874, 34.9559, 35.01992, 35.16126, 35.32012, 35.54401, 35.70615, 
    35.81544, 35.74836, 35.80758, 35.74139, 35.71043, 36.05655, 35.8616, 
    36.15468, 36.13837, 36.00539, 36.14021, 34.85536, 34.81929, 34.6945, 
    34.7921, 34.61456, 34.71379, 34.77103, 34.99316, 35.04223, 35.08783, 
    35.17815, 35.29456, 35.50014, 35.68045, 35.84622, 35.83403, 35.83832, 
    35.8755, 35.78352, 35.89064, 35.90867, 35.86156, 36.13618, 36.05741, 
    36.13802, 36.0867, 34.83101, 34.89175, 34.85891, 34.92071, 34.87716, 
    35.07144, 35.13, 35.40589, 35.29227, 35.47334, 35.31059, 35.33935, 
    35.4793, 35.31936, 35.67049, 35.4319, 35.87695, 35.63669, 35.89209, 
    35.8455, 35.92268, 35.99202, 36.07952, 36.24183, 36.20415, 36.3405, 
    34.9826, 35.06193, 35.05492, 35.13819, 35.19995, 35.33437, 35.55154, 
    35.46964, 35.6202, 35.65054, 35.42188, 35.56203, 35.11515, 35.18681, 
    35.14411, 34.98885, 35.48851, 35.23079, 35.70884, 35.5676, 35.98212, 
    35.7751, 36.18343, 36.36015, 36.52758, 36.7248, 35.10532, 35.05129, 
    35.1481, 35.28271, 35.40826, 35.5762, 35.59344, 35.62506, 35.70713, 
    35.77637, 35.63507, 35.79375, 35.20348, 35.511, 35.03091, 35.17449, 
    35.27475, 35.23071, 35.4603, 35.51473, 35.73721, 35.62194, 36.31643, 
    36.00671, 36.876, 36.62993, 35.03245, 35.10513, 35.35982, 35.2383, 
    35.58744, 35.67417, 35.74489, 35.83562, 35.84542, 35.89936, 35.81104, 
    35.89586, 35.57656, 35.71872, 35.33056, 35.42447, 35.38122, 35.33387, 
    35.48029, 35.6373, 35.64064, 35.69121, 35.83432, 35.58887, 36.35673, 
    35.87968, 35.18463, 35.32574, 35.34594, 35.29114, 35.66546, 35.52916, 
    35.89804, 35.79779, 35.96227, 35.8804, 35.86837, 35.76368, 35.69872, 
    35.5354, 35.40331, 35.29908, 35.32327, 35.43792, 35.64693, 35.84632, 
    35.80251, 35.94973, 35.56196, 35.72381, 35.66113, 35.8249, 35.46747, 
    35.77157, 35.39036, 35.42354, 35.52646, 35.73484, 35.78116, 35.83075, 
    35.80013, 35.65226, 35.62811, 35.52395, 35.49529, 35.41631, 35.35114, 
    35.41068, 35.47338, 35.65231, 35.81471, 35.99301, 36.03684, 36.24728, 
    36.07586, 36.35942, 36.11818, 36.53728, 35.78928, 36.11107, 35.53115, 
    35.59296, 35.70518, 35.96449, 35.82413, 35.98835, 35.62716, 35.44189, 
    35.39416, 35.3054, 35.39619, 35.3888, 35.47597, 35.44792, 35.65827, 
    35.54505, 35.86808, 35.98705, 36.32619, 36.53647, 36.75237, 36.84832, 
    36.87759, 36.88984,
  60.67866, 61.07138, 60.99464, 61.31427, 61.13654, 61.34644, 60.75787, 
    61.08709, 60.87651, 60.71379, 61.94415, 61.3286, 62.59654, 62.19429, 
    63.21474, 62.53363, 63.35389, 63.19484, 63.67592, 63.53733, 64.16097, 
    63.74009, 64.48915, 64.05992, 64.12669, 63.72631, 61.45146, 61.86686, 
    61.42703, 61.48588, 61.45945, 61.14022, 60.9806, 60.64882, 60.70879, 
    60.95258, 61.51238, 61.32119, 61.80522, 61.7942, 62.34192, 62.09377, 
    63.02899, 62.76031, 63.54311, 63.34439, 63.53375, 63.4762, 63.5345, 
    63.24357, 63.36789, 63.11309, 62.1401, 62.42293, 61.58691, 61.09489, 
    60.77224, 60.54533, 60.5773, 60.63837, 60.95401, 61.2537, 61.48405, 
    61.6391, 61.79262, 62.26212, 62.51342, 63.08363, 62.97991, 63.15579, 
    63.32469, 63.61038, 63.56317, 63.68969, 63.15111, 63.50803, 62.92099, 
    63.08046, 61.83464, 61.37265, 61.17846, 61.00938, 60.60192, 60.88274, 
    60.77174, 61.03644, 61.20583, 61.12193, 61.64335, 61.4396, 62.52837, 
    62.05472, 63.30494, 63.00117, 63.37819, 63.18523, 63.5166, 63.21821, 
    63.7369, 63.85101, 63.77299, 64.07372, 63.20175, 63.53376, 61.11959, 
    61.13326, 61.197, 60.91779, 60.90078, 60.64719, 60.87272, 60.96927, 
    61.21567, 61.36237, 61.50245, 61.81269, 62.16289, 62.65925, 63.02077, 
    63.26548, 63.11519, 63.24784, 63.0996, 63.03035, 63.80822, 63.36906, 
    64.03029, 63.99333, 63.69271, 63.99749, 61.14286, 61.06427, 60.79298, 
    61.00508, 60.61969, 60.83485, 60.95924, 61.44387, 61.55134, 61.65136, 
    61.84983, 62.10643, 62.56173, 62.96335, 63.33453, 63.30719, 63.31681, 
    63.40031, 63.19391, 63.43432, 63.47487, 63.36899, 63.98838, 63.81017, 
    63.99254, 63.87637, 61.08979, 61.22225, 61.1506, 61.28547, 61.19041, 
    61.6154, 61.74396, 62.35265, 62.10136, 62.5022, 62.14183, 62.20539, 
    62.51543, 62.16119, 62.9411, 62.41028, 63.40356, 62.86567, 63.43758, 
    63.33292, 63.50638, 63.66257, 63.86015, 64.22809, 64.14249, 64.45267, 
    61.42075, 61.59453, 61.57916, 61.76195, 61.89783, 62.19437, 62.67599, 
    62.494, 62.8289, 62.89658, 62.38808, 62.69933, 61.71135, 61.86889, 
    61.77497, 61.43444, 62.53588, 61.96577, 63.02679, 62.71173, 63.64025, 
    63.17506, 64.09548, 64.49747, 64.88044, 65.3342, 61.68975, 61.57121, 
    61.78375, 62.08028, 62.35789, 62.73087, 62.76926, 62.83974, 63.02298, 
    63.1779, 62.86208, 63.21685, 61.9056, 62.58585, 61.52654, 61.84178, 
    62.06271, 61.96557, 62.47326, 62.59414, 63.09025, 62.83279, 64.3978, 
    63.6957, 65.68405, 65.11556, 61.5299, 61.68932, 62.25066, 61.98231, 
    62.75591, 62.94933, 63.10743, 63.31075, 63.33276, 63.45393, 63.25561, 
    63.44606, 62.73167, 63.04889, 62.18595, 62.39381, 62.298, 62.19328, 
    62.51765, 62.86703, 62.87449, 62.9874, 63.30784, 62.75908, 64.48967, 
    63.4097, 61.8641, 62.17531, 62.21996, 62.09887, 62.92989, 62.62622, 
    63.45097, 63.22589, 63.59551, 63.4113, 63.38429, 63.14947, 63.00418, 
    62.64008, 62.34694, 62.1164, 62.16985, 62.42362, 62.88852, 63.33477, 
    63.23648, 63.56726, 62.69917, 63.06026, 62.92022, 63.2867, 62.48919, 
    63.16716, 62.31825, 62.39175, 62.62022, 63.08494, 63.18863, 63.2998, 
    63.23115, 62.90041, 62.84653, 62.61464, 62.55093, 62.37573, 62.23145, 
    62.36326, 62.5023, 62.90052, 63.26383, 63.6648, 63.7637, 64.24046, 
    63.85188, 64.4958, 63.9476, 64.90269, 63.20683, 63.93153, 62.63064, 
    62.7682, 63.0186, 63.60052, 63.28497, 63.6543, 62.84442, 62.43243, 
    62.32666, 62.13037, 62.33117, 62.31479, 62.50804, 62.4458, 62.91383, 
    62.66155, 63.38363, 63.65136, 64.42004, 64.90083, 65.39787, 65.61987, 
    65.68774, 65.71616,
  116.3177, 117.5456, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.1711, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3958, 122.2342, 124.1728, 123.8164, 124.4217, 
    125.0078, 126.01, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.8839, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4582, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9566, 
    124.8018, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.3901, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3966, 123.7596, 125.0421, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2484, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6645, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7011, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3602, 121.7737, 121.2941, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8678, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1653, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.0212997, -0.02095049, -0.0210179, -0.0207397, -0.02089354, -0.02071207, 
    -0.02122841, -0.02093674, -0.02112245, -0.02126801, -0.02021082, 
    -0.02072738, -0.01968869, -0.02000757, -0.01921673, -0.01973795, 
    -0.01911341, -0.01923157, -0.0188783, -0.0189788, -0.01853446, 
    -0.01883211, -0.0183085, -0.01860509, -0.01855835, -0.01884201, 
    -0.02062232, -0.02027438, -0.02064313, -0.02059308, -0.02061552, 
    -0.02089035, -0.0210303, -0.02132664, -0.02127252, -0.02105502, 
    -0.02057061, -0.02073372, -0.02032526, -0.02033439, -0.01988942, 
    -0.02008876, -0.01935626, -0.01956153, -0.01897459, -0.01912041, 
    -0.01898141, -0.01902345, -0.01898086, -0.01919522, -0.01910306, 
    -0.01929284, -0.02005126, -0.01982514, -0.02050765, -0.02092995, 
    -0.02121552, -0.02142066, -0.02139153, -0.02133612, -0.02105376, 
    -0.02079188, -0.02059462, -0.02046377, -0.0203357, -0.01995317, 
    -0.01975381, -0.01931503, -0.01939345, -0.0192608, -0.01913499, 
    -0.01892571, -0.01895999, -0.01886838, -0.01926429, -0.01900019, 
    -0.01943827, -0.01931739, -0.020301, -0.02068959, -0.0208571, 
    -0.02100492, -0.02136916, -0.02111692, -0.02121598, -0.02098112, 
    -0.0208333, -0.02090627, -0.0204602, -0.02063242, -0.01974206, 
    -0.02012048, -0.01914962, -0.01937733, -0.01909546, -0.01923874, 
    -0.01899393, -0.01921411, -0.01883441, -0.01875279, -0.01880852, 
    -0.01859539, -0.01922639, -0.01898141, -0.02090832, -0.0208964, 
    -0.02084096, -0.02108582, -0.0211009, -0.02132813, -0.02112581, 
    -0.02104027, -0.02082477, -0.02069839, -0.02057901, -0.02031908, 
    -0.02003288, -0.01963981, -0.01936248, -0.0191789, -0.01929125, 
    -0.01919203, -0.01930298, -0.01935522, -0.01878332, -0.0191022, 
    -0.01862588, -0.01865191, -0.0188662, -0.01864897, -0.02088803, 
    -0.0209567, -0.02119695, -0.02100869, -0.02135303, -0.02115955, 
    -0.02104914, -0.0206288, -0.02053764, -0.02045349, -0.02028836, 
    -0.0200785, -0.01971589, -0.01940604, -0.01912769, -0.01914795, 
    -0.01914081, -0.01907917, -0.01923225, -0.01905416, -0.01902444, 
    -0.01910225, -0.0186554, -0.01878191, -0.01865246, -0.01873472, 
    -0.02093435, -0.02081908, -0.02088129, -0.02076447, -0.02084669, 
    -0.0204837, -0.02037617, -0.0198809, -0.02008261, -0.01976261, 
    -0.02004986, -0.01999864, -0.01975225, -0.02003423, -0.01942298, 
    -0.01983518, -0.01907677, -0.01948059, -0.01905177, -0.01912889, 
    -0.01900138, -0.01888795, -0.01874627, -0.01848779, -0.01854731, 
    -0.01833334, -0.02064848, -0.02050124, -0.02051417, -0.02036117, 
    -0.0202488, -0.02000749, -0.01962679, -0.01976905, -0.01950873, 
    -0.01945691, -0.01985273, -0.0196087, -0.02040333, -0.02027266, 
    -0.02035036, -0.02063682, -0.01973616, -0.02019307, -0.01935793, 
    -0.01959907, -0.01890408, -0.01924637, -0.01858016, -0.01830287, 
    -0.01804595, -0.01775054, -0.02042136, -0.02052087, -0.02034306, 
    -0.02009972, -0.01987671, -0.01958427, -0.01955462, -0.01950042, 
    -0.0193608, -0.01924423, -0.01948332, -0.01921512, -0.02024247, 
    -0.01969702, -0.02055862, -0.02029505, -0.02011398, -0.02019321, 
    -0.01978538, -0.01969053, -0.01931004, -0.01950575, -0.01837089, 
    -0.01886407, -0.01752911, -0.01789171, -0.02055576, -0.02042171, 
    -0.01996231, -0.02017951, -0.01956492, -0.0194167, -0.01929709, 
    -0.01914532, -0.01912902, -0.01903977, -0.01918624, -0.01904554, 
    -0.01958366, -0.01934122, -0.02001427, -0.01984819, -0.01992441, 
    -0.02000837, -0.01975045, -0.01947953, -0.01947379, -0.01938778, 
    -0.01914756, -0.01956247, -0.01830822, -0.01907233, -0.02027658, 
    -0.02002288, -0.01998693, -0.02008461, -0.0194315, -0.01966551, 
    -0.01904194, -0.01920838, -0.01893649, -0.01907108, -0.01909096, 
    -0.01926552, -0.01937504, -0.01965471, -0.01988542, -0.02007042, 
    -0.02002724, -0.01982459, -0.01946308, -0.01912753, -0.01920051, 
    -0.018957, -0.01960881, -0.01933264, -0.01943888, -0.01916315, 
    -0.01977284, -0.01925235, -0.01990826, -0.01984981, -0.01967018, 
    -0.01931405, -0.0192362, -0.01915343, -0.01920446, -0.019454, 
    -0.01949522, -0.01967453, -0.01972434, -0.01986253, -0.0199777, 
    -0.01987244, -0.01976253, -0.0194539, -0.01918014, -0.01888634, 
    -0.01881517, -0.01847926, -0.0187522, -0.01830406, -0.01868431, 
    -0.01803131, -0.01922265, -0.01869564, -0.01966205, -0.01955544, 
    -0.01936414, -0.01893288, -0.01916443, -0.01889393, -0.01949683, 
    -0.01981763, -0.01990155, -0.02005912, -0.01989797, -0.01991102, 
    -0.019758, -0.01980704, -0.01944374, -0.019638, -0.01909146, -0.01889606, 
    -0.01835564, -0.0180325, -0.01770981, -0.01756931, -0.01752679, 
    -0.01750904,
  -0.05476891, -0.0537186, -0.05392112, -0.05308613, -0.05354765, 
    -0.05300333, -0.05455427, -0.0536773, -0.05423543, -0.05467353, 
    -0.05150439, -0.05304921, -0.04995042, -0.05089871, -0.04855207, 
    -0.05009669, -0.0482468, -0.048596, -0.04755323, -0.04784952, 
    -0.04654148, -0.04741713, -0.04587856, -0.04674907, -0.04661171, 
    -0.0474463, -0.05273452, -0.05169407, -0.05279684, -0.05264694, 
    -0.05271417, -0.05353804, -0.05395831, -0.05485014, -0.0546871, 
    -0.05403267, -0.05257969, -0.05306828, -0.05184618, -0.05187345, 
    -0.05054706, -0.0511406, -0.0489649, -0.04957313, -0.04783711, 
    -0.04826753, -0.04785722, -0.04798126, -0.04785561, -0.04848853, 
    -0.04821627, -0.04877722, -0.05102886, -0.05035588, -0.05239131, 
    -0.05365682, -0.05451547, -0.05513351, -0.05504569, -0.05487866, 
    -0.05402886, -0.05324265, -0.0526516, -0.0522601, -0.05187737, 
    -0.05073662, -0.05014383, -0.04884284, -0.04907503, -0.04868242, 
    -0.04831058, -0.04769294, -0.04779403, -0.04752396, -0.04869279, 
    -0.0479126, -0.04920779, -0.04884988, -0.05177351, -0.05293601, 
    -0.05343818, -0.05388211, -0.05497826, -0.05421878, -0.05451683, 
    -0.05381063, -0.0533669, -0.05358589, -0.05224944, -0.05276476, 
    -0.05010893, -0.05123511, -0.04835379, -0.04902728, -0.04819384, 
    -0.04861724, -0.04789413, -0.04854441, -0.04742388, -0.04718352, 
    -0.04734763, -0.0467206, -0.04858072, -0.0478572, -0.05359202, 
    -0.05355624, -0.05338988, -0.05412524, -0.05417059, -0.0548546, 
    -0.05424555, -0.05398835, -0.05334132, -0.0529624, -0.05260487, 
    -0.05182771, -0.05097406, -0.04980535, -0.04898332, -0.04844035, 
    -0.04877255, -0.04847913, -0.04880725, -0.04896186, -0.04727341, 
    -0.04821372, -0.04681024, -0.04688677, -0.04751755, -0.04687814, 
    -0.05353113, -0.05373731, -0.05445958, -0.05389347, -0.05492964, 
    -0.05434703, -0.05401497, -0.05275387, -0.05248107, -0.05222934, 
    -0.051736, -0.05111004, -0.05003124, -0.04911228, -0.04828905, 
    -0.04834887, -0.0483278, -0.04814572, -0.04859804, -0.04807189, 
    -0.04798415, -0.04821387, -0.04689702, -0.0472693, -0.0468884, 
    -0.04713039, -0.0536702, -0.05332423, -0.05351088, -0.05316045, 
    -0.05340705, -0.05231962, -0.05199817, -0.05052167, -0.05112227, 
    -0.05017002, -0.05102469, -0.05087212, -0.05013914, -0.05097814, 
    -0.04916242, -0.05038567, -0.04813866, -0.04933306, -0.04806483, 
    -0.04829258, -0.04791615, -0.04758163, -0.04716436, -0.04640451, 
    -0.04657931, -0.0459514, -0.05281287, -0.05237213, -0.05241084, 
    -0.05195345, -0.05161789, -0.05089851, -0.04976675, -0.05018919, 
    -0.0494166, -0.049263, -0.05043795, -0.04971302, -0.05207938, 
    -0.05168906, -0.05192113, -0.05277792, -0.05009143, -0.05145154, 
    -0.04896984, -0.0496845, -0.04762917, -0.04863975, -0.04667582, 
    -0.04586198, -0.04511005, -0.04424763, -0.0521333, -0.05243089, 
    -0.05189935, -0.05117322, -0.05050927, -0.04964058, -0.04955264, 
    -0.04939195, -0.04897837, -0.04863345, -0.04934121, -0.0485474, 
    -0.05159886, -0.04997521, -0.05254382, -0.05175588, -0.05121575, 
    -0.05145201, -0.05023773, -0.04995597, -0.04882808, -0.04940775, 
    -0.04606139, -0.04751121, -0.04360292, -0.04465941, -0.05253528, 
    -0.05213435, -0.05076393, -0.05141117, -0.04958319, -0.04914387, 
    -0.04878982, -0.04834108, -0.04829294, -0.04802942, -0.04846204, 
    -0.04804645, -0.04963876, -0.04892038, -0.0509187, -0.05042445, 
    -0.05065121, -0.05090114, -0.05013394, -0.04932996, -0.04931303, 
    -0.04905821, -0.04834748, -0.04957593, -0.04587755, -0.04812535, 
    -0.05170083, -0.05094425, -0.05083726, -0.05112827, -0.04918772, 
    -0.04988166, -0.04803584, -0.04852746, -0.04772474, -0.04812184, 
    -0.04818055, -0.04869642, -0.04902052, -0.0498496, -0.05053518, 
    -0.05108597, -0.05095734, -0.05035426, -0.04928125, -0.04828854, 
    -0.04850416, -0.04778525, -0.04971339, -0.04889497, -0.04920955, 
    -0.04839377, -0.05020045, -0.04865726, -0.05060314, -0.0504293, 
    -0.04989554, -0.04883992, -0.04860972, -0.04836504, -0.04851589, 
    -0.04925435, -0.04937651, -0.04990847, -0.05005636, -0.0504671, 
    -0.0508098, -0.05049656, -0.05016979, -0.04925407, -0.04844397, 
    -0.04757687, -0.04736723, -0.04637936, -0.04718173, -0.04586533, 
    -0.04698179, -0.04506709, -0.04856953, -0.04701524, -0.04987143, 
    -0.04955509, -0.0489882, -0.04771402, -0.04839757, -0.04759923, 
    -0.0493813, -0.05033354, -0.05058319, -0.05105228, -0.05057252, 
    -0.05061136, -0.05015637, -0.05030211, -0.04922397, -0.04980003, 
    -0.04818201, -0.0476055, -0.04601675, -0.04507068, -0.04412901, 
    -0.04371991, -0.04359621, -0.0435446,
  -0.07892428, -0.07727004, -0.07758883, -0.07627513, -0.07700105, 
    -0.07614495, -0.07858603, -0.07720505, -0.07808375, -0.07877396, 
    -0.073791, -0.07621709, -0.07135644, -0.07284144, -0.0691708, 
    -0.07158534, -0.06869433, -0.06923942, -0.06761269, -0.06807461, 
    -0.06603707, -0.0674006, -0.06500623, -0.06636015, -0.06614637, 
    -0.06744605, -0.07572243, -0.07408857, -0.07582036, -0.07558481, 
    -0.07569045, -0.07698593, -0.07764736, -0.07905233, -0.07879534, 
    -0.07776444, -0.07547913, -0.07624708, -0.07432733, -0.07437014, 
    -0.07229052, -0.07322058, -0.06981556, -0.07076627, -0.06805527, 
    -0.06872669, -0.06808663, -0.06828007, -0.06808411, -0.06907163, 
    -0.06864671, -0.0695224, -0.07304543, -0.07199111, -0.07518321, 
    -0.07717281, -0.0785249, -0.07949911, -0.07936063, -0.07909729, 
    -0.07775845, -0.07652127, -0.07559214, -0.07497714, -0.07437629, 
    -0.07258743, -0.07165914, -0.06962487, -0.06998763, -0.06937435, 
    -0.06879387, -0.06783047, -0.06798809, -0.06756707, -0.06939055, 
    -0.06817298, -0.07019511, -0.06963589, -0.07421324, -0.07603914, 
    -0.07682879, -0.07752742, -0.07925431, -0.07805751, -0.07852703, 
    -0.07741491, -0.07671668, -0.07706122, -0.0749604, -0.07576996, 
    -0.07160451, -0.07336874, -0.06886131, -0.06991302, -0.0686117, 
    -0.06927259, -0.06814418, -0.06915887, -0.06741111, -0.06703661, 
    -0.06729229, -0.06631586, -0.06921556, -0.06808658, -0.07707087, 
    -0.07701456, -0.07675284, -0.07791021, -0.07798163, -0.07905935, 
    -0.0780997, -0.07769466, -0.07667646, -0.07608062, -0.0755187, 
    -0.07429834, -0.07295953, -0.07112948, -0.06984434, -0.06899641, 
    -0.06951511, -0.06905696, -0.0695693, -0.06981082, -0.06717665, 
    -0.06864272, -0.06645539, -0.06657451, -0.06755707, -0.06656108, 
    -0.07697506, -0.0772995, -0.07843683, -0.0775453, -0.07917766, 
    -0.07825952, -0.07773657, -0.07575282, -0.07532421, -0.07492884, 
    -0.07415442, -0.07317267, -0.07148293, -0.07004584, -0.06876028, 
    -0.06885364, -0.06882075, -0.06853662, -0.0692426, -0.06842145, 
    -0.06828458, -0.06864296, -0.06659049, -0.06717025, -0.06657705, 
    -0.06695388, -0.07719389, -0.07664958, -0.0769432, -0.076392, 
    -0.07677985, -0.0750706, -0.07456587, -0.07225073, -0.07319184, 
    -0.07170014, -0.07303889, -0.07279976, -0.07165178, -0.07296593, 
    -0.07012418, -0.07203773, -0.0685256, -0.07039087, -0.06841043, 
    -0.06876578, -0.06817853, -0.06765696, -0.06700679, -0.06582401, 
    -0.06609597, -0.06511945, -0.07584558, -0.07515308, -0.07521389, 
    -0.0744957, -0.07396911, -0.07284113, -0.07106909, -0.07173017, 
    -0.07052151, -0.0702814, -0.07211965, -0.07098505, -0.07469337, 
    -0.07408075, -0.07444496, -0.07579064, -0.07157712, -0.07370815, 
    -0.06982328, -0.07094045, -0.06773105, -0.0693077, -0.06624616, 
    -0.06498045, -0.06381272, -0.06247527, -0.07477803, -0.0752454, 
    -0.0744108, -0.07327171, -0.07223132, -0.07087176, -0.07073423, 
    -0.07048298, -0.06983662, -0.06929789, -0.07040363, -0.06916353, 
    -0.0739392, -0.07139524, -0.07542279, -0.07418559, -0.0733384, 
    -0.0737089, -0.07180616, -0.07136515, -0.06960183, -0.07050768, 
    -0.06529039, -0.06754718, -0.06147688, -0.06311359, -0.07540938, 
    -0.07477969, -0.07263025, -0.07364484, -0.07078201, -0.0700952, 
    -0.06954208, -0.06884147, -0.06876635, -0.0683552, -0.06903028, 
    -0.06838176, -0.07086889, -0.06974602, -0.07287277, -0.07209849, 
    -0.07245366, -0.07284526, -0.07164369, -0.07038605, -0.0703596, 
    -0.06996135, -0.06885138, -0.07077065, -0.06500461, -0.06850478, 
    -0.07409925, -0.07291279, -0.07274515, -0.07320126, -0.07016374, 
    -0.07124888, -0.06836521, -0.0691324, -0.06788005, -0.06849937, 
    -0.06859098, -0.06939621, -0.06990246, -0.07119872, -0.0722719, 
    -0.07313494, -0.07293332, -0.07198858, -0.07030991, -0.06875947, 
    -0.06909601, -0.0679744, -0.07098564, -0.06970631, -0.07019785, 
    -0.06892371, -0.07174778, -0.069335, -0.07237836, -0.07210609, 
    -0.0712706, -0.0696203, -0.06926084, -0.06887887, -0.06911433, 
    -0.07026786, -0.07045882, -0.07129083, -0.07152226, -0.07216529, 
    -0.07270213, -0.07221143, -0.07169978, -0.07026744, -0.06900206, 
    -0.06764954, -0.06732284, -0.06578485, -0.0670338, -0.06498562, 
    -0.06672239, -0.06374598, -0.06919804, -0.06677451, -0.07123288, 
    -0.07073805, -0.06985194, -0.06786332, -0.06892965, -0.06768437, 
    -0.07046633, -0.07195613, -0.0723471, -0.07308214, -0.07233039, 
    -0.07239124, -0.07167879, -0.07190695, -0.0702204, -0.07112117, 
    -0.06859323, -0.06769416, -0.06522103, -0.06375159, -0.0622915, 
    -0.06165798, -0.0614665, -0.06138663,
  -0.08614824, -0.08423898, -0.08460681, -0.08309136, -0.08392866, 
    -0.08294123, -0.08575773, -0.084164, -0.08517796, -0.08597469, 
    -0.08022814, -0.08302442, -0.07742525, -0.07913453, -0.07491174, 
    -0.07768865, -0.07436416, -0.07499061, -0.07312158, -0.07365216, 
    -0.07131279, -0.07287802, -0.07013021, -0.07168356, -0.07143821, 
    -0.07293022, -0.08245404, -0.08057095, -0.08256695, -0.08229536, 
    -0.08241716, -0.08391121, -0.08467435, -0.08629609, -0.08599938, 
    -0.08480946, -0.08217353, -0.08305901, -0.08084605, -0.08089536, 
    -0.07850026, -0.07957114, -0.07565295, -0.07674628, -0.07362994, 
    -0.07440135, -0.07366596, -0.07388819, -0.07366307, -0.07479776, 
    -0.07430944, -0.07531591, -0.07936942, -0.07815563, -0.08183241, 
    -0.0841268, -0.08568716, -0.08681201, -0.08665208, -0.086348, 
    -0.08480255, -0.08337523, -0.08230381, -0.08159489, -0.08090246, 
    -0.07884208, -0.07777357, -0.0754337, -0.07585079, -0.07514571, 
    -0.07447854, -0.07337172, -0.07355276, -0.07306919, -0.07516434, 
    -0.07376516, -0.07608937, -0.07544637, -0.08071458, -0.08281921, 
    -0.08372995, -0.08453596, -0.08652931, -0.08514768, -0.08568963, 
    -0.08440614, -0.08360063, -0.08399807, -0.08157559, -0.08250884, 
    -0.0777107, -0.07974178, -0.07455605, -0.07576501, -0.07426922, 
    -0.07502873, -0.07373207, -0.07489803, -0.07289009, -0.07246009, 
    -0.07275365, -0.07163272, -0.07496319, -0.0736659, -0.0840092, 
    -0.08394424, -0.08364233, -0.08497768, -0.0850601, -0.0863042, 
    -0.08519637, -0.08472893, -0.08355423, -0.08286705, -0.08221915, 
    -0.08081265, -0.07927051, -0.07716412, -0.07568603, -0.07471132, 
    -0.07530752, -0.0747809, -0.07536982, -0.0756475, -0.07262086, 
    -0.07430486, -0.07179286, -0.0719296, -0.0730577, -0.07191418, 
    -0.08389866, -0.08427297, -0.0855855, -0.08455659, -0.08644081, 
    -0.08538084, -0.0847773, -0.08248908, -0.08199494, -0.08153921, 
    -0.08064682, -0.07951596, -0.0775708, -0.07591772, -0.07443994, 
    -0.07454723, -0.07450944, -0.07418295, -0.07499427, -0.07405061, 
    -0.07389336, -0.07430514, -0.07194793, -0.07261352, -0.07193251, 
    -0.0723651, -0.08415113, -0.08352323, -0.08386192, -0.08322614, 
    -0.08367349, -0.08170261, -0.08112092, -0.07845446, -0.07953803, 
    -0.07782076, -0.0793619, -0.07908655, -0.07776511, -0.07927787, 
    -0.07600781, -0.0782093, -0.07417028, -0.07631451, -0.07403796, 
    -0.07444627, -0.07377153, -0.07317243, -0.07242583, -0.07106831, 
    -0.07138037, -0.07026006, -0.08259602, -0.08179767, -0.08186778, 
    -0.08104005, -0.08043332, -0.07913418, -0.07709464, -0.07785531, 
    -0.07646476, -0.07618861, -0.07830358, -0.07699796, -0.08126785, 
    -0.08056194, -0.08098157, -0.08253268, -0.07767919, -0.08013271, 
    -0.07566182, -0.07694665, -0.07325753, -0.0750691, -0.07155272, 
    -0.07010064, -0.06876185, -0.06722955, -0.08136541, -0.0819041, 
    -0.08094221, -0.07963002, -0.07843213, -0.07686763, -0.07670942, 
    -0.07642043, -0.07567715, -0.07505782, -0.07632918, -0.07490338, 
    -0.08039887, -0.0774699, -0.08210858, -0.08068273, -0.07970682, 
    -0.08013356, -0.07794276, -0.07743527, -0.07540721, -0.07644885, 
    -0.07045613, -0.07304636, -0.06608647, -0.06796072, -0.08209313, 
    -0.08136731, -0.07889137, -0.08005978, -0.07676439, -0.07597449, 
    -0.07533853, -0.07453325, -0.07444692, -0.07397449, -0.07475024, 
    -0.07400502, -0.07686433, -0.07557299, -0.07917061, -0.07827923, 
    -0.07868807, -0.07913893, -0.07775579, -0.07630896, -0.07627854, 
    -0.07582057, -0.07454465, -0.07675132, -0.07012835, -0.07414637, 
    -0.08058326, -0.07921669, -0.07902367, -0.07954888, -0.0760533, 
    -0.07730149, -0.07398599, -0.07486761, -0.07342867, -0.07414015, 
    -0.0742454, -0.07517084, -0.07575286, -0.07724378, -0.07847883, 
    -0.07947251, -0.07924034, -0.07815272, -0.0762214, -0.07443902, 
    -0.07482579, -0.07353704, -0.07699863, -0.07552733, -0.07609252, 
    -0.07462776, -0.07787558, -0.07510048, -0.07860138, -0.07828797, 
    -0.07732648, -0.07542845, -0.07501523, -0.07457622, -0.07484685, 
    -0.07617304, -0.07639266, -0.07734975, -0.07761605, -0.07835611, 
    -0.07897414, -0.07840923, -0.07782035, -0.07617255, -0.07471781, 
    -0.0731639, -0.07278872, -0.07102337, -0.07245685, -0.07010657, 
    -0.07209934, -0.06868537, -0.07494306, -0.07215918, -0.07728308, 
    -0.07671383, -0.07569478, -0.07340945, -0.07463458, -0.07320391, 
    -0.07640129, -0.07811537, -0.07856541, -0.0794117, -0.07854617, 
    -0.07861622, -0.07779619, -0.07805876, -0.07611845, -0.07715455, 
    -0.074248, -0.07321515, -0.07037656, -0.06869179, -0.0670191, 
    -0.06629376, -0.06607459, -0.06598318,
  -0.06724861, -0.0657028, -0.06600061, -0.06477361, -0.06545154, 
    -0.06465206, -0.06693244, -0.0656421, -0.06646304, -0.06710809, 
    -0.06245529, -0.06471941, -0.0601857, -0.06156976, -0.05815042, 
    -0.06039899, -0.05770702, -0.05821428, -0.05670086, -0.05713048, 
    -0.05523624, -0.05650364, -0.05427869, -0.05553646, -0.05533779, 
    -0.05654591, -0.06425758, -0.06273286, -0.06434901, -0.06412911, 
    -0.06422772, -0.06543741, -0.0660553, -0.06736831, -0.06712808, 
    -0.06616469, -0.06403047, -0.06474742, -0.0629556, -0.06299553, 
    -0.06105618, -0.06192329, -0.0587506, -0.05963592, -0.05711249, 
    -0.05773713, -0.05714166, -0.05732161, -0.05713932, -0.05805812, 
    -0.05766271, -0.05847768, -0.06175996, -0.06077712, -0.06375425, 
    -0.06561197, -0.0668753, -0.06778599, -0.06765652, -0.06741033, 
    -0.06615909, -0.06500345, -0.06413595, -0.06356194, -0.06300128, 
    -0.06133296, -0.06046775, -0.05857307, -0.0589108, -0.05833987, 
    -0.05779964, -0.0569034, -0.05705, -0.05665844, -0.05835495, -0.05722198, 
    -0.05910399, -0.05858333, -0.06284916, -0.06455325, -0.06529065, 
    -0.06594324, -0.06755712, -0.06643853, -0.0668773, -0.06583814, 
    -0.06518595, -0.06550775, -0.06354631, -0.06430195, -0.06041684, 
    -0.06206146, -0.0578624, -0.05884134, -0.05763014, -0.05824515, 
    -0.05719519, -0.05813931, -0.05651341, -0.05616523, -0.05640293, 
    -0.05549529, -0.05819207, -0.05714162, -0.06551675, -0.06546416, 
    -0.06521972, -0.06630088, -0.06636762, -0.06737488, -0.06647795, 
    -0.06609949, -0.06514838, -0.06459199, -0.0640674, -0.06292856, 
    -0.06167986, -0.05997426, -0.05877739, -0.05798813, -0.05847089, 
    -0.05804447, -0.05852134, -0.05874619, -0.05629541, -0.057659, 
    -0.05562495, -0.05573568, -0.05664914, -0.05572319, -0.06542726, 
    -0.06573032, -0.066793, -0.06595995, -0.06748547, -0.0666273, 
    -0.06613865, -0.06428596, -0.06388586, -0.06351686, -0.06279428, 
    -0.06187861, -0.06030356, -0.058965, -0.05776838, -0.05785526, 
    -0.05782466, -0.05756028, -0.05821724, -0.05745313, -0.0573258, 
    -0.05765922, -0.05575052, -0.05628947, -0.05573804, -0.05608831, 
    -0.06563167, -0.06512328, -0.06539751, -0.06488274, -0.06524494, 
    -0.06364916, -0.06317817, -0.06101909, -0.06189648, -0.06050596, 
    -0.06175387, -0.0615309, -0.0604609, -0.06168583, -0.05903795, 
    -0.06082057, -0.05755003, -0.0592863, -0.05744288, -0.05777351, 
    -0.05722715, -0.05674203, -0.05613749, -0.05503828, -0.05529096, 
    -0.05438383, -0.06437255, -0.06372613, -0.06378289, -0.06311268, 
    -0.06262141, -0.06156947, -0.059918, -0.06053393, -0.05940795, 
    -0.05918435, -0.06089691, -0.05983971, -0.06329714, -0.06272556, 
    -0.06306534, -0.06432126, -0.06039132, -0.062378, -0.05875779, 
    -0.05979816, -0.05681094, -0.05827784, -0.05543052, -0.05425476, 
    -0.05317075, -0.05193013, -0.06337613, -0.0638123, -0.06303347, 
    -0.06197096, -0.061001, -0.05973418, -0.05960607, -0.05937206, 
    -0.0587702, -0.0582687, -0.05929817, -0.05814365, -0.06259353, 
    -0.06022185, -0.06397787, -0.06282336, -0.06203315, -0.0623787, 
    -0.06060475, -0.06019381, -0.05855162, -0.05939507, -0.0545426, 
    -0.05663995, -0.05100467, -0.05252212, -0.06396536, -0.06337767, 
    -0.06137287, -0.06231895, -0.05965058, -0.05901096, -0.058496, 
    -0.05784394, -0.05777403, -0.05739149, -0.05801964, -0.05741621, 
    -0.05973151, -0.05868585, -0.06159898, -0.0608772, -0.06120825, 
    -0.06157332, -0.06045335, -0.0592818, -0.05925717, -0.05888633, 
    -0.05785317, -0.05964, -0.05427719, -0.05753067, -0.06274281, 
    -0.06163629, -0.06147999, -0.06190527, -0.05907478, -0.06008549, 
    -0.0574008, -0.05811468, -0.05694951, -0.05752563, -0.05761085, 
    -0.05836022, -0.0588315, -0.06003875, -0.06103882, -0.06184343, 
    -0.06165544, -0.06077475, -0.0592109, -0.05776764, -0.05808081, 
    -0.05703726, -0.05984025, -0.05864888, -0.05910654, -0.05792047, 
    -0.06055035, -0.05830326, -0.06113806, -0.06088427, -0.06010573, 
    -0.05856882, -0.05823422, -0.05787873, -0.05809787, -0.05917174, 
    -0.05934957, -0.06012457, -0.0603402, -0.06093945, -0.06143988, 
    -0.06098246, -0.06050562, -0.05917135, -0.05799339, -0.05673513, 
    -0.05643133, -0.0550019, -0.05616261, -0.05425956, -0.05587313, 
    -0.05310883, -0.05817578, -0.05592158, -0.06007058, -0.05960964, 
    -0.05878447, -0.05693395, -0.05792599, -0.05676753, -0.05935656, 
    -0.06074451, -0.06110892, -0.06179419, -0.06109335, -0.06115006, 
    -0.06048606, -0.06069868, -0.05912754, -0.05996651, -0.05761296, 
    -0.05677662, -0.05447817, -0.05311403, -0.05175973, -0.05117249, 
    -0.05099506, -0.05092105,
  -0.0638878, -0.06219571, -0.06252145, -0.06118011, -0.06192097, 
    -0.06104734, -0.06354146, -0.06212931, -0.06302749, -0.06373387, 
    -0.05865141, -0.0611209, -0.05618335, -0.05768754, -0.0539767, 
    -0.05641496, -0.05349683, -0.05404584, -0.05240909, -0.05287335, 
    -0.05082871, -0.05219607, -0.04979745, -0.05115236, -0.05093817, 
    -0.05224172, -0.06061661, -0.05895377, -0.06071642, -0.06047637, 
    -0.06058401, -0.06190552, -0.06258129, -0.06401896, -0.06375577, 
    -0.06270097, -0.06036871, -0.0611515, -0.05919648, -0.05924, -0.05712904, 
    -0.0580722, -0.05462674, -0.05558664, -0.0528539, -0.05352941, 
    -0.05288543, -0.05307997, -0.0528829, -0.05387678, -0.05344889, 
    -0.05433109, -0.05789446, -0.05682575, -0.06006733, -0.06209638, 
    -0.06347889, -0.06447678, -0.06433484, -0.06406501, -0.06269485, 
    -0.06143122, -0.06048384, -0.05985754, -0.05924626, -0.05742998, 
    -0.05648965, -0.05443441, -0.05480035, -0.05418183, -0.05359704, 
    -0.05262792, -0.05278635, -0.05236326, -0.05419816, -0.05297226, 
    -0.05500976, -0.05444552, -0.05908049, -0.06093944, -0.06174509, 
    -0.06245869, -0.06422589, -0.06300066, -0.06348107, -0.06234372, 
    -0.06163065, -0.06198241, -0.0598405, -0.06066505, -0.05643435, 
    -0.05822259, -0.05366496, -0.05472507, -0.05341366, -0.05407926, 
    -0.0529433, -0.05396467, -0.05220662, -0.0518307, -0.05208732, 
    -0.05110797, -0.0540218, -0.05288538, -0.06199227, -0.06193476, 
    -0.06166755, -0.06285001, -0.06292305, -0.06402616, -0.06304381, 
    -0.06262964, -0.06158959, -0.06098174, -0.06040902, -0.05916701, 
    -0.05780732, -0.0559538, -0.05465577, -0.05380102, -0.05432373, 
    -0.05386201, -0.05437837, -0.05462196, -0.05197123, -0.05344488, 
    -0.05124779, -0.05136721, -0.05235322, -0.05135375, -0.06189442, 
    -0.0622258, -0.06338875, -0.06247697, -0.06414735, -0.06320732, 
    -0.06267248, -0.06064758, -0.06021091, -0.05980838, -0.05902069, 
    -0.05802358, -0.05631132, -0.05485909, -0.05356322, -0.05365723, 
    -0.05362411, -0.0533381, -0.05404904, -0.05322219, -0.0530845, 
    -0.05344512, -0.05138322, -0.05196482, -0.05136976, -0.05174769, 
    -0.06211792, -0.06156216, -0.0618619, -0.06129932, -0.06169512, 
    -0.05995268, -0.05943907, -0.05708873, -0.05804303, -0.05653114, 
    -0.05788784, -0.05764527, -0.0564822, -0.05781381, -0.05493817, 
    -0.05687296, -0.05332701, -0.05520742, -0.05321112, -0.05356877, 
    -0.05297784, -0.05245356, -0.05180077, -0.05061537, -0.05088769, 
    -0.0499106, -0.06074211, -0.06003665, -0.06009857, -0.05936769, 
    -0.05883235, -0.05768723, -0.05589274, -0.05656153, -0.05533936, 
    -0.05509688, -0.05695593, -0.05580777, -0.05956878, -0.05894582, 
    -0.05931609, -0.06068613, -0.05640663, -0.05856724, -0.05463453, 
    -0.05576269, -0.05252801, -0.05411466, -0.05103813, -0.04977169, 
    -0.04860622, -0.04727497, -0.05965491, -0.06013065, -0.05928135, 
    -0.0581241, -0.05706907, -0.05569325, -0.05555426, -0.05530043, 
    -0.05464798, -0.05410477, -0.0552203, -0.05396937, -0.05880198, 
    -0.0562226, -0.06031131, -0.05905238, -0.05819178, -0.05856799, 
    -0.05663846, -0.05619216, -0.05441117, -0.05532539, -0.05008151, 
    -0.05234329, -0.04628376, -0.04790984, -0.06029766, -0.05965659, 
    -0.05747338, -0.05850293, -0.05560255, -0.05490891, -0.05435093, 
    -0.05364498, -0.05356934, -0.05315554, -0.05383513, -0.05318227, 
    -0.05569036, -0.05455659, -0.05771932, -0.0569345, -0.05729437, 
    -0.05769141, -0.056474, -0.05520255, -0.05517584, -0.05477383, 
    -0.05365497, -0.05559107, -0.04979584, -0.05330606, -0.05896461, 
    -0.05775991, -0.05758988, -0.05805259, -0.05497809, -0.05607455, 
    -0.05316561, -0.05393801, -0.05267775, -0.05330061, -0.0533928, 
    -0.05420387, -0.05471441, -0.05602381, -0.05711018, -0.05798529, 
    -0.05778074, -0.05682318, -0.05512566, -0.05356242, -0.05390135, 
    -0.05277259, -0.05580836, -0.05451654, -0.05501252, -0.05372779, 
    -0.05657937, -0.05414218, -0.05721806, -0.05694219, -0.05609652, 
    -0.0544298, -0.05406743, -0.05368263, -0.05391981, -0.05508321, 
    -0.05527604, -0.05611697, -0.05635111, -0.05700216, -0.05754626, 
    -0.05704891, -0.05653078, -0.05508278, -0.05380671, -0.05244611, 
    -0.05211799, -0.05057618, -0.05182788, -0.04977685, -0.05151549, 
    -0.04853971, -0.05400416, -0.05156777, -0.05605836, -0.05555813, 
    -0.05466345, -0.05266094, -0.05373377, -0.05248111, -0.05528362, 
    -0.05679032, -0.05718638, -0.05793171, -0.05716945, -0.05723111, 
    -0.05650954, -0.05674052, -0.05503529, -0.05594539, -0.05339507, 
    -0.05249094, -0.05001215, -0.04854529, -0.04709235, -0.04646339, 
    -0.04627347, -0.04619428,
  -0.04035017, -0.03907184, -0.03931778, -0.03830553, -0.03886447, 
    -0.0382054, -0.04008836, -0.03902173, -0.03969999, -0.0402338, 
    -0.03640078, -0.03826088, -0.03454657, -0.03567605, -0.0328932, 
    -0.03472036, -0.03253425, -0.03294493, -0.03172141, -0.03206819, 
    -0.03054259, -0.03156237, -0.0297748, -0.03078379, -0.03062415, 
    -0.03159644, -0.03788066, -0.03662828, -0.0379559, -0.03777496, 
    -0.03785609, -0.03885281, -0.03936297, -0.04044933, -0.04025035, 
    -0.03945336, -0.03769382, -0.03828395, -0.03681095, -0.03684371, 
    -0.03525646, -0.03596519, -0.0333798, -0.03409905, -0.03205366, 
    -0.03255861, -0.03207722, -0.0322226, -0.03207533, -0.03281844, 
    -0.0324984, -0.03315843, -0.03583157, -0.0350287, -0.03746673, 
    -0.03899687, -0.04004107, -0.04079557, -0.04068821, -0.04048416, 
    -0.03944873, -0.03849493, -0.03778059, -0.03730871, -0.03684842, 
    -0.03548251, -0.03477641, -0.03323578, -0.03350982, -0.03304671, 
    -0.03260919, -0.03188484, -0.03200319, -0.03168719, -0.03305893, 
    -0.03214211, -0.03366669, -0.0332441, -0.03672365, -0.03812404, 
    -0.03873174, -0.0392704, -0.04060581, -0.03967972, -0.04004272, 
    -0.03918359, -0.03864539, -0.03891084, -0.03729587, -0.03791717, 
    -0.03473491, -0.03607827, -0.03265998, -0.03345343, -0.03247205, 
    -0.03296995, -0.03212046, -0.0328842, -0.03157025, -0.03128969, 
    -0.03148119, -0.0307507, -0.03292695, -0.03207719, -0.03891828, 
    -0.03887488, -0.03867324, -0.03956592, -0.0396211, -0.04045478, 
    -0.03971232, -0.03939948, -0.03861441, -0.03815594, -0.0377242, 
    -0.03678877, -0.03576607, -0.03437437, -0.03340153, -0.03276176, 
    -0.03315292, -0.03280739, -0.03319383, -0.03337621, -0.03139455, 
    -0.0324954, -0.03085493, -0.03094397, -0.03167969, -0.03093393, 
    -0.03884443, -0.03909456, -0.03997295, -0.03928419, -0.04054642, 
    -0.03983586, -0.03943183, -0.03790401, -0.03757491, -0.03727167, 
    -0.03667865, -0.03592864, -0.03464259, -0.03355382, -0.03258389, 
    -0.0326542, -0.03262943, -0.03241555, -0.03294734, -0.03232891, 
    -0.03222599, -0.03249558, -0.03095591, -0.03138977, -0.03094587, 
    -0.03122775, -0.03901313, -0.03859372, -0.03881989, -0.03839545, 
    -0.03869404, -0.03738037, -0.03699358, -0.03522618, -0.03594326, 
    -0.03480756, -0.03582659, -0.03564429, -0.03477082, -0.03577095, 
    -0.03361305, -0.03506416, -0.03240727, -0.0338148, -0.03232063, 
    -0.03258804, -0.03214628, -0.03175462, -0.03126735, -0.03038366, 
    -0.03058653, -0.02985898, -0.03797527, -0.03744363, -0.03749027, 
    -0.03693983, -0.03653692, -0.03567582, -0.03432857, -0.03483037, 
    -0.03391368, -0.03373196, -0.03512646, -0.03426485, -0.03709124, 
    -0.0366223, -0.03690099, -0.03793306, -0.03471411, -0.03633747, 
    -0.03338563, -0.03423104, -0.03181022, -0.03299643, -0.03069865, 
    -0.02975564, -0.0288894, -0.02790193, -0.03715609, -0.03751444, 
    -0.03687483, -0.0360042, -0.03521141, -0.03417898, -0.03407476, 
    -0.0338845, -0.0333957, -0.03298903, -0.03382445, -0.03288772, 
    -0.03651407, -0.03457602, -0.03765057, -0.0367025, -0.0360551, 
    -0.03633804, -0.03488811, -0.03455318, -0.03321838, -0.03390321, 
    -0.02998617, -0.03167228, -0.02716813, -0.02837259, -0.03764028, 
    -0.03715736, -0.03551513, -0.0362891, -0.03411097, -0.03359114, 
    -0.03317328, -0.03264504, -0.03258847, -0.03227909, -0.03278728, 
    -0.03229907, -0.03417681, -0.03332726, -0.03569993, -0.03511037, 
    -0.03538064, -0.03567896, -0.03476467, -0.03381115, -0.03379113, 
    -0.03348995, -0.03265251, -0.03410237, -0.0297736, -0.03239161, 
    -0.03663645, -0.03573044, -0.03560267, -0.03595044, -0.03364296, 
    -0.03446495, -0.03228661, -0.03286425, -0.03192206, -0.03238753, 
    -0.03245645, -0.0330632, -0.03344545, -0.03442689, -0.03524229, 
    -0.03589985, -0.03574609, -0.03502678, -0.03375353, -0.03258329, 
    -0.03283682, -0.03199291, -0.03426529, -0.03329727, -0.03366876, 
    -0.03270698, -0.03484375, -0.03301704, -0.03532331, -0.03511614, 
    -0.03448142, -0.03323233, -0.03296109, -0.0326732, -0.03285063, 
    -0.03372172, -0.03386622, -0.03449677, -0.03467245, -0.03516117, 
    -0.03556988, -0.03519628, -0.03480728, -0.0337214, -0.03276602, 
    -0.03174906, -0.03150408, -0.03035447, -0.03128758, -0.02975948, 
    -0.03105455, -0.02884002, -0.03291374, -0.03109354, -0.0344528, 
    -0.03407767, -0.03340728, -0.03190951, -0.03271146, -0.0317752, 
    -0.0338719, -0.0350021, -0.03529953, -0.03585957, -0.03528681, 
    -0.03533312, -0.03479134, -0.03496472, -0.03368582, -0.03436807, 
    -0.03245816, -0.03178254, -0.02993454, -0.02884416, -0.02776664, 
    -0.02730101, -0.02716052, -0.02710195,
  -0.01970495, -0.01870051, -0.01889313, -0.01810233, -0.01853834, 
    -0.01802441, -0.01949858, -0.0186613, -0.01919307, -0.01961318, 
    -0.01662921, -0.01806758, -0.01521542, -0.01607413, -0.01397334, 
    -0.01534703, -0.01370616, -0.01401192, -0.01310461, -0.01336065, 
    -0.01224113, -0.01298748, -0.01168475, -0.01241691, -0.01230052, 
    -0.01301256, -0.01777202, -0.01680408, -0.01783044, -0.01768999, 
    -0.01775294, -0.01852923, -0.01892854, -0.0197832, -0.01962623, 
    -0.01899943, -0.01762706, -0.01808554, -0.01694472, -0.01696996, 
    -0.0157542, -0.01629521, -0.01433697, -0.01487742, -0.01334991, 
    -0.01372426, -0.01336733, -0.01347495, -0.01336593, -0.01391762, 
    -0.01367953, -0.01417134, -0.01619298, -0.015581, -0.01745114, 
    -0.01864185, -0.01946134, -0.02005678, -0.01997189, -0.01981069, 
    -0.0189958, -0.0182499, -0.01769435, -0.01732889, -0.01697359, 
    -0.01592643, -0.01538952, -0.01422918, -0.01443441, -0.01408788, 
    -0.01376187, -0.01322516, -0.01331259, -0.01307939, -0.01409701, 
    -0.01341534, -0.01455213, -0.0142354, -0.01687748, -0.01796112, 
    -0.01843466, -0.01885599, -0.01990677, -0.01917714, -0.01946264, 
    -0.01878799, -0.01836725, -0.01857458, -0.01731896, -0.01780037, 
    -0.01535806, -0.0163818, -0.01379965, -0.01439214, -0.01365996, 
    -0.01403058, -0.01339933, -0.01396663, -0.01299328, -0.01278711, 
    -0.01292777, -0.01239277, -0.0139985, -0.0133673, -0.0185804, 
    -0.01854647, -0.01838898, -0.01908777, -0.01913109, -0.0197875, 
    -0.01920275, -0.01895718, -0.01834308, -0.01798592, -0.01765062, 
    -0.01692763, -0.01614291, -0.01508521, -0.01435325, -0.0138754, 
    -0.01416722, -0.01390938, -0.0141978, -0.01433429, -0.0128641, 
    -0.0136773, -0.01246885, -0.01253391, -0.01307387, -0.01252657, 
    -0.01852268, -0.01871829, -0.01940772, -0.0188668, -0.01985986, 
    -0.01929986, -0.01898255, -0.01779014, -0.01753491, -0.01730026, 
    -0.01684284, -0.01626723, -0.01528811, -0.01446741, -0.01374306, 
    -0.01379535, -0.01377692, -0.01361802, -0.01401371, -0.01355374, 
    -0.01347746, -0.01367744, -0.01254264, -0.01286059, -0.0125353, 
    -0.01274168, -0.01865457, -0.01832693, -0.0185035, -0.01817236, 
    -0.01840522, -0.01738431, -0.01708551, -0.01573116, -0.01627842, 
    -0.01541313, -0.01618917, -0.01604987, -0.01538528, -0.01614663, 
    -0.01451186, -0.01560794, -0.01361187, -0.01466342, -0.0135476, 
    -0.01374614, -0.01341843, -0.01312909, -0.01277073, -0.01212556, 
    -0.01227312, -0.01174552, -0.01784549, -0.01743325, -0.01746936, 
    -0.01704405, -0.01673382, -0.01607395, -0.01505061, -0.01543043, 
    -0.0147378, -0.01460116, -0.0156553, -0.0150025, -0.01716087, 
    -0.01679948, -0.0170141, -0.0178127, -0.01534229, -0.01658059, 
    -0.01434134, -0.01497698, -0.0131701, -0.01405035, -0.01235481, 
    -0.01167093, -0.01104941, -0.0103492, -0.01721095, -0.01748808, 
    -0.01699394, -0.01632508, -0.01571992, -0.0149377, -0.01485912, 
    -0.01471585, -0.01434888, -0.01404482, -0.01467068, -0.01396925, 
    -0.01671625, -0.01523771, -0.01759354, -0.01686119, -0.01636406, 
    -0.01658102, -0.01547424, -0.01522042, -0.01421617, -0.01472993, 
    -0.01183743, -0.0130684, -0.009834953, -0.01068181, -0.01758556, 
    -0.01721193, -0.0159513, -0.01654346, -0.01488641, -0.01449541, 
    -0.01418244, -0.01378853, -0.01374646, -0.0135168, -0.01389441, 
    -0.01353161, -0.01493606, -0.01429764, -0.01609237, -0.01564306, 
    -0.01584878, -0.01607635, -0.01538061, -0.01466068, -0.01464562, 
    -0.01441952, -0.01379409, -0.01487992, -0.01168389, -0.01360025, 
    -0.01681037, -0.01611568, -0.0160181, -0.01628392, -0.01453431, 
    -0.01515368, -0.01352238, -0.01395176, -0.01325265, -0.01359722, 
    -0.01364838, -0.0141002, -0.01438616, -0.0151249, -0.01574342, 
    -0.01624521, -0.01612764, -0.01557954, -0.01461737, -0.01374261, 
    -0.01393131, -0.01330499, -0.01500283, -0.01427519, -0.01455368, 
    -0.01383462, -0.01544059, -0.01406572, -0.01580511, -0.01564746, 
    -0.01516614, -0.0142266, -0.01402398, -0.01380948, -0.01394161, 
    -0.01459346, -0.0147021, -0.01517775, -0.01531073, -0.0156817, 
    -0.01599308, -0.01570841, -0.01541293, -0.01459322, -0.01387857, 
    -0.01312499, -0.0129446, -0.01210436, -0.01278557, -0.0116737, 
    -0.0126148, -0.01101418, -0.01398866, -0.01264334, -0.0151445, 
    -0.01486131, -0.01435756, -0.01324338, -0.01383795, -0.01314426, 
    -0.01470637, -0.01556079, -0.01578699, -0.0162144, -0.01577731, 
    -0.01581258, -0.01540083, -0.0155324, -0.01456649, -0.01508045, 
    -0.01364964, -0.01314967, -0.01180011, -0.01101713, -0.01025399, 
    -0.009927681, -0.009829647, -0.009788836,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  363.612, 365.4624, 365.1021, 366.5885, 365.7677, 366.7354, 363.9866, 
    365.5361, 364.5464, 363.7782, 369.4446, 366.654, 372.3569, 370.5666, 
    375.0744, 372.0781, 375.6804, 374.9874, 377.0748, 376.476, 379.1507, 
    377.3513, 380.5399, 378.7206, 379.0049, 377.292, 367.2142, 369.0965, 
    367.1029, 367.3709, 367.2506, 365.7849, 365.0363, 363.4707, 363.7545, 
    364.9045, 367.4914, 366.6201, 368.8181, 368.7684, 371.2256, 370.1164, 
    374.2621, 373.0807, 376.501, 375.639, 376.4605, 376.2112, 376.4638, 
    375.2, 375.7411, 374.6303, 370.324, 371.5863, 367.83, 365.5727, 364.0545, 
    362.9798, 363.1316, 363.4212, 364.9112, 366.3096, 367.3625, 368.0666, 
    368.7613, 370.8698, 371.9884, 374.5014, 374.0469, 374.817, 375.5533, 
    376.7919, 376.5878, 377.1342, 374.7964, 376.3492, 373.7881, 374.4875, 
    368.9512, 366.855, 365.9625, 365.1714, 363.2484, 364.5757, 364.0521, 
    365.2984, 366.0888, 365.6993, 368.0859, 367.1602, 372.0548, 369.9413, 
    375.4673, 374.1401, 375.7859, 374.9455, 376.3863, 375.0894, 377.3376, 
    377.828, 377.493, 378.7793, 375.0176, 376.4606, 365.6883, 365.7523, 
    366.048, 364.7408, 364.6607, 363.463, 364.5285, 364.9829, 366.1342, 
    366.808, 367.4462, 368.8519, 370.4261, 372.6344, 374.2261, 375.2955, 
    374.6394, 375.2186, 374.5712, 374.268, 377.6446, 375.7463, 378.5942, 
    378.4365, 377.1473, 378.4543, 365.7973, 365.429, 364.1524, 365.1512, 
    363.3327, 364.35, 364.9358, 367.1797, 367.6684, 368.1223, 369.0195, 
    370.1731, 372.2027, 373.9742, 375.5961, 375.4771, 375.519, 375.882, 
    374.9834, 376.0296, 376.2055, 375.7459, 378.4154, 377.6529, 378.4332, 
    377.9366, 365.5486, 366.1646, 365.8335, 366.4561, 366.0176, 367.9593, 
    368.5415, 371.2735, 370.1505, 371.9386, 370.3318, 370.6162, 371.9974, 
    370.4184, 373.8766, 371.5302, 375.8961, 373.5451, 376.0438, 375.5891, 
    376.342, 377.0172, 377.8671, 379.4357, 379.0721, 380.386, 367.0743, 
    367.8645, 367.7947, 368.6227, 369.2359, 370.5669, 372.7084, 371.9021, 
    373.383, 373.6808, 371.4312, 372.8116, 368.3939, 369.1055, 368.6816, 
    367.1367, 372.0881, 369.5417, 374.2524, 372.8663, 376.9209, 374.9012, 
    378.872, 380.5751, 382.1815, 384.0653, 368.2961, 367.7586, 368.7212, 
    370.056, 371.2968, 372.9508, 373.1202, 373.4308, 374.2357, 374.9135, 
    373.5292, 375.0835, 369.271, 372.3095, 367.5557, 368.9832, 369.9771, 
    369.5408, 371.81, 372.3462, 374.5304, 373.4001, 380.1544, 377.1602, 
    385.503, 383.1603, 367.571, 368.2942, 370.8185, 369.616, 373.0613, 
    373.9126, 374.6055, 375.4926, 375.5884, 376.1147, 375.2525, 376.0806, 
    372.9543, 374.3493, 370.5292, 371.4568, 371.0298, 370.562, 372.0071, 
    373.551, 373.5837, 374.0797, 375.4803, 373.0753, 380.5424, 375.923, 
    369.0838, 370.4817, 370.6813, 370.1393, 373.8272, 372.4883, 376.1018, 
    375.1229, 376.7276, 375.9297, 375.8124, 374.7893, 374.1533, 372.5496, 
    371.248, 370.2178, 370.4572, 371.5894, 373.6455, 375.5972, 375.1691, 
    376.6055, 372.8108, 374.3991, 373.7848, 375.3879, 371.8808, 374.8669, 
    371.1201, 371.4476, 372.4617, 374.5072, 374.9603, 375.445, 375.1458, 
    373.6977, 373.4607, 372.437, 372.1548, 371.3762, 370.7326, 371.3207, 
    371.939, 373.6982, 375.2884, 377.0269, 377.453, 379.4883, 377.8318, 
    380.5683, 378.2416, 382.2747, 375.0399, 378.1727, 372.5078, 373.1155, 
    374.2166, 376.7494, 375.3804, 376.9817, 373.4514, 371.6286, 371.1576, 
    370.2804, 371.1777, 371.1046, 371.9644, 371.688, 373.7567, 372.6445, 
    375.8095, 376.9689, 380.2483, 382.2667, 384.3278, 385.2401, 385.5181, 
    385.6343 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.190983e-08, 6.218286e-08, 6.212978e-08, 6.234999e-08, 6.222784e-08, 
    6.237203e-08, 6.196519e-08, 6.219368e-08, 6.204782e-08, 6.193441e-08, 
    6.277735e-08, 6.235982e-08, 6.321117e-08, 6.294484e-08, 6.361391e-08, 
    6.316971e-08, 6.370349e-08, 6.360111e-08, 6.390928e-08, 6.382099e-08, 
    6.421514e-08, 6.395003e-08, 6.44195e-08, 6.415184e-08, 6.41937e-08, 
    6.394128e-08, 6.244386e-08, 6.272536e-08, 6.242718e-08, 6.246731e-08, 
    6.244931e-08, 6.223036e-08, 6.212002e-08, 6.188898e-08, 6.193092e-08, 
    6.210062e-08, 6.248537e-08, 6.235477e-08, 6.268395e-08, 6.267651e-08, 
    6.3043e-08, 6.287775e-08, 6.349378e-08, 6.331869e-08, 6.382468e-08, 
    6.369742e-08, 6.38187e-08, 6.378193e-08, 6.381918e-08, 6.363254e-08, 
    6.371251e-08, 6.354828e-08, 6.29087e-08, 6.309665e-08, 6.253609e-08, 
    6.219904e-08, 6.197521e-08, 6.181637e-08, 6.183883e-08, 6.188163e-08, 
    6.210161e-08, 6.230846e-08, 6.246609e-08, 6.257154e-08, 6.267544e-08, 
    6.298992e-08, 6.315641e-08, 6.352918e-08, 6.346192e-08, 6.357588e-08, 
    6.368477e-08, 6.386757e-08, 6.383748e-08, 6.391802e-08, 6.357288e-08, 
    6.380225e-08, 6.34236e-08, 6.352716e-08, 6.270364e-08, 6.239001e-08, 
    6.225666e-08, 6.213998e-08, 6.185609e-08, 6.205214e-08, 6.197485e-08, 
    6.215873e-08, 6.227556e-08, 6.221778e-08, 6.257442e-08, 6.243577e-08, 
    6.316627e-08, 6.28516e-08, 6.367206e-08, 6.347572e-08, 6.371913e-08, 
    6.359492e-08, 6.380773e-08, 6.361621e-08, 6.394799e-08, 6.402023e-08, 
    6.397087e-08, 6.416053e-08, 6.360559e-08, 6.38187e-08, 6.221616e-08, 
    6.222558e-08, 6.226949e-08, 6.207648e-08, 6.206467e-08, 6.188782e-08, 
    6.204519e-08, 6.21122e-08, 6.228234e-08, 6.238297e-08, 6.247863e-08, 
    6.268897e-08, 6.292388e-08, 6.325241e-08, 6.348845e-08, 6.364667e-08, 
    6.354966e-08, 6.363531e-08, 6.353956e-08, 6.349468e-08, 6.399316e-08, 
    6.371325e-08, 6.413325e-08, 6.411001e-08, 6.391993e-08, 6.411263e-08, 
    6.22322e-08, 6.217797e-08, 6.198967e-08, 6.213703e-08, 6.186856e-08, 
    6.201883e-08, 6.210523e-08, 6.243865e-08, 6.251192e-08, 6.257985e-08, 
    6.271402e-08, 6.288621e-08, 6.318828e-08, 6.345113e-08, 6.36911e-08, 
    6.367352e-08, 6.367971e-08, 6.373331e-08, 6.360052e-08, 6.375511e-08, 
    6.378105e-08, 6.371322e-08, 6.41069e-08, 6.399443e-08, 6.410952e-08, 
    6.403629e-08, 6.21956e-08, 6.228685e-08, 6.223754e-08, 6.233027e-08, 
    6.226494e-08, 6.255542e-08, 6.264251e-08, 6.305007e-08, 6.288282e-08, 
    6.314902e-08, 6.290986e-08, 6.295224e-08, 6.315769e-08, 6.292279e-08, 
    6.343662e-08, 6.308824e-08, 6.373539e-08, 6.338745e-08, 6.37572e-08, 
    6.369006e-08, 6.380122e-08, 6.390078e-08, 6.402603e-08, 6.425714e-08, 
    6.420363e-08, 6.439692e-08, 6.24229e-08, 6.254125e-08, 6.253084e-08, 
    6.265472e-08, 6.274633e-08, 6.294491e-08, 6.326341e-08, 6.314364e-08, 
    6.336354e-08, 6.340768e-08, 6.307361e-08, 6.327871e-08, 6.262048e-08, 
    6.272681e-08, 6.266351e-08, 6.243223e-08, 6.317123e-08, 6.279195e-08, 
    6.349235e-08, 6.328687e-08, 6.388658e-08, 6.358832e-08, 6.417417e-08, 
    6.442461e-08, 6.466037e-08, 6.493585e-08, 6.260586e-08, 6.252544e-08, 
    6.266945e-08, 6.286869e-08, 6.305359e-08, 6.32994e-08, 6.332456e-08, 
    6.33706e-08, 6.348989e-08, 6.359019e-08, 6.338515e-08, 6.361533e-08, 
    6.275145e-08, 6.320415e-08, 6.249503e-08, 6.270854e-08, 6.285696e-08, 
    6.279186e-08, 6.312996e-08, 6.320965e-08, 6.353348e-08, 6.336608e-08, 
    6.436279e-08, 6.39218e-08, 6.514564e-08, 6.480359e-08, 6.249734e-08, 
    6.260559e-08, 6.298236e-08, 6.28031e-08, 6.331581e-08, 6.344202e-08, 
    6.354463e-08, 6.367578e-08, 6.368995e-08, 6.376766e-08, 6.364031e-08, 
    6.376263e-08, 6.329992e-08, 6.35067e-08, 6.293931e-08, 6.307739e-08, 
    6.301387e-08, 6.294419e-08, 6.315926e-08, 6.338838e-08, 6.339329e-08, 
    6.346676e-08, 6.367377e-08, 6.331789e-08, 6.441968e-08, 6.373919e-08, 
    6.272364e-08, 6.293214e-08, 6.296194e-08, 6.288117e-08, 6.342937e-08, 
    6.323073e-08, 6.376577e-08, 6.362117e-08, 6.38581e-08, 6.374036e-08, 
    6.372304e-08, 6.357183e-08, 6.347768e-08, 6.323983e-08, 6.304632e-08, 
    6.289289e-08, 6.292857e-08, 6.309711e-08, 6.34024e-08, 6.369122e-08, 
    6.362795e-08, 6.384009e-08, 6.327863e-08, 6.351405e-08, 6.342306e-08, 
    6.366032e-08, 6.314046e-08, 6.358311e-08, 6.302731e-08, 6.307604e-08, 
    6.322679e-08, 6.353001e-08, 6.359712e-08, 6.366874e-08, 6.362455e-08, 
    6.341015e-08, 6.337503e-08, 6.322313e-08, 6.318118e-08, 6.306544e-08, 
    6.296961e-08, 6.305716e-08, 6.31491e-08, 6.341025e-08, 6.364559e-08, 
    6.390219e-08, 6.3965e-08, 6.426479e-08, 6.402072e-08, 6.442347e-08, 
    6.408103e-08, 6.467384e-08, 6.360878e-08, 6.407099e-08, 6.323365e-08, 
    6.332385e-08, 6.3487e-08, 6.386124e-08, 6.365921e-08, 6.389548e-08, 
    6.337365e-08, 6.310292e-08, 6.303289e-08, 6.290222e-08, 6.303588e-08, 
    6.302501e-08, 6.315292e-08, 6.311182e-08, 6.341892e-08, 6.325396e-08, 
    6.37226e-08, 6.389362e-08, 6.437666e-08, 6.467278e-08, 6.497426e-08, 
    6.510736e-08, 6.514787e-08, 6.516481e-08 ;

 SOM_C_LEACHED =
  1.901379e-20, 7.966147e-20, 3.717541e-20, 3.391367e-21, -5.970066e-20, 
    -6.803741e-20, -6.361204e-21, 5.21695e-20, 3.274475e-21, -4.359097e-21, 
    -3.803636e-20, -8.197168e-20, -2.896278e-20, 3.437594e-20, 6.121997e-20, 
    -6.119233e-20, -9.231051e-21, -2.104595e-20, 2.451709e-20, 1.044391e-21, 
    -3.181237e-20, 5.529554e-20, -4.32328e-20, -3.744575e-20, -2.381505e-20, 
    -8.713728e-21, -5.640072e-20, 1.3618e-21, -2.560845e-20, 4.02167e-21, 
    2.534358e-20, 1.74214e-20, -1.587115e-20, 1.671824e-20, 3.015938e-20, 
    1.207607e-20, -7.382811e-20, -1.521761e-20, -2.675106e-20, -1.518307e-20, 
    -4.397901e-20, 2.444069e-20, -2.79059e-20, -5.114637e-21, 2.00387e-21, 
    -1.110592e-19, -5.662536e-20, 7.872418e-21, 7.723169e-21, -2.777038e-20, 
    -4.435189e-21, -2.686042e-20, 8.936775e-21, 1.605617e-20, -1.83772e-20, 
    -5.898651e-20, -2.289942e-20, 2.305124e-20, 2.512272e-20, 4.450246e-21, 
    3.471969e-20, -3.570283e-20, 1.939359e-20, 3.832378e-20, -2.106534e-21, 
    -5.694721e-20, 3.192324e-20, -3.446372e-20, 7.697484e-20, -4.208612e-20, 
    -2.962246e-20, 1.615009e-20, -3.939531e-20, 1.259805e-20, -1.048774e-20, 
    3.86832e-20, 5.260086e-21, 7.615705e-20, -8.557702e-21, -4.690645e-20, 
    -6.286806e-20, -2.128973e-21, 1.945636e-22, -4.347333e-20, 5.384927e-20, 
    -3.179942e-20, 3.457576e-20, -3.12483e-20, 9.45383e-20, -9.584202e-21, 
    4.559086e-21, 2.367859e-21, 2.481093e-20, -4.921299e-20, 1.29007e-20, 
    -4.028188e-20, 6.543742e-21, 7.259442e-20, 2.552523e-21, 1.562173e-21, 
    2.285965e-20, -3.804616e-21, -4.433078e-20, 1.643117e-20, -3.220197e-20, 
    3.355215e-20, 3.576174e-20, 5.700768e-20, 1.921264e-20, -2.154986e-20, 
    6.530911e-20, -1.508543e-20, -2.423926e-21, 1.150309e-20, 3.256609e-20, 
    -1.194721e-20, -4.604023e-20, -3.446768e-20, 1.316625e-20, -1.797865e-20, 
    -3.810864e-20, -1.820253e-21, -4.167427e-20, -2.983773e-20, 
    -1.197799e-20, -2.441213e-21, -3.83313e-20, -5.061652e-20, 1.362604e-20, 
    -1.275621e-20, -2.026118e-20, -4.759978e-20, 3.116482e-20, 1.059783e-20, 
    -8.248343e-21, 2.612406e-20, -1.988515e-20, 1.000714e-20, -1.773569e-20, 
    -9.192375e-21, 3.820041e-20, 4.849014e-20, -3.00039e-20, 6.297912e-21, 
    2.209561e-20, 1.256283e-20, -9.264347e-20, -3.140321e-20, -5.697092e-21, 
    -7.118776e-20, -2.988995e-20, 3.643055e-20, -1.072051e-20, -8.996137e-20, 
    -1.412978e-20, 3.92262e-20, -1.061223e-20, 4.38921e-20, 2.72497e-20, 
    2.624065e-21, -5.964228e-20, -4.253225e-20, -1.414599e-20, -6.447274e-20, 
    -1.181452e-20, -2.376276e-20, -1.972536e-21, 8.192234e-21, -2.392836e-20, 
    9.384974e-21, 2.427931e-20, -4.733808e-20, 8.827981e-21, 3.351072e-20, 
    -3.468338e-20, 3.33042e-20, -4.368846e-20, 3.733225e-20, -2.260004e-20, 
    -4.827802e-20, -2.086899e-21, 1.16985e-20, 2.974612e-20, 6.493208e-21, 
    -6.840384e-20, 3.318032e-20, 1.970923e-20, -4.330293e-20, 1.961912e-20, 
    -3.09563e-20, 5.946856e-20, -2.721978e-20, -9.844298e-21, 4.193037e-20, 
    3.595345e-21, -1.094588e-20, 2.177123e-20, -9.566509e-21, 2.502063e-20, 
    -5.866553e-20, 2.246528e-20, -2.05286e-20, -8.848903e-20, -1.278634e-20, 
    -4.065381e-20, 1.687646e-20, 1.290883e-20, 3.551526e-20, -5.777194e-20, 
    8.221464e-20, -3.2671e-20, -1.269456e-20, -5.567709e-21, -1.79081e-20, 
    3.157749e-20, 1.254514e-20, 5.223525e-21, -2.08403e-20, -1.919515e-20, 
    3.980347e-20, -1.056592e-20, -8.929504e-21, 3.029155e-20, -9.648795e-21, 
    6.259462e-20, 5.325014e-20, -3.703843e-20, 7.526246e-20, -1.4028e-20, 
    2.282261e-20, 3.958275e-20, 2.239166e-20, 3.227932e-20, -4.829831e-20, 
    -2.02462e-20, 4.45548e-20, -5.848754e-22, 1.753356e-20, 4.396805e-20, 
    1.475752e-20, 2.838967e-20, -1.143456e-20, 7.231228e-20, -1.631038e-20, 
    -1.314104e-20, -5.092829e-20, 6.15578e-20, -4.789485e-20, 4.15292e-21, 
    -2.17885e-20, -4.037203e-20, -5.453586e-20, 1.120172e-21, 1.06976e-20, 
    -7.625418e-21, 1.031273e-20, -8.976092e-21, -2.549064e-20, 7.068656e-20, 
    -2.119023e-20, -5.872666e-20, 2.411349e-20, 3.802481e-20, 3.9656e-20, 
    8.058171e-20, 6.538376e-21, 6.912861e-20, 1.322579e-21, -2.264342e-20, 
    -1.513401e-20, 5.722904e-20, 7.022605e-21, -6.29132e-20, -3.728482e-20, 
    -5.537131e-20, -2.986193e-20, -6.25852e-20, -1.936711e-20, -5.392956e-20, 
    3.884838e-20, -5.142991e-20, 2.495772e-20, -6.539166e-20, 3.090264e-20, 
    7.334605e-20, 5.89084e-20, -8.195965e-20, -1.721241e-20, -2.196552e-20, 
    -1.608081e-20, -2.878163e-20, -2.360907e-20, 2.676231e-21, -5.383244e-20, 
    -2.191138e-21, 4.043485e-20, 4.375235e-21, -3.427655e-20, -3.604844e-20, 
    -4.784653e-21, 5.818566e-20, 1.442349e-20, -4.387874e-21, -2.310855e-20, 
    6.611111e-20, -2.27952e-20, 3.082987e-20, 3.124934e-20, -4.320503e-20, 
    1.519638e-20, -8.036607e-20, -4.555636e-20, -2.563021e-21, -4.595284e-20, 
    -2.775955e-20, -4.176972e-21, 9.956745e-22, 2.6878e-21, 2.426667e-20, 
    2.264516e-20, -1.184436e-20, -3.103501e-20, 6.875593e-20, -3.800497e-21, 
    5.073869e-20, -8.63863e-20, -8.17246e-20, -5.156077e-20, 1.439384e-20, 
    -3.018139e-20, 8.131292e-21, 5.876923e-21, -4.619698e-21, 2.257825e-20, 
    -1.984811e-20, -4.914792e-20, -3.467586e-20, -3.011617e-20 ;

 SR =
  6.191079e-08, 6.218382e-08, 6.213074e-08, 6.235096e-08, 6.22288e-08, 
    6.2373e-08, 6.196615e-08, 6.219464e-08, 6.204878e-08, 6.193537e-08, 
    6.277832e-08, 6.236078e-08, 6.321213e-08, 6.294581e-08, 6.361488e-08, 
    6.317068e-08, 6.370446e-08, 6.360209e-08, 6.391026e-08, 6.382197e-08, 
    6.421612e-08, 6.395101e-08, 6.442048e-08, 6.415281e-08, 6.419468e-08, 
    6.394226e-08, 6.244482e-08, 6.272633e-08, 6.242814e-08, 6.246828e-08, 
    6.245027e-08, 6.223132e-08, 6.212098e-08, 6.188993e-08, 6.193188e-08, 
    6.210158e-08, 6.248633e-08, 6.235573e-08, 6.268491e-08, 6.267748e-08, 
    6.304396e-08, 6.287872e-08, 6.349475e-08, 6.331966e-08, 6.382565e-08, 
    6.369839e-08, 6.381968e-08, 6.378291e-08, 6.382015e-08, 6.363351e-08, 
    6.371348e-08, 6.354926e-08, 6.290966e-08, 6.309762e-08, 6.253705e-08, 
    6.219999e-08, 6.197617e-08, 6.181733e-08, 6.183978e-08, 6.188259e-08, 
    6.210257e-08, 6.230942e-08, 6.246706e-08, 6.25725e-08, 6.267641e-08, 
    6.299089e-08, 6.315737e-08, 6.353015e-08, 6.346289e-08, 6.357685e-08, 
    6.368574e-08, 6.386854e-08, 6.383846e-08, 6.391899e-08, 6.357385e-08, 
    6.380323e-08, 6.342457e-08, 6.352813e-08, 6.270461e-08, 6.239097e-08, 
    6.225762e-08, 6.214094e-08, 6.185705e-08, 6.20531e-08, 6.197581e-08, 
    6.215969e-08, 6.227652e-08, 6.221874e-08, 6.257539e-08, 6.243673e-08, 
    6.316724e-08, 6.285257e-08, 6.367303e-08, 6.34767e-08, 6.37201e-08, 
    6.35959e-08, 6.380871e-08, 6.361718e-08, 6.394897e-08, 6.402121e-08, 
    6.397185e-08, 6.416151e-08, 6.360656e-08, 6.381967e-08, 6.221712e-08, 
    6.222654e-08, 6.227045e-08, 6.207744e-08, 6.206563e-08, 6.188878e-08, 
    6.204615e-08, 6.211316e-08, 6.22833e-08, 6.238393e-08, 6.247959e-08, 
    6.268994e-08, 6.292485e-08, 6.325337e-08, 6.348942e-08, 6.364765e-08, 
    6.355063e-08, 6.363629e-08, 6.354053e-08, 6.349565e-08, 6.399414e-08, 
    6.371423e-08, 6.413423e-08, 6.411099e-08, 6.392091e-08, 6.411361e-08, 
    6.223316e-08, 6.217893e-08, 6.199063e-08, 6.213799e-08, 6.186952e-08, 
    6.201979e-08, 6.210619e-08, 6.243962e-08, 6.251289e-08, 6.258082e-08, 
    6.271499e-08, 6.288717e-08, 6.318925e-08, 6.34521e-08, 6.369208e-08, 
    6.367449e-08, 6.368068e-08, 6.373428e-08, 6.36015e-08, 6.375608e-08, 
    6.378202e-08, 6.37142e-08, 6.410788e-08, 6.39954e-08, 6.411049e-08, 
    6.403727e-08, 6.219656e-08, 6.228781e-08, 6.22385e-08, 6.233122e-08, 
    6.22659e-08, 6.255637e-08, 6.264347e-08, 6.305104e-08, 6.288379e-08, 
    6.315e-08, 6.291083e-08, 6.295321e-08, 6.315866e-08, 6.292376e-08, 
    6.34376e-08, 6.30892e-08, 6.373637e-08, 6.338842e-08, 6.375817e-08, 
    6.369104e-08, 6.38022e-08, 6.390175e-08, 6.402701e-08, 6.425812e-08, 
    6.420461e-08, 6.43979e-08, 6.242386e-08, 6.254222e-08, 6.253181e-08, 
    6.265568e-08, 6.27473e-08, 6.294588e-08, 6.326439e-08, 6.314462e-08, 
    6.336451e-08, 6.340865e-08, 6.307459e-08, 6.327969e-08, 6.262145e-08, 
    6.272778e-08, 6.266447e-08, 6.243319e-08, 6.31722e-08, 6.279292e-08, 
    6.349332e-08, 6.328784e-08, 6.388755e-08, 6.358929e-08, 6.417515e-08, 
    6.442559e-08, 6.466136e-08, 6.493683e-08, 6.260683e-08, 6.25264e-08, 
    6.267042e-08, 6.286966e-08, 6.305456e-08, 6.330037e-08, 6.332552e-08, 
    6.337157e-08, 6.349087e-08, 6.359117e-08, 6.338612e-08, 6.361631e-08, 
    6.275242e-08, 6.320513e-08, 6.249599e-08, 6.27095e-08, 6.285792e-08, 
    6.279282e-08, 6.313093e-08, 6.321061e-08, 6.353445e-08, 6.336705e-08, 
    6.436377e-08, 6.392277e-08, 6.514664e-08, 6.480458e-08, 6.24983e-08, 
    6.260656e-08, 6.298333e-08, 6.280406e-08, 6.331678e-08, 6.3443e-08, 
    6.354561e-08, 6.367676e-08, 6.369093e-08, 6.376864e-08, 6.364129e-08, 
    6.376361e-08, 6.33009e-08, 6.350767e-08, 6.294027e-08, 6.307836e-08, 
    6.301484e-08, 6.294515e-08, 6.316022e-08, 6.338935e-08, 6.339426e-08, 
    6.346773e-08, 6.367474e-08, 6.331886e-08, 6.442066e-08, 6.374017e-08, 
    6.272461e-08, 6.293312e-08, 6.296292e-08, 6.288214e-08, 6.343034e-08, 
    6.32317e-08, 6.376674e-08, 6.362214e-08, 6.385908e-08, 6.374134e-08, 
    6.372401e-08, 6.35728e-08, 6.347865e-08, 6.32408e-08, 6.30473e-08, 
    6.289386e-08, 6.292954e-08, 6.309808e-08, 6.340337e-08, 6.36922e-08, 
    6.362893e-08, 6.384107e-08, 6.327961e-08, 6.351502e-08, 6.342403e-08, 
    6.36613e-08, 6.314143e-08, 6.358408e-08, 6.302828e-08, 6.307702e-08, 
    6.322776e-08, 6.353098e-08, 6.359809e-08, 6.366972e-08, 6.362552e-08, 
    6.341112e-08, 6.337601e-08, 6.322409e-08, 6.318215e-08, 6.306641e-08, 
    6.297058e-08, 6.305813e-08, 6.315008e-08, 6.341122e-08, 6.364657e-08, 
    6.390317e-08, 6.396598e-08, 6.426577e-08, 6.402171e-08, 6.442445e-08, 
    6.408201e-08, 6.467483e-08, 6.360975e-08, 6.407196e-08, 6.323462e-08, 
    6.332483e-08, 6.348797e-08, 6.386221e-08, 6.366019e-08, 6.389647e-08, 
    6.337463e-08, 6.310389e-08, 6.303387e-08, 6.290318e-08, 6.303685e-08, 
    6.302598e-08, 6.315389e-08, 6.311279e-08, 6.341989e-08, 6.325493e-08, 
    6.372358e-08, 6.38946e-08, 6.437764e-08, 6.467376e-08, 6.497525e-08, 
    6.510835e-08, 6.514885e-08, 6.516579e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3396222, -0.3396269, -0.339626, -0.3396298, -0.3396277, -0.3396302, 
    -0.3396232, -0.3396271, -0.3396246, -0.3396227, -0.3396372, -0.33963, 
    -0.3396452, -0.3396405, -0.3396525, -0.3396444, -0.3396542, -0.3396524, 
    -0.339658, -0.3396564, -0.3396634, -0.3396588, -0.3396672, -0.3396624, 
    -0.3396631, -0.3396586, -0.3396315, -0.3396362, -0.3396312, -0.3396319, 
    -0.3396316, -0.3396277, -0.3396257, -0.3396219, -0.3396226, -0.3396255, 
    -0.3396322, -0.3396299, -0.3396358, -0.3396357, -0.3396423, -0.3396393, 
    -0.3396504, -0.3396473, -0.3396565, -0.3396541, -0.3396564, -0.3396557, 
    -0.3396564, -0.339653, -0.3396544, -0.3396514, -0.3396398, -0.3396432, 
    -0.3396331, -0.3396271, -0.3396233, -0.3396206, -0.339621, -0.3396217, 
    -0.3396255, -0.3396291, -0.3396319, -0.3396338, -0.3396356, -0.3396411, 
    -0.3396442, -0.339651, -0.3396499, -0.3396519, -0.3396539, -0.3396572, 
    -0.3396567, -0.3396581, -0.3396519, -0.339656, -0.3396492, -0.339651, 
    -0.3396358, -0.3396305, -0.3396281, -0.3396262, -0.3396213, -0.3396246, 
    -0.3396233, -0.3396266, -0.3396286, -0.3396276, -0.3396338, -0.3396313, 
    -0.3396444, -0.3396387, -0.3396537, -0.3396501, -0.3396546, -0.3396523, 
    -0.3396561, -0.3396527, -0.3396587, -0.33966, -0.3396591, -0.3396626, 
    -0.3396525, -0.3396563, -0.3396275, -0.3396277, -0.3396285, -0.3396251, 
    -0.3396249, -0.3396219, -0.3396246, -0.3396257, -0.3396287, -0.3396304, 
    -0.3396321, -0.3396358, -0.3396401, -0.339646, -0.3396503, -0.3396533, 
    -0.3396515, -0.339653, -0.3396513, -0.3396505, -0.3396595, -0.3396544, 
    -0.3396621, -0.3396617, -0.3396582, -0.3396617, -0.3396278, -0.3396269, 
    -0.3396236, -0.3396262, -0.3396215, -0.3396241, -0.3396255, -0.3396313, 
    -0.3396327, -0.3396339, -0.3396363, -0.3396394, -0.3396448, -0.3396496, 
    -0.3396541, -0.3396537, -0.3396538, -0.3396548, -0.3396524, -0.3396552, 
    -0.3396556, -0.3396544, -0.3396616, -0.3396596, -0.3396617, -0.3396603, 
    -0.3396272, -0.3396288, -0.3396279, -0.3396295, -0.3396284, -0.3396334, 
    -0.3396349, -0.3396423, -0.3396393, -0.3396441, -0.3396399, -0.3396406, 
    -0.3396441, -0.3396401, -0.3396493, -0.3396429, -0.3396548, -0.3396483, 
    -0.3396552, -0.339654, -0.3396561, -0.3396578, -0.3396601, -0.3396643, 
    -0.3396633, -0.3396668, -0.3396311, -0.3396332, -0.339633, -0.3396353, 
    -0.3396369, -0.3396405, -0.3396463, -0.3396441, -0.3396481, -0.3396489, 
    -0.3396429, -0.3396465, -0.3396346, -0.3396364, -0.3396354, -0.3396313, 
    -0.3396445, -0.3396376, -0.3396504, -0.3396467, -0.3396576, -0.3396521, 
    -0.3396628, -0.3396672, -0.3396717, -0.3396766, -0.3396344, -0.339633, 
    -0.3396356, -0.339639, -0.3396424, -0.3396469, -0.3396474, -0.3396482, 
    -0.3396504, -0.3396522, -0.3396484, -0.3396527, -0.3396367, -0.3396451, 
    -0.3396324, -0.3396361, -0.3396389, -0.3396377, -0.3396439, -0.3396453, 
    -0.3396511, -0.3396482, -0.3396661, -0.3396581, -0.3396805, -0.3396742, 
    -0.3396325, -0.3396344, -0.3396411, -0.3396379, -0.3396472, -0.3396495, 
    -0.3396514, -0.3396537, -0.339654, -0.3396554, -0.3396531, -0.3396553, 
    -0.3396469, -0.3396507, -0.3396404, -0.3396429, -0.3396418, -0.3396405, 
    -0.3396444, -0.3396485, -0.3396486, -0.3396499, -0.3396533, -0.3396473, 
    -0.3396669, -0.3396546, -0.3396365, -0.3396401, -0.3396408, -0.3396394, 
    -0.3396493, -0.3396457, -0.3396554, -0.3396528, -0.3396571, -0.3396549, 
    -0.3396546, -0.3396519, -0.3396502, -0.3396458, -0.3396423, -0.3396396, 
    -0.3396402, -0.3396432, -0.3396487, -0.339654, -0.3396528, -0.3396568, 
    -0.3396465, -0.3396508, -0.3396491, -0.3396535, -0.339644, -0.3396518, 
    -0.339642, -0.3396429, -0.3396456, -0.339651, -0.3396523, -0.3396536, 
    -0.3396528, -0.3396489, -0.3396483, -0.3396456, -0.3396448, -0.3396427, 
    -0.339641, -0.3396425, -0.3396442, -0.3396489, -0.3396532, -0.3396578, 
    -0.339659, -0.3396643, -0.3396599, -0.339667, -0.3396607, -0.3396716, 
    -0.3396524, -0.3396607, -0.3396457, -0.3396474, -0.3396502, -0.339657, 
    -0.3396535, -0.3396577, -0.3396482, -0.3396433, -0.3396421, -0.3396397, 
    -0.3396422, -0.339642, -0.3396443, -0.3396435, -0.3396491, -0.3396461, 
    -0.3396546, -0.3396576, -0.3396665, -0.3396718, -0.3396774, -0.3396799, 
    -0.3396806, -0.3396809 ;

 TAUY =
  -0.3396222, -0.3396269, -0.339626, -0.3396298, -0.3396277, -0.3396302, 
    -0.3396232, -0.3396271, -0.3396246, -0.3396227, -0.3396372, -0.33963, 
    -0.3396452, -0.3396405, -0.3396525, -0.3396444, -0.3396542, -0.3396524, 
    -0.339658, -0.3396564, -0.3396634, -0.3396588, -0.3396672, -0.3396624, 
    -0.3396631, -0.3396586, -0.3396315, -0.3396362, -0.3396312, -0.3396319, 
    -0.3396316, -0.3396277, -0.3396257, -0.3396219, -0.3396226, -0.3396255, 
    -0.3396322, -0.3396299, -0.3396358, -0.3396357, -0.3396423, -0.3396393, 
    -0.3396504, -0.3396473, -0.3396565, -0.3396541, -0.3396564, -0.3396557, 
    -0.3396564, -0.339653, -0.3396544, -0.3396514, -0.3396398, -0.3396432, 
    -0.3396331, -0.3396271, -0.3396233, -0.3396206, -0.339621, -0.3396217, 
    -0.3396255, -0.3396291, -0.3396319, -0.3396338, -0.3396356, -0.3396411, 
    -0.3396442, -0.339651, -0.3396499, -0.3396519, -0.3396539, -0.3396572, 
    -0.3396567, -0.3396581, -0.3396519, -0.339656, -0.3396492, -0.339651, 
    -0.3396358, -0.3396305, -0.3396281, -0.3396262, -0.3396213, -0.3396246, 
    -0.3396233, -0.3396266, -0.3396286, -0.3396276, -0.3396338, -0.3396313, 
    -0.3396444, -0.3396387, -0.3396537, -0.3396501, -0.3396546, -0.3396523, 
    -0.3396561, -0.3396527, -0.3396587, -0.33966, -0.3396591, -0.3396626, 
    -0.3396525, -0.3396563, -0.3396275, -0.3396277, -0.3396285, -0.3396251, 
    -0.3396249, -0.3396219, -0.3396246, -0.3396257, -0.3396287, -0.3396304, 
    -0.3396321, -0.3396358, -0.3396401, -0.339646, -0.3396503, -0.3396533, 
    -0.3396515, -0.339653, -0.3396513, -0.3396505, -0.3396595, -0.3396544, 
    -0.3396621, -0.3396617, -0.3396582, -0.3396617, -0.3396278, -0.3396269, 
    -0.3396236, -0.3396262, -0.3396215, -0.3396241, -0.3396255, -0.3396313, 
    -0.3396327, -0.3396339, -0.3396363, -0.3396394, -0.3396448, -0.3396496, 
    -0.3396541, -0.3396537, -0.3396538, -0.3396548, -0.3396524, -0.3396552, 
    -0.3396556, -0.3396544, -0.3396616, -0.3396596, -0.3396617, -0.3396603, 
    -0.3396272, -0.3396288, -0.3396279, -0.3396295, -0.3396284, -0.3396334, 
    -0.3396349, -0.3396423, -0.3396393, -0.3396441, -0.3396399, -0.3396406, 
    -0.3396441, -0.3396401, -0.3396493, -0.3396429, -0.3396548, -0.3396483, 
    -0.3396552, -0.339654, -0.3396561, -0.3396578, -0.3396601, -0.3396643, 
    -0.3396633, -0.3396668, -0.3396311, -0.3396332, -0.339633, -0.3396353, 
    -0.3396369, -0.3396405, -0.3396463, -0.3396441, -0.3396481, -0.3396489, 
    -0.3396429, -0.3396465, -0.3396346, -0.3396364, -0.3396354, -0.3396313, 
    -0.3396445, -0.3396376, -0.3396504, -0.3396467, -0.3396576, -0.3396521, 
    -0.3396628, -0.3396672, -0.3396717, -0.3396766, -0.3396344, -0.339633, 
    -0.3396356, -0.339639, -0.3396424, -0.3396469, -0.3396474, -0.3396482, 
    -0.3396504, -0.3396522, -0.3396484, -0.3396527, -0.3396367, -0.3396451, 
    -0.3396324, -0.3396361, -0.3396389, -0.3396377, -0.3396439, -0.3396453, 
    -0.3396511, -0.3396482, -0.3396661, -0.3396581, -0.3396805, -0.3396742, 
    -0.3396325, -0.3396344, -0.3396411, -0.3396379, -0.3396472, -0.3396495, 
    -0.3396514, -0.3396537, -0.339654, -0.3396554, -0.3396531, -0.3396553, 
    -0.3396469, -0.3396507, -0.3396404, -0.3396429, -0.3396418, -0.3396405, 
    -0.3396444, -0.3396485, -0.3396486, -0.3396499, -0.3396533, -0.3396473, 
    -0.3396669, -0.3396546, -0.3396365, -0.3396401, -0.3396408, -0.3396394, 
    -0.3396493, -0.3396457, -0.3396554, -0.3396528, -0.3396571, -0.3396549, 
    -0.3396546, -0.3396519, -0.3396502, -0.3396458, -0.3396423, -0.3396396, 
    -0.3396402, -0.3396432, -0.3396487, -0.339654, -0.3396528, -0.3396568, 
    -0.3396465, -0.3396508, -0.3396491, -0.3396535, -0.339644, -0.3396518, 
    -0.339642, -0.3396429, -0.3396456, -0.339651, -0.3396523, -0.3396536, 
    -0.3396528, -0.3396489, -0.3396483, -0.3396456, -0.3396448, -0.3396427, 
    -0.339641, -0.3396425, -0.3396442, -0.3396489, -0.3396532, -0.3396578, 
    -0.339659, -0.3396643, -0.3396599, -0.339667, -0.3396607, -0.3396716, 
    -0.3396524, -0.3396607, -0.3396457, -0.3396474, -0.3396502, -0.339657, 
    -0.3396535, -0.3396577, -0.3396482, -0.3396433, -0.3396421, -0.3396397, 
    -0.3396422, -0.339642, -0.3396443, -0.3396435, -0.3396491, -0.3396461, 
    -0.3396546, -0.3396576, -0.3396665, -0.3396718, -0.3396774, -0.3396799, 
    -0.3396806, -0.3396809 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.7812, 261.8008, 261.797, 261.8128, 261.804, 261.8144, 261.7852, 
    261.8016, 261.7911, 261.783, 261.8434, 261.8135, 261.8745, 261.8554, 
    261.9033, 261.8715, 261.9098, 261.9024, 261.9245, 261.9182, 261.9464, 
    261.9274, 261.9611, 261.9419, 261.9449, 261.9268, 261.8195, 261.8396, 
    261.8183, 261.8212, 261.8199, 261.8042, 261.7963, 261.7798, 261.7828, 
    261.7949, 261.8225, 261.8131, 261.8367, 261.8362, 261.8624, 261.8506, 
    261.8947, 261.8822, 261.9185, 261.9093, 261.918, 261.9154, 261.9181, 
    261.9047, 261.9104, 261.8987, 261.8528, 261.8663, 261.8261, 261.8019, 
    261.7859, 261.7746, 261.7762, 261.7792, 261.795, 261.8098, 261.8211, 
    261.8287, 261.8361, 261.8586, 261.8705, 261.8973, 261.8925, 261.9006, 
    261.9084, 261.9215, 261.9194, 261.9251, 261.9004, 261.9168, 261.8897, 
    261.8971, 261.8381, 261.8156, 261.8061, 261.7977, 261.7774, 261.7914, 
    261.7859, 261.7991, 261.8075, 261.8033, 261.8289, 261.8189, 261.8712, 
    261.8487, 261.9075, 261.8935, 261.9109, 261.902, 261.9172, 261.9035, 
    261.9273, 261.9325, 261.9289, 261.9425, 261.9028, 261.918, 261.8032, 
    261.8039, 261.807, 261.7932, 261.7923, 261.7797, 261.791, 261.7957, 
    261.808, 261.8152, 261.822, 261.8371, 261.8539, 261.8774, 261.8943, 
    261.9057, 261.8987, 261.9049, 261.898, 261.8948, 261.9305, 261.9105, 
    261.9406, 261.9389, 261.9253, 261.9391, 261.8044, 261.8005, 261.787, 
    261.7975, 261.7783, 261.7891, 261.7952, 261.8191, 261.8244, 261.8293, 
    261.8389, 261.8512, 261.8728, 261.8917, 261.9089, 261.9076, 261.9081, 
    261.9119, 261.9024, 261.9135, 261.9153, 261.9105, 261.9387, 261.9306, 
    261.9389, 261.9336, 261.8017, 261.8083, 261.8047, 261.8114, 261.8067, 
    261.8275, 261.8337, 261.8629, 261.851, 261.87, 261.8529, 261.8559, 
    261.8706, 261.8538, 261.8906, 261.8657, 261.912, 261.8871, 261.9136, 
    261.9088, 261.9168, 261.9239, 261.9329, 261.9494, 261.9456, 261.9594, 
    261.818, 261.8265, 261.8257, 261.8346, 261.8412, 261.8554, 261.8782, 
    261.8697, 261.8854, 261.8886, 261.8647, 261.8793, 261.8322, 261.8398, 
    261.8352, 261.8187, 261.8716, 261.8445, 261.8947, 261.8799, 261.9229, 
    261.9015, 261.9435, 261.9614, 261.9783, 261.998, 261.8311, 261.8254, 
    261.8357, 261.8499, 261.8632, 261.8808, 261.8826, 261.8859, 261.8945, 
    261.9016, 261.887, 261.9034, 261.8415, 261.874, 261.8232, 261.8385, 
    261.8491, 261.8445, 261.8687, 261.8744, 261.8976, 261.8856, 261.957, 
    261.9254, 262.0131, 261.9886, 261.8234, 261.8311, 261.8581, 261.8452, 
    261.882, 261.891, 261.8984, 261.9078, 261.9088, 261.9144, 261.9052, 
    261.914, 261.8809, 261.8957, 261.855, 261.8649, 261.8604, 261.8554, 
    261.8708, 261.8872, 261.8875, 261.8928, 261.9076, 261.8821, 261.961, 
    261.9123, 261.8396, 261.8545, 261.8566, 261.8509, 261.8901, 261.8759, 
    261.9142, 261.9039, 261.9208, 261.9124, 261.9112, 261.9003, 261.8936, 
    261.8766, 261.8627, 261.8517, 261.8542, 261.8663, 261.8882, 261.9089, 
    261.9044, 261.9196, 261.8793, 261.8962, 261.8897, 261.9067, 261.8694, 
    261.9011, 261.8613, 261.8648, 261.8756, 261.8973, 261.9022, 261.9073, 
    261.9041, 261.8887, 261.8862, 261.8754, 261.8723, 261.864, 261.8572, 
    261.8635, 261.87, 261.8888, 261.9056, 261.924, 261.9285, 261.95, 
    261.9325, 261.9613, 261.9368, 261.9792, 261.903, 261.9361, 261.8761, 
    261.8826, 261.8943, 261.9211, 261.9066, 261.9235, 261.8861, 261.8667, 
    261.8617, 261.8524, 261.8619, 261.8611, 261.8703, 261.8674, 261.8894, 
    261.8776, 261.9111, 261.9234, 261.958, 261.9792, 262.0008, 262.0103, 
    262.0132, 262.0144 ;

 TG_R =
  261.7812, 261.8008, 261.797, 261.8128, 261.804, 261.8144, 261.7852, 
    261.8016, 261.7911, 261.783, 261.8434, 261.8135, 261.8745, 261.8554, 
    261.9033, 261.8715, 261.9098, 261.9024, 261.9245, 261.9182, 261.9464, 
    261.9274, 261.9611, 261.9419, 261.9449, 261.9268, 261.8195, 261.8396, 
    261.8183, 261.8212, 261.8199, 261.8042, 261.7963, 261.7798, 261.7828, 
    261.7949, 261.8225, 261.8131, 261.8367, 261.8362, 261.8624, 261.8506, 
    261.8947, 261.8822, 261.9185, 261.9093, 261.918, 261.9154, 261.9181, 
    261.9047, 261.9104, 261.8987, 261.8528, 261.8663, 261.8261, 261.8019, 
    261.7859, 261.7746, 261.7762, 261.7792, 261.795, 261.8098, 261.8211, 
    261.8287, 261.8361, 261.8586, 261.8705, 261.8973, 261.8925, 261.9006, 
    261.9084, 261.9215, 261.9194, 261.9251, 261.9004, 261.9168, 261.8897, 
    261.8971, 261.8381, 261.8156, 261.8061, 261.7977, 261.7774, 261.7914, 
    261.7859, 261.7991, 261.8075, 261.8033, 261.8289, 261.8189, 261.8712, 
    261.8487, 261.9075, 261.8935, 261.9109, 261.902, 261.9172, 261.9035, 
    261.9273, 261.9325, 261.9289, 261.9425, 261.9028, 261.918, 261.8032, 
    261.8039, 261.807, 261.7932, 261.7923, 261.7797, 261.791, 261.7957, 
    261.808, 261.8152, 261.822, 261.8371, 261.8539, 261.8774, 261.8943, 
    261.9057, 261.8987, 261.9049, 261.898, 261.8948, 261.9305, 261.9105, 
    261.9406, 261.9389, 261.9253, 261.9391, 261.8044, 261.8005, 261.787, 
    261.7975, 261.7783, 261.7891, 261.7952, 261.8191, 261.8244, 261.8293, 
    261.8389, 261.8512, 261.8728, 261.8917, 261.9089, 261.9076, 261.9081, 
    261.9119, 261.9024, 261.9135, 261.9153, 261.9105, 261.9387, 261.9306, 
    261.9389, 261.9336, 261.8017, 261.8083, 261.8047, 261.8114, 261.8067, 
    261.8275, 261.8337, 261.8629, 261.851, 261.87, 261.8529, 261.8559, 
    261.8706, 261.8538, 261.8906, 261.8657, 261.912, 261.8871, 261.9136, 
    261.9088, 261.9168, 261.9239, 261.9329, 261.9494, 261.9456, 261.9594, 
    261.818, 261.8265, 261.8257, 261.8346, 261.8412, 261.8554, 261.8782, 
    261.8697, 261.8854, 261.8886, 261.8647, 261.8793, 261.8322, 261.8398, 
    261.8352, 261.8187, 261.8716, 261.8445, 261.8947, 261.8799, 261.9229, 
    261.9015, 261.9435, 261.9614, 261.9783, 261.998, 261.8311, 261.8254, 
    261.8357, 261.8499, 261.8632, 261.8808, 261.8826, 261.8859, 261.8945, 
    261.9016, 261.887, 261.9034, 261.8415, 261.874, 261.8232, 261.8385, 
    261.8491, 261.8445, 261.8687, 261.8744, 261.8976, 261.8856, 261.957, 
    261.9254, 262.0131, 261.9886, 261.8234, 261.8311, 261.8581, 261.8452, 
    261.882, 261.891, 261.8984, 261.9078, 261.9088, 261.9144, 261.9052, 
    261.914, 261.8809, 261.8957, 261.855, 261.8649, 261.8604, 261.8554, 
    261.8708, 261.8872, 261.8875, 261.8928, 261.9076, 261.8821, 261.961, 
    261.9123, 261.8396, 261.8545, 261.8566, 261.8509, 261.8901, 261.8759, 
    261.9142, 261.9039, 261.9208, 261.9124, 261.9112, 261.9003, 261.8936, 
    261.8766, 261.8627, 261.8517, 261.8542, 261.8663, 261.8882, 261.9089, 
    261.9044, 261.9196, 261.8793, 261.8962, 261.8897, 261.9067, 261.8694, 
    261.9011, 261.8613, 261.8648, 261.8756, 261.8973, 261.9022, 261.9073, 
    261.9041, 261.8887, 261.8862, 261.8754, 261.8723, 261.864, 261.8572, 
    261.8635, 261.87, 261.8888, 261.9056, 261.924, 261.9285, 261.95, 
    261.9325, 261.9613, 261.9368, 261.9792, 261.903, 261.9361, 261.8761, 
    261.8826, 261.8943, 261.9211, 261.9066, 261.9235, 261.8861, 261.8667, 
    261.8617, 261.8524, 261.8619, 261.8611, 261.8703, 261.8674, 261.8894, 
    261.8776, 261.9111, 261.9234, 261.958, 261.9792, 262.0008, 262.0103, 
    262.0132, 262.0144 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  255.2182, 255.218, 255.218, 255.218, 255.218, 255.2179, 255.2181, 255.218, 
    255.2181, 255.2182, 255.2177, 255.2179, 255.2176, 255.2177, 255.2175, 
    255.2176, 255.2175, 255.2175, 255.2174, 255.2175, 255.2173, 255.2174, 
    255.2173, 255.2173, 255.2173, 255.2174, 255.2179, 255.2178, 255.2179, 
    255.2179, 255.2179, 255.218, 255.218, 255.2182, 255.2182, 255.2181, 
    255.2179, 255.218, 255.2178, 255.2178, 255.2177, 255.2178, 255.2175, 
    255.2176, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 
    255.2175, 255.2175, 255.2177, 255.2177, 255.2179, 255.218, 255.2181, 
    255.2182, 255.2182, 255.2182, 255.2181, 255.218, 255.2179, 255.2179, 
    255.2178, 255.2177, 255.2176, 255.2175, 255.2176, 255.2175, 255.2175, 
    255.2174, 255.2174, 255.2174, 255.2175, 255.2174, 255.2176, 255.2175, 
    255.2178, 255.2179, 255.218, 255.218, 255.2182, 255.2181, 255.2181, 
    255.218, 255.218, 255.218, 255.2179, 255.2179, 255.2176, 255.2178, 
    255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 255.2174, 
    255.2174, 255.2174, 255.2174, 255.2175, 255.2174, 255.218, 255.218, 
    255.218, 255.2181, 255.2181, 255.2182, 255.2181, 255.2181, 255.218, 
    255.2179, 255.2179, 255.2178, 255.2177, 255.2176, 255.2175, 255.2175, 
    255.2175, 255.2175, 255.2175, 255.2175, 255.2174, 255.2175, 255.2174, 
    255.2174, 255.2174, 255.2174, 255.218, 255.218, 255.2181, 255.2181, 
    255.2182, 255.2181, 255.2181, 255.2179, 255.2179, 255.2179, 255.2178, 
    255.2177, 255.2176, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 
    255.2175, 255.2175, 255.2175, 255.2175, 255.2174, 255.2174, 255.2174, 
    255.2174, 255.218, 255.218, 255.218, 255.218, 255.218, 255.2179, 
    255.2178, 255.2177, 255.2177, 255.2176, 255.2177, 255.2177, 255.2176, 
    255.2177, 255.2175, 255.2177, 255.2175, 255.2175, 255.2175, 255.2175, 
    255.2175, 255.2174, 255.2174, 255.2173, 255.2173, 255.2173, 255.2179, 
    255.2179, 255.2179, 255.2178, 255.2178, 255.2177, 255.2176, 255.2177, 
    255.2176, 255.2176, 255.2177, 255.2176, 255.2178, 255.2178, 255.2178, 
    255.2179, 255.2176, 255.2178, 255.2175, 255.2176, 255.2174, 255.2175, 
    255.2173, 255.2173, 255.2173, 255.2172, 255.2178, 255.2179, 255.2178, 
    255.2177, 255.2177, 255.2176, 255.2176, 255.2176, 255.2175, 255.2175, 
    255.2176, 255.2175, 255.2178, 255.2176, 255.2179, 255.2178, 255.2177, 
    255.2178, 255.2177, 255.2176, 255.2175, 255.2176, 255.2173, 255.2174, 
    255.2172, 255.2172, 255.2179, 255.2179, 255.2177, 255.2178, 255.2176, 
    255.2176, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 255.2175, 
    255.2176, 255.2175, 255.2177, 255.2177, 255.2177, 255.2177, 255.2177, 
    255.2176, 255.2176, 255.2175, 255.2174, 255.2176, 255.2172, 255.2174, 
    255.2178, 255.2177, 255.2177, 255.2178, 255.2176, 255.2176, 255.2175, 
    255.2175, 255.2174, 255.2175, 255.2175, 255.2175, 255.2175, 255.2176, 
    255.2177, 255.2178, 255.2177, 255.2177, 255.2176, 255.2175, 255.2175, 
    255.2175, 255.2176, 255.2175, 255.2176, 255.2175, 255.2177, 255.2175, 
    255.2177, 255.2177, 255.2176, 255.2175, 255.2175, 255.2175, 255.2175, 
    255.2176, 255.2176, 255.2176, 255.2176, 255.2177, 255.2177, 255.2177, 
    255.2177, 255.2176, 255.2175, 255.2174, 255.2174, 255.2173, 255.2174, 
    255.2172, 255.2173, 255.2172, 255.2175, 255.2173, 255.2176, 255.2176, 
    255.2175, 255.2174, 255.2175, 255.2174, 255.2176, 255.2177, 255.2177, 
    255.2177, 255.2177, 255.2177, 255.2177, 255.2177, 255.2176, 255.2176, 
    255.2175, 255.2174, 255.2173, 255.2172, 255.2172, 255.2172, 255.2172, 
    255.2172 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24018, 18.24017, 18.24019, 
    18.24018, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24017, 18.24016, 18.24016, 18.24018, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 
    18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.2401, 18.24012, 
    18.24011, 18.24015, 18.24017, 18.24017, 18.24018, 18.24019, 18.24018, 
    18.24019, 18.24018, 18.24017, 18.24018, 18.24016, 18.24016, 18.24013, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24018, 
    18.24018, 18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24017, 18.24017, 18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 
    18.24011, 18.24011, 18.24011, 18.24011, 18.24011, 18.24009, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24019, 
    18.24018, 18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24008, 18.24009, 18.24018, 18.24017, 18.24017, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24014, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24014, 18.24012, 18.24013, 18.2401, 18.24012, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24008, 18.24008, 18.24007, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.24012, 18.24013, 18.24012, 18.24016, 18.24015, 
    18.24015, 18.24016, 18.24013, 18.24015, 18.24011, 18.24012, 18.2401, 
    18.24011, 18.24008, 18.24007, 18.24006, 18.24005, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24014, 18.24012, 18.24012, 18.24012, 18.24011, 
    18.24011, 18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 
    18.24014, 18.24015, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 
    18.24009, 18.24003, 18.24005, 18.24016, 18.24016, 18.24014, 18.24015, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 
    18.2401, 18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 
    18.2401, 18.24015, 18.24014, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 18.24011, 
    18.24013, 18.24014, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 
    18.24011, 18.2401, 18.24012, 18.24011, 18.24012, 18.24011, 18.24013, 
    18.24011, 18.24014, 18.24013, 18.24013, 18.24011, 18.24011, 18.2401, 
    18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24014, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.2401, 18.24009, 18.24008, 
    18.24009, 18.24007, 18.24009, 18.24006, 18.24011, 18.24009, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24011, 18.2401, 18.24012, 18.24013, 
    18.24014, 18.24014, 18.24014, 18.24014, 18.24013, 18.24013, 18.24012, 
    18.24013, 18.2401, 18.2401, 18.24007, 18.24006, 18.24004, 18.24004, 
    18.24003, 18.24003 ;

 TOTCOLCH4 =
  4.77247e-06, 4.633464e-06, 4.660348e-06, 4.549268e-06, 4.610744e-06, 
    4.538219e-06, 4.744147e-06, 4.627979e-06, 4.701994e-06, 4.759889e-06, 
    4.337125e-06, 4.544342e-06, 4.126591e-06, 4.255308e-06, 3.935448e-06, 
    4.146495e-06, 3.893515e-06, 3.941476e-06, 3.797986e-06, 3.838838e-06, 
    3.658026e-06, 3.779201e-06, 3.565947e-06, 3.686799e-06, 3.667763e-06, 
    3.783229e-06, 4.502303e-06, 4.362681e-06, 4.510634e-06, 4.490587e-06, 
    4.49958e-06, 4.609466e-06, 4.665281e-06, 4.783177e-06, 4.761679e-06, 
    4.675139e-06, 4.481586e-06, 4.546886e-06, 4.383151e-06, 4.386819e-06, 
    4.207664e-06, 4.28802e-06, 3.992041e-06, 4.075172e-06, 3.837129e-06, 
    3.896364e-06, 3.8399e-06, 3.856982e-06, 3.839678e-06, 3.926725e-06, 
    3.889317e-06, 3.966329e-06, 4.272915e-06, 4.181717e-06, 4.456352e-06, 
    4.625258e-06, 4.739023e-06, 4.820482e-06, 4.808928e-06, 4.786936e-06, 
    4.674635e-06, 4.570138e-06, 4.49121e-06, 4.438756e-06, 4.387347e-06, 
    4.233362e-06, 4.152905e-06, 3.975322e-06, 4.007114e-06, 3.953332e-06, 
    3.902281e-06, 3.817257e-06, 3.831193e-06, 3.793948e-06, 3.954753e-06, 
    3.847529e-06, 4.025273e-06, 3.976287e-06, 4.373377e-06, 4.52923e-06, 
    4.59618e-06, 4.655173e-06, 4.800053e-06, 4.69979e-06, 4.739202e-06, 
    4.645686e-06, 4.58669e-06, 4.615828e-06, 4.437326e-06, 4.506346e-06, 
    4.148158e-06, 4.300788e-06, 3.908219e-06, 4.00058e-06, 3.886232e-06, 
    3.94439e-06, 3.844985e-06, 3.934395e-06, 3.780133e-06, 3.746924e-06, 
    3.769602e-06, 3.682854e-06, 3.939379e-06, 3.839897e-06, 4.616644e-06, 
    4.611885e-06, 4.58975e-06, 4.687405e-06, 4.693411e-06, 4.783765e-06, 
    4.703334e-06, 4.669263e-06, 4.583283e-06, 4.532754e-06, 4.484956e-06, 
    4.380667e-06, 4.265504e-06, 4.106834e-06, 3.994563e-06, 3.920108e-06, 
    3.965688e-06, 3.925434e-06, 3.970444e-06, 3.991624e-06, 3.759349e-06, 
    3.888967e-06, 3.695272e-06, 3.705869e-06, 3.793063e-06, 3.704674e-06, 
    4.608546e-06, 4.635949e-06, 4.731638e-06, 4.656679e-06, 4.793651e-06, 
    4.716759e-06, 4.672793e-06, 4.50489e-06, 4.468378e-06, 4.43463e-06, 
    4.368324e-06, 4.28389e-06, 4.137591e-06, 4.012212e-06, 3.899322e-06, 
    3.907543e-06, 3.904647e-06, 3.879614e-06, 3.941755e-06, 3.869457e-06, 
    3.857381e-06, 3.888987e-06, 3.707289e-06, 3.75878e-06, 3.706095e-06, 
    3.739578e-06, 4.627035e-06, 4.581008e-06, 4.605853e-06, 4.559181e-06, 
    4.592036e-06, 4.446741e-06, 4.403588e-06, 4.204221e-06, 4.285542e-06, 
    4.156465e-06, 4.272351e-06, 4.251709e-06, 4.152269e-06, 4.266054e-06, 
    4.019071e-06, 4.185763e-06, 3.878642e-06, 4.042397e-06, 3.868485e-06, 
    3.899806e-06, 3.848017e-06, 3.801905e-06, 3.744275e-06, 3.639024e-06, 
    3.66327e-06, 3.576077e-06, 4.512777e-06, 4.453781e-06, 4.458968e-06, 
    4.397576e-06, 4.352419e-06, 4.255281e-06, 4.101573e-06, 4.159071e-06, 
    4.053806e-06, 4.032821e-06, 4.19286e-06, 4.09425e-06, 4.414499e-06, 
    4.362006e-06, 4.393231e-06, 4.508106e-06, 4.145778e-06, 4.329997e-06, 
    3.992718e-06, 4.090362e-06, 3.808463e-06, 3.947478e-06, 3.676649e-06, 
    3.563643e-06, 3.458864e-06, 3.338296e-06, 4.421738e-06, 4.461657e-06, 
    4.390303e-06, 4.292428e-06, 4.202537e-06, 4.084374e-06, 4.072376e-06, 
    4.05044e-06, 3.993885e-06, 3.946614e-06, 4.043508e-06, 3.934805e-06, 
    4.349857e-06, 4.129965e-06, 4.476783e-06, 4.371001e-06, 4.298173e-06, 
    4.33006e-06, 4.165668e-06, 4.127345e-06, 3.973299e-06, 4.052598e-06, 
    3.591371e-06, 3.79219e-06, 3.24791e-06, 3.395914e-06, 4.47564e-06, 
    4.421879e-06, 4.23706e-06, 4.324551e-06, 4.076545e-06, 4.016532e-06, 
    3.968055e-06, 3.906473e-06, 3.899857e-06, 3.863612e-06, 3.923088e-06, 
    3.865956e-06, 4.084124e-06, 3.985945e-06, 4.258012e-06, 4.191027e-06, 
    4.221785e-06, 4.255636e-06, 4.151559e-06, 4.041973e-06, 4.039658e-06, 
    4.004814e-06, 3.907356e-06, 4.075554e-06, 3.565812e-06, 3.876816e-06, 
    4.36359e-06, 4.261471e-06, 4.24699e-06, 4.286353e-06, 4.02253e-06, 
    4.117228e-06, 3.864495e-06, 3.932069e-06, 3.821642e-06, 3.876329e-06, 
    3.884405e-06, 3.95525e-06, 3.999655e-06, 4.112862e-06, 4.206051e-06, 
    4.280635e-06, 4.26324e-06, 4.181497e-06, 4.035317e-06, 3.899253e-06, 
    3.928871e-06, 3.829982e-06, 4.0943e-06, 3.982464e-06, 4.025515e-06, 
    3.913711e-06, 4.160601e-06, 3.949883e-06, 4.215268e-06, 4.191684e-06, 
    4.119119e-06, 3.974922e-06, 3.943358e-06, 3.909765e-06, 3.93048e-06, 
    4.031639e-06, 4.04833e-06, 4.120878e-06, 4.141008e-06, 4.196815e-06, 
    4.243271e-06, 4.200813e-06, 4.156434e-06, 4.031601e-06, 3.920607e-06, 
    3.801249e-06, 3.772309e-06, 3.635535e-06, 3.746678e-06, 3.564112e-06, 
    3.719028e-06, 3.452871e-06, 3.937845e-06, 3.723654e-06, 4.115835e-06, 
    4.07271e-06, 3.995232e-06, 3.820166e-06, 3.914234e-06, 3.804334e-06, 
    4.048986e-06, 4.178684e-06, 4.212563e-06, 4.276082e-06, 4.211116e-06, 
    4.216383e-06, 4.154609e-06, 4.174415e-06, 4.027487e-06, 4.106108e-06, 
    3.884606e-06, 3.8052e-06, 3.585164e-06, 3.45337e-06, 3.321678e-06, 
    3.264326e-06, 3.246967e-06, 3.239724e-06 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24018, 18.24017, 18.24019, 
    18.24018, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24017, 18.24016, 18.24016, 18.24018, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 
    18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.2401, 18.24012, 
    18.24011, 18.24015, 18.24017, 18.24017, 18.24018, 18.24019, 18.24018, 
    18.24019, 18.24018, 18.24017, 18.24018, 18.24016, 18.24016, 18.24013, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24018, 
    18.24018, 18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24017, 18.24017, 18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 
    18.24011, 18.24011, 18.24011, 18.24011, 18.24011, 18.24009, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24019, 
    18.24018, 18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24008, 18.24009, 18.24018, 18.24017, 18.24017, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24014, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24014, 18.24012, 18.24013, 18.2401, 18.24012, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24008, 18.24008, 18.24007, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.24012, 18.24013, 18.24012, 18.24016, 18.24015, 
    18.24015, 18.24016, 18.24013, 18.24015, 18.24011, 18.24012, 18.2401, 
    18.24011, 18.24008, 18.24007, 18.24006, 18.24005, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24014, 18.24012, 18.24012, 18.24012, 18.24011, 
    18.24011, 18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 
    18.24014, 18.24015, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 
    18.24009, 18.24003, 18.24005, 18.24016, 18.24016, 18.24014, 18.24015, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 
    18.2401, 18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 
    18.2401, 18.24015, 18.24014, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 18.24011, 
    18.24013, 18.24014, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 
    18.24011, 18.2401, 18.24012, 18.24011, 18.24012, 18.24011, 18.24013, 
    18.24011, 18.24014, 18.24013, 18.24013, 18.24011, 18.24011, 18.2401, 
    18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24014, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.2401, 18.24009, 18.24008, 
    18.24009, 18.24007, 18.24009, 18.24006, 18.24011, 18.24009, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24011, 18.2401, 18.24012, 18.24013, 
    18.24014, 18.24014, 18.24014, 18.24014, 18.24013, 18.24013, 18.24012, 
    18.24013, 18.2401, 18.2401, 18.24007, 18.24006, 18.24004, 18.24004, 
    18.24003, 18.24003 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976299e-05, 5.976284e-05, 5.976287e-05, 5.976275e-05, 5.976282e-05, 
    5.976274e-05, 5.976296e-05, 5.976284e-05, 5.976292e-05, 5.976298e-05, 
    5.976252e-05, 5.976275e-05, 5.976229e-05, 5.976243e-05, 5.976207e-05, 
    5.976231e-05, 5.976202e-05, 5.976207e-05, 5.976191e-05, 5.976195e-05, 
    5.976174e-05, 5.976189e-05, 5.976163e-05, 5.976178e-05, 5.976175e-05, 
    5.976189e-05, 5.97627e-05, 5.976255e-05, 5.976271e-05, 5.976269e-05, 
    5.97627e-05, 5.976282e-05, 5.976288e-05, 5.9763e-05, 5.976298e-05, 
    5.976289e-05, 5.976268e-05, 5.976275e-05, 5.976257e-05, 5.976257e-05, 
    5.976238e-05, 5.976246e-05, 5.976213e-05, 5.976223e-05, 5.976195e-05, 
    5.976202e-05, 5.976195e-05, 5.976198e-05, 5.976195e-05, 5.976206e-05, 
    5.976201e-05, 5.97621e-05, 5.976245e-05, 5.976235e-05, 5.976265e-05, 
    5.976284e-05, 5.976296e-05, 5.976304e-05, 5.976303e-05, 5.976301e-05, 
    5.976289e-05, 5.976277e-05, 5.976269e-05, 5.976263e-05, 5.976258e-05, 
    5.976241e-05, 5.976231e-05, 5.976211e-05, 5.976215e-05, 5.976209e-05, 
    5.976203e-05, 5.976193e-05, 5.976195e-05, 5.97619e-05, 5.976209e-05, 
    5.976197e-05, 5.976217e-05, 5.976211e-05, 5.976256e-05, 5.976273e-05, 
    5.97628e-05, 5.976286e-05, 5.976302e-05, 5.976291e-05, 5.976296e-05, 
    5.976286e-05, 5.976279e-05, 5.976282e-05, 5.976263e-05, 5.97627e-05, 
    5.976231e-05, 5.976248e-05, 5.976203e-05, 5.976214e-05, 5.976201e-05, 
    5.976208e-05, 5.976196e-05, 5.976207e-05, 5.976189e-05, 5.976185e-05, 
    5.976187e-05, 5.976177e-05, 5.976207e-05, 5.976195e-05, 5.976282e-05, 
    5.976282e-05, 5.976279e-05, 5.97629e-05, 5.976291e-05, 5.9763e-05, 
    5.976292e-05, 5.976288e-05, 5.976279e-05, 5.976273e-05, 5.976268e-05, 
    5.976257e-05, 5.976244e-05, 5.976226e-05, 5.976214e-05, 5.976205e-05, 
    5.97621e-05, 5.976206e-05, 5.976211e-05, 5.976213e-05, 5.976186e-05, 
    5.976201e-05, 5.976179e-05, 5.97618e-05, 5.97619e-05, 5.97618e-05, 
    5.976282e-05, 5.976285e-05, 5.976295e-05, 5.976287e-05, 5.976301e-05, 
    5.976293e-05, 5.976289e-05, 5.97627e-05, 5.976266e-05, 5.976263e-05, 
    5.976255e-05, 5.976246e-05, 5.97623e-05, 5.976215e-05, 5.976202e-05, 
    5.976203e-05, 5.976203e-05, 5.9762e-05, 5.976207e-05, 5.976199e-05, 
    5.976198e-05, 5.976201e-05, 5.97618e-05, 5.976186e-05, 5.97618e-05, 
    5.976184e-05, 5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976276e-05, 
    5.97628e-05, 5.976264e-05, 5.976259e-05, 5.976237e-05, 5.976246e-05, 
    5.976232e-05, 5.976245e-05, 5.976242e-05, 5.976231e-05, 5.976244e-05, 
    5.976216e-05, 5.976235e-05, 5.9762e-05, 5.976219e-05, 5.976199e-05, 
    5.976203e-05, 5.976197e-05, 5.976191e-05, 5.976185e-05, 5.976172e-05, 
    5.976175e-05, 5.976165e-05, 5.976271e-05, 5.976265e-05, 5.976265e-05, 
    5.976259e-05, 5.976254e-05, 5.976243e-05, 5.976226e-05, 5.976232e-05, 
    5.97622e-05, 5.976218e-05, 5.976236e-05, 5.976225e-05, 5.976261e-05, 
    5.976255e-05, 5.976258e-05, 5.976271e-05, 5.976231e-05, 5.976251e-05, 
    5.976213e-05, 5.976224e-05, 5.976192e-05, 5.976208e-05, 5.976177e-05, 
    5.976163e-05, 5.97615e-05, 5.976135e-05, 5.976261e-05, 5.976266e-05, 
    5.976258e-05, 5.976247e-05, 5.976237e-05, 5.976224e-05, 5.976222e-05, 
    5.97622e-05, 5.976213e-05, 5.976208e-05, 5.976219e-05, 5.976207e-05, 
    5.976253e-05, 5.976229e-05, 5.976267e-05, 5.976256e-05, 5.976247e-05, 
    5.976251e-05, 5.976233e-05, 5.976229e-05, 5.976211e-05, 5.97622e-05, 
    5.976166e-05, 5.97619e-05, 5.976124e-05, 5.976142e-05, 5.976267e-05, 
    5.976261e-05, 5.976241e-05, 5.97625e-05, 5.976223e-05, 5.976216e-05, 
    5.97621e-05, 5.976203e-05, 5.976203e-05, 5.976198e-05, 5.976205e-05, 
    5.976199e-05, 5.976224e-05, 5.976213e-05, 5.976243e-05, 5.976236e-05, 
    5.976239e-05, 5.976243e-05, 5.976231e-05, 5.976219e-05, 5.976219e-05, 
    5.976215e-05, 5.976203e-05, 5.976223e-05, 5.976163e-05, 5.9762e-05, 
    5.976255e-05, 5.976243e-05, 5.976242e-05, 5.976246e-05, 5.976217e-05, 
    5.976227e-05, 5.976198e-05, 5.976206e-05, 5.976194e-05, 5.9762e-05, 
    5.976201e-05, 5.976209e-05, 5.976214e-05, 5.976227e-05, 5.976237e-05, 
    5.976246e-05, 5.976244e-05, 5.976235e-05, 5.976218e-05, 5.976202e-05, 
    5.976206e-05, 5.976194e-05, 5.976225e-05, 5.976212e-05, 5.976217e-05, 
    5.976204e-05, 5.976232e-05, 5.976208e-05, 5.976238e-05, 5.976236e-05, 
    5.976227e-05, 5.976211e-05, 5.976207e-05, 5.976204e-05, 5.976206e-05, 
    5.976218e-05, 5.976219e-05, 5.976228e-05, 5.97623e-05, 5.976236e-05, 
    5.976242e-05, 5.976237e-05, 5.976232e-05, 5.976218e-05, 5.976205e-05, 
    5.976191e-05, 5.976188e-05, 5.976171e-05, 5.976185e-05, 5.976163e-05, 
    5.976182e-05, 5.97615e-05, 5.976207e-05, 5.976182e-05, 5.976227e-05, 
    5.976222e-05, 5.976214e-05, 5.976193e-05, 5.976204e-05, 5.976191e-05, 
    5.97622e-05, 5.976234e-05, 5.976238e-05, 5.976245e-05, 5.976238e-05, 
    5.976238e-05, 5.976231e-05, 5.976234e-05, 5.976217e-05, 5.976226e-05, 
    5.976201e-05, 5.976191e-05, 5.976166e-05, 5.97615e-05, 5.976133e-05, 
    5.976126e-05, 5.976124e-05, 5.976123e-05 ;

 TOTLITC_1m =
  5.976299e-05, 5.976284e-05, 5.976287e-05, 5.976275e-05, 5.976282e-05, 
    5.976274e-05, 5.976296e-05, 5.976284e-05, 5.976292e-05, 5.976298e-05, 
    5.976252e-05, 5.976275e-05, 5.976229e-05, 5.976243e-05, 5.976207e-05, 
    5.976231e-05, 5.976202e-05, 5.976207e-05, 5.976191e-05, 5.976195e-05, 
    5.976174e-05, 5.976189e-05, 5.976163e-05, 5.976178e-05, 5.976175e-05, 
    5.976189e-05, 5.97627e-05, 5.976255e-05, 5.976271e-05, 5.976269e-05, 
    5.97627e-05, 5.976282e-05, 5.976288e-05, 5.9763e-05, 5.976298e-05, 
    5.976289e-05, 5.976268e-05, 5.976275e-05, 5.976257e-05, 5.976257e-05, 
    5.976238e-05, 5.976246e-05, 5.976213e-05, 5.976223e-05, 5.976195e-05, 
    5.976202e-05, 5.976195e-05, 5.976198e-05, 5.976195e-05, 5.976206e-05, 
    5.976201e-05, 5.97621e-05, 5.976245e-05, 5.976235e-05, 5.976265e-05, 
    5.976284e-05, 5.976296e-05, 5.976304e-05, 5.976303e-05, 5.976301e-05, 
    5.976289e-05, 5.976277e-05, 5.976269e-05, 5.976263e-05, 5.976258e-05, 
    5.976241e-05, 5.976231e-05, 5.976211e-05, 5.976215e-05, 5.976209e-05, 
    5.976203e-05, 5.976193e-05, 5.976195e-05, 5.97619e-05, 5.976209e-05, 
    5.976197e-05, 5.976217e-05, 5.976211e-05, 5.976256e-05, 5.976273e-05, 
    5.97628e-05, 5.976286e-05, 5.976302e-05, 5.976291e-05, 5.976296e-05, 
    5.976286e-05, 5.976279e-05, 5.976282e-05, 5.976263e-05, 5.97627e-05, 
    5.976231e-05, 5.976248e-05, 5.976203e-05, 5.976214e-05, 5.976201e-05, 
    5.976208e-05, 5.976196e-05, 5.976207e-05, 5.976189e-05, 5.976185e-05, 
    5.976187e-05, 5.976177e-05, 5.976207e-05, 5.976195e-05, 5.976282e-05, 
    5.976282e-05, 5.976279e-05, 5.97629e-05, 5.976291e-05, 5.9763e-05, 
    5.976292e-05, 5.976288e-05, 5.976279e-05, 5.976273e-05, 5.976268e-05, 
    5.976257e-05, 5.976244e-05, 5.976226e-05, 5.976214e-05, 5.976205e-05, 
    5.97621e-05, 5.976206e-05, 5.976211e-05, 5.976213e-05, 5.976186e-05, 
    5.976201e-05, 5.976179e-05, 5.97618e-05, 5.97619e-05, 5.97618e-05, 
    5.976282e-05, 5.976285e-05, 5.976295e-05, 5.976287e-05, 5.976301e-05, 
    5.976293e-05, 5.976289e-05, 5.97627e-05, 5.976266e-05, 5.976263e-05, 
    5.976255e-05, 5.976246e-05, 5.97623e-05, 5.976215e-05, 5.976202e-05, 
    5.976203e-05, 5.976203e-05, 5.9762e-05, 5.976207e-05, 5.976199e-05, 
    5.976198e-05, 5.976201e-05, 5.97618e-05, 5.976186e-05, 5.97618e-05, 
    5.976184e-05, 5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976276e-05, 
    5.97628e-05, 5.976264e-05, 5.976259e-05, 5.976237e-05, 5.976246e-05, 
    5.976232e-05, 5.976245e-05, 5.976242e-05, 5.976231e-05, 5.976244e-05, 
    5.976216e-05, 5.976235e-05, 5.9762e-05, 5.976219e-05, 5.976199e-05, 
    5.976203e-05, 5.976197e-05, 5.976191e-05, 5.976185e-05, 5.976172e-05, 
    5.976175e-05, 5.976165e-05, 5.976271e-05, 5.976265e-05, 5.976265e-05, 
    5.976259e-05, 5.976254e-05, 5.976243e-05, 5.976226e-05, 5.976232e-05, 
    5.97622e-05, 5.976218e-05, 5.976236e-05, 5.976225e-05, 5.976261e-05, 
    5.976255e-05, 5.976258e-05, 5.976271e-05, 5.976231e-05, 5.976251e-05, 
    5.976213e-05, 5.976224e-05, 5.976192e-05, 5.976208e-05, 5.976177e-05, 
    5.976163e-05, 5.97615e-05, 5.976135e-05, 5.976261e-05, 5.976266e-05, 
    5.976258e-05, 5.976247e-05, 5.976237e-05, 5.976224e-05, 5.976222e-05, 
    5.97622e-05, 5.976213e-05, 5.976208e-05, 5.976219e-05, 5.976207e-05, 
    5.976253e-05, 5.976229e-05, 5.976267e-05, 5.976256e-05, 5.976247e-05, 
    5.976251e-05, 5.976233e-05, 5.976229e-05, 5.976211e-05, 5.97622e-05, 
    5.976166e-05, 5.97619e-05, 5.976124e-05, 5.976142e-05, 5.976267e-05, 
    5.976261e-05, 5.976241e-05, 5.97625e-05, 5.976223e-05, 5.976216e-05, 
    5.97621e-05, 5.976203e-05, 5.976203e-05, 5.976198e-05, 5.976205e-05, 
    5.976199e-05, 5.976224e-05, 5.976213e-05, 5.976243e-05, 5.976236e-05, 
    5.976239e-05, 5.976243e-05, 5.976231e-05, 5.976219e-05, 5.976219e-05, 
    5.976215e-05, 5.976203e-05, 5.976223e-05, 5.976163e-05, 5.9762e-05, 
    5.976255e-05, 5.976243e-05, 5.976242e-05, 5.976246e-05, 5.976217e-05, 
    5.976227e-05, 5.976198e-05, 5.976206e-05, 5.976194e-05, 5.9762e-05, 
    5.976201e-05, 5.976209e-05, 5.976214e-05, 5.976227e-05, 5.976237e-05, 
    5.976246e-05, 5.976244e-05, 5.976235e-05, 5.976218e-05, 5.976202e-05, 
    5.976206e-05, 5.976194e-05, 5.976225e-05, 5.976212e-05, 5.976217e-05, 
    5.976204e-05, 5.976232e-05, 5.976208e-05, 5.976238e-05, 5.976236e-05, 
    5.976227e-05, 5.976211e-05, 5.976207e-05, 5.976204e-05, 5.976206e-05, 
    5.976218e-05, 5.976219e-05, 5.976228e-05, 5.97623e-05, 5.976236e-05, 
    5.976242e-05, 5.976237e-05, 5.976232e-05, 5.976218e-05, 5.976205e-05, 
    5.976191e-05, 5.976188e-05, 5.976171e-05, 5.976185e-05, 5.976163e-05, 
    5.976182e-05, 5.97615e-05, 5.976207e-05, 5.976182e-05, 5.976227e-05, 
    5.976222e-05, 5.976214e-05, 5.976193e-05, 5.976204e-05, 5.976191e-05, 
    5.97622e-05, 5.976234e-05, 5.976238e-05, 5.976245e-05, 5.976238e-05, 
    5.976238e-05, 5.976231e-05, 5.976234e-05, 5.976217e-05, 5.976226e-05, 
    5.976201e-05, 5.976191e-05, 5.976166e-05, 5.97615e-05, 5.976133e-05, 
    5.976126e-05, 5.976124e-05, 5.976123e-05 ;

 TOTLITN =
  1.375956e-06, 1.375952e-06, 1.375953e-06, 1.375949e-06, 1.375951e-06, 
    1.375949e-06, 1.375955e-06, 1.375952e-06, 1.375954e-06, 1.375956e-06, 
    1.375943e-06, 1.375949e-06, 1.375936e-06, 1.37594e-06, 1.37593e-06, 
    1.375937e-06, 1.375929e-06, 1.37593e-06, 1.375926e-06, 1.375927e-06, 
    1.375921e-06, 1.375925e-06, 1.375918e-06, 1.375922e-06, 1.375921e-06, 
    1.375925e-06, 1.375948e-06, 1.375944e-06, 1.375948e-06, 1.375947e-06, 
    1.375948e-06, 1.375951e-06, 1.375953e-06, 1.375956e-06, 1.375956e-06, 
    1.375953e-06, 1.375947e-06, 1.375949e-06, 1.375944e-06, 1.375944e-06, 
    1.375939e-06, 1.375941e-06, 1.375932e-06, 1.375935e-06, 1.375927e-06, 
    1.375929e-06, 1.375927e-06, 1.375927e-06, 1.375927e-06, 1.37593e-06, 
    1.375929e-06, 1.375931e-06, 1.375941e-06, 1.375938e-06, 1.375946e-06, 
    1.375952e-06, 1.375955e-06, 1.375957e-06, 1.375957e-06, 1.375956e-06, 
    1.375953e-06, 1.37595e-06, 1.375948e-06, 1.375946e-06, 1.375944e-06, 
    1.37594e-06, 1.375937e-06, 1.375931e-06, 1.375932e-06, 1.375931e-06, 
    1.375929e-06, 1.375926e-06, 1.375927e-06, 1.375925e-06, 1.375931e-06, 
    1.375927e-06, 1.375933e-06, 1.375931e-06, 1.375944e-06, 1.375949e-06, 
    1.375951e-06, 1.375952e-06, 1.375957e-06, 1.375954e-06, 1.375955e-06, 
    1.375952e-06, 1.37595e-06, 1.375951e-06, 1.375946e-06, 1.375948e-06, 
    1.375937e-06, 1.375942e-06, 1.375929e-06, 1.375932e-06, 1.375928e-06, 
    1.37593e-06, 1.375927e-06, 1.37593e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.375922e-06, 1.37593e-06, 1.375927e-06, 1.375951e-06, 
    1.375951e-06, 1.375951e-06, 1.375954e-06, 1.375954e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.37595e-06, 1.375949e-06, 1.375947e-06, 
    1.375944e-06, 1.375941e-06, 1.375936e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.37593e-06, 1.375931e-06, 1.375932e-06, 1.375924e-06, 
    1.375928e-06, 1.375922e-06, 1.375922e-06, 1.375925e-06, 1.375922e-06, 
    1.375951e-06, 1.375952e-06, 1.375955e-06, 1.375953e-06, 1.375957e-06, 
    1.375954e-06, 1.375953e-06, 1.375948e-06, 1.375947e-06, 1.375946e-06, 
    1.375944e-06, 1.375941e-06, 1.375937e-06, 1.375933e-06, 1.375929e-06, 
    1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 1.375928e-06, 
    1.375927e-06, 1.375928e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375924e-06, 1.375952e-06, 1.37595e-06, 1.375951e-06, 1.37595e-06, 
    1.375951e-06, 1.375946e-06, 1.375945e-06, 1.375939e-06, 1.375941e-06, 
    1.375937e-06, 1.375941e-06, 1.37594e-06, 1.375937e-06, 1.375941e-06, 
    1.375933e-06, 1.375938e-06, 1.375928e-06, 1.375933e-06, 1.375928e-06, 
    1.375929e-06, 1.375927e-06, 1.375926e-06, 1.375924e-06, 1.37592e-06, 
    1.375921e-06, 1.375918e-06, 1.375948e-06, 1.375946e-06, 1.375947e-06, 
    1.375945e-06, 1.375943e-06, 1.37594e-06, 1.375935e-06, 1.375937e-06, 
    1.375934e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375945e-06, 
    1.375944e-06, 1.375945e-06, 1.375948e-06, 1.375937e-06, 1.375943e-06, 
    1.375932e-06, 1.375935e-06, 1.375926e-06, 1.37593e-06, 1.375922e-06, 
    1.375918e-06, 1.375914e-06, 1.37591e-06, 1.375945e-06, 1.375947e-06, 
    1.375944e-06, 1.375941e-06, 1.375939e-06, 1.375935e-06, 1.375934e-06, 
    1.375934e-06, 1.375932e-06, 1.37593e-06, 1.375933e-06, 1.37593e-06, 
    1.375943e-06, 1.375936e-06, 1.375947e-06, 1.375944e-06, 1.375942e-06, 
    1.375943e-06, 1.375937e-06, 1.375936e-06, 1.375931e-06, 1.375934e-06, 
    1.375919e-06, 1.375925e-06, 1.375907e-06, 1.375912e-06, 1.375947e-06, 
    1.375945e-06, 1.37594e-06, 1.375942e-06, 1.375935e-06, 1.375933e-06, 
    1.375931e-06, 1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 
    1.375928e-06, 1.375935e-06, 1.375932e-06, 1.37594e-06, 1.375938e-06, 
    1.375939e-06, 1.37594e-06, 1.375937e-06, 1.375933e-06, 1.375933e-06, 
    1.375932e-06, 1.375929e-06, 1.375935e-06, 1.375918e-06, 1.375928e-06, 
    1.375944e-06, 1.37594e-06, 1.37594e-06, 1.375941e-06, 1.375933e-06, 
    1.375936e-06, 1.375928e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 
    1.375928e-06, 1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375939e-06, 
    1.375941e-06, 1.375941e-06, 1.375938e-06, 1.375933e-06, 1.375929e-06, 
    1.37593e-06, 1.375927e-06, 1.375935e-06, 1.375932e-06, 1.375933e-06, 
    1.375929e-06, 1.375937e-06, 1.375931e-06, 1.375939e-06, 1.375938e-06, 
    1.375936e-06, 1.375931e-06, 1.37593e-06, 1.375929e-06, 1.37593e-06, 
    1.375933e-06, 1.375934e-06, 1.375936e-06, 1.375937e-06, 1.375938e-06, 
    1.37594e-06, 1.375938e-06, 1.375937e-06, 1.375933e-06, 1.37593e-06, 
    1.375926e-06, 1.375925e-06, 1.37592e-06, 1.375924e-06, 1.375918e-06, 
    1.375923e-06, 1.375914e-06, 1.37593e-06, 1.375923e-06, 1.375936e-06, 
    1.375935e-06, 1.375932e-06, 1.375926e-06, 1.375929e-06, 1.375926e-06, 
    1.375934e-06, 1.375938e-06, 1.375939e-06, 1.375941e-06, 1.375939e-06, 
    1.375939e-06, 1.375937e-06, 1.375938e-06, 1.375933e-06, 1.375936e-06, 
    1.375928e-06, 1.375926e-06, 1.375918e-06, 1.375914e-06, 1.375909e-06, 
    1.375907e-06, 1.375907e-06, 1.375907e-06 ;

 TOTLITN_1m =
  1.375956e-06, 1.375952e-06, 1.375953e-06, 1.375949e-06, 1.375951e-06, 
    1.375949e-06, 1.375955e-06, 1.375952e-06, 1.375954e-06, 1.375956e-06, 
    1.375943e-06, 1.375949e-06, 1.375936e-06, 1.37594e-06, 1.37593e-06, 
    1.375937e-06, 1.375929e-06, 1.37593e-06, 1.375926e-06, 1.375927e-06, 
    1.375921e-06, 1.375925e-06, 1.375918e-06, 1.375922e-06, 1.375921e-06, 
    1.375925e-06, 1.375948e-06, 1.375944e-06, 1.375948e-06, 1.375947e-06, 
    1.375948e-06, 1.375951e-06, 1.375953e-06, 1.375956e-06, 1.375956e-06, 
    1.375953e-06, 1.375947e-06, 1.375949e-06, 1.375944e-06, 1.375944e-06, 
    1.375939e-06, 1.375941e-06, 1.375932e-06, 1.375935e-06, 1.375927e-06, 
    1.375929e-06, 1.375927e-06, 1.375927e-06, 1.375927e-06, 1.37593e-06, 
    1.375929e-06, 1.375931e-06, 1.375941e-06, 1.375938e-06, 1.375946e-06, 
    1.375952e-06, 1.375955e-06, 1.375957e-06, 1.375957e-06, 1.375956e-06, 
    1.375953e-06, 1.37595e-06, 1.375948e-06, 1.375946e-06, 1.375944e-06, 
    1.37594e-06, 1.375937e-06, 1.375931e-06, 1.375932e-06, 1.375931e-06, 
    1.375929e-06, 1.375926e-06, 1.375927e-06, 1.375925e-06, 1.375931e-06, 
    1.375927e-06, 1.375933e-06, 1.375931e-06, 1.375944e-06, 1.375949e-06, 
    1.375951e-06, 1.375952e-06, 1.375957e-06, 1.375954e-06, 1.375955e-06, 
    1.375952e-06, 1.37595e-06, 1.375951e-06, 1.375946e-06, 1.375948e-06, 
    1.375937e-06, 1.375942e-06, 1.375929e-06, 1.375932e-06, 1.375928e-06, 
    1.37593e-06, 1.375927e-06, 1.37593e-06, 1.375925e-06, 1.375924e-06, 
    1.375925e-06, 1.375922e-06, 1.37593e-06, 1.375927e-06, 1.375951e-06, 
    1.375951e-06, 1.375951e-06, 1.375954e-06, 1.375954e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.37595e-06, 1.375949e-06, 1.375947e-06, 
    1.375944e-06, 1.375941e-06, 1.375936e-06, 1.375932e-06, 1.37593e-06, 
    1.375931e-06, 1.37593e-06, 1.375931e-06, 1.375932e-06, 1.375924e-06, 
    1.375928e-06, 1.375922e-06, 1.375922e-06, 1.375925e-06, 1.375922e-06, 
    1.375951e-06, 1.375952e-06, 1.375955e-06, 1.375953e-06, 1.375957e-06, 
    1.375954e-06, 1.375953e-06, 1.375948e-06, 1.375947e-06, 1.375946e-06, 
    1.375944e-06, 1.375941e-06, 1.375937e-06, 1.375933e-06, 1.375929e-06, 
    1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 1.375928e-06, 
    1.375927e-06, 1.375928e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375924e-06, 1.375952e-06, 1.37595e-06, 1.375951e-06, 1.37595e-06, 
    1.375951e-06, 1.375946e-06, 1.375945e-06, 1.375939e-06, 1.375941e-06, 
    1.375937e-06, 1.375941e-06, 1.37594e-06, 1.375937e-06, 1.375941e-06, 
    1.375933e-06, 1.375938e-06, 1.375928e-06, 1.375933e-06, 1.375928e-06, 
    1.375929e-06, 1.375927e-06, 1.375926e-06, 1.375924e-06, 1.37592e-06, 
    1.375921e-06, 1.375918e-06, 1.375948e-06, 1.375946e-06, 1.375947e-06, 
    1.375945e-06, 1.375943e-06, 1.37594e-06, 1.375935e-06, 1.375937e-06, 
    1.375934e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375945e-06, 
    1.375944e-06, 1.375945e-06, 1.375948e-06, 1.375937e-06, 1.375943e-06, 
    1.375932e-06, 1.375935e-06, 1.375926e-06, 1.37593e-06, 1.375922e-06, 
    1.375918e-06, 1.375914e-06, 1.37591e-06, 1.375945e-06, 1.375947e-06, 
    1.375944e-06, 1.375941e-06, 1.375939e-06, 1.375935e-06, 1.375934e-06, 
    1.375934e-06, 1.375932e-06, 1.37593e-06, 1.375933e-06, 1.37593e-06, 
    1.375943e-06, 1.375936e-06, 1.375947e-06, 1.375944e-06, 1.375942e-06, 
    1.375943e-06, 1.375937e-06, 1.375936e-06, 1.375931e-06, 1.375934e-06, 
    1.375919e-06, 1.375925e-06, 1.375907e-06, 1.375912e-06, 1.375947e-06, 
    1.375945e-06, 1.37594e-06, 1.375942e-06, 1.375935e-06, 1.375933e-06, 
    1.375931e-06, 1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 
    1.375928e-06, 1.375935e-06, 1.375932e-06, 1.37594e-06, 1.375938e-06, 
    1.375939e-06, 1.37594e-06, 1.375937e-06, 1.375933e-06, 1.375933e-06, 
    1.375932e-06, 1.375929e-06, 1.375935e-06, 1.375918e-06, 1.375928e-06, 
    1.375944e-06, 1.37594e-06, 1.37594e-06, 1.375941e-06, 1.375933e-06, 
    1.375936e-06, 1.375928e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 
    1.375928e-06, 1.375931e-06, 1.375932e-06, 1.375936e-06, 1.375939e-06, 
    1.375941e-06, 1.375941e-06, 1.375938e-06, 1.375933e-06, 1.375929e-06, 
    1.37593e-06, 1.375927e-06, 1.375935e-06, 1.375932e-06, 1.375933e-06, 
    1.375929e-06, 1.375937e-06, 1.375931e-06, 1.375939e-06, 1.375938e-06, 
    1.375936e-06, 1.375931e-06, 1.37593e-06, 1.375929e-06, 1.37593e-06, 
    1.375933e-06, 1.375934e-06, 1.375936e-06, 1.375937e-06, 1.375938e-06, 
    1.37594e-06, 1.375938e-06, 1.375937e-06, 1.375933e-06, 1.37593e-06, 
    1.375926e-06, 1.375925e-06, 1.37592e-06, 1.375924e-06, 1.375918e-06, 
    1.375923e-06, 1.375914e-06, 1.37593e-06, 1.375923e-06, 1.375936e-06, 
    1.375935e-06, 1.375932e-06, 1.375926e-06, 1.375929e-06, 1.375926e-06, 
    1.375934e-06, 1.375938e-06, 1.375939e-06, 1.375941e-06, 1.375939e-06, 
    1.375939e-06, 1.375937e-06, 1.375938e-06, 1.375933e-06, 1.375936e-06, 
    1.375928e-06, 1.375926e-06, 1.375918e-06, 1.375914e-06, 1.375909e-06, 
    1.375907e-06, 1.375907e-06, 1.375907e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 TOTSOMC_1m =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34476, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 TOTSOMN =
  1.773786, 1.773785, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773785, 1.773785, 1.773786, 1.773781, 1.773783, 1.773778, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773774, 1.773771, 
    1.773773, 1.773769, 1.773771, 1.773771, 1.773773, 1.773783, 1.773781, 
    1.773783, 1.773783, 1.773783, 1.773784, 1.773785, 1.773787, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773779, 1.77378, 
    1.773776, 1.773777, 1.773773, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773775, 1.773774, 1.773775, 1.77378, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773787, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773773, 1.773775, 1.773774, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773787, 1.773785, 
    1.773786, 1.773785, 1.773784, 1.773784, 1.773782, 1.773783, 1.773778, 
    1.77378, 1.773775, 1.773776, 1.773774, 1.773775, 1.773774, 1.773775, 
    1.773773, 1.773772, 1.773772, 1.773771, 1.773775, 1.773774, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773787, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773783, 1.773781, 1.77378, 1.773777, 1.773776, 
    1.773775, 1.773775, 1.773775, 1.773775, 1.773776, 1.773772, 1.773774, 
    1.773771, 1.773772, 1.773773, 1.773772, 1.773784, 1.773785, 1.773786, 
    1.773785, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773776, 1.773774, 1.773775, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773774, 1.773774, 1.773772, 1.773772, 
    1.773772, 1.773772, 1.773785, 1.773784, 1.773784, 1.773784, 1.773784, 
    1.773782, 1.773781, 1.773779, 1.77378, 1.773778, 1.77378, 1.773779, 
    1.773778, 1.77378, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773774, 1.773773, 1.773772, 1.773771, 1.773771, 1.77377, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.773781, 1.773779, 1.773777, 
    1.773778, 1.773777, 1.773776, 1.773779, 1.773777, 1.773782, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773776, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773768, 1.773766, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773779, 1.773777, 1.773777, 1.773777, 1.773776, 
    1.773775, 1.773776, 1.773775, 1.773781, 1.773778, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773778, 1.773775, 1.773777, 1.77377, 
    1.773773, 1.773765, 1.773767, 1.773782, 1.773782, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773775, 
    1.773774, 1.773777, 1.773776, 1.773779, 1.773779, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.77378, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773776, 
    1.773777, 1.773779, 1.77378, 1.77378, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773776, 1.773776, 1.773775, 1.773778, 
    1.773775, 1.773779, 1.773779, 1.773777, 1.773775, 1.773775, 1.773775, 
    1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 1.773779, 
    1.773779, 1.773778, 1.773776, 1.773775, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773772, 1.773768, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773776, 1.773773, 1.773775, 1.773773, 1.773777, 1.773778, 
    1.773779, 1.77378, 1.773779, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.77377, 1.773768, 1.773766, 1.773765, 
    1.773764, 1.773764 ;

 TOTSOMN_1m =
  1.773786, 1.773785, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773785, 1.773785, 1.773786, 1.773781, 1.773783, 1.773778, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773774, 1.773771, 
    1.773773, 1.773769, 1.773771, 1.773771, 1.773773, 1.773783, 1.773781, 
    1.773783, 1.773783, 1.773783, 1.773784, 1.773785, 1.773787, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773779, 1.77378, 
    1.773776, 1.773777, 1.773773, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773775, 1.773774, 1.773775, 1.77378, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773787, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773773, 1.773775, 1.773774, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773787, 1.773785, 
    1.773786, 1.773785, 1.773784, 1.773784, 1.773782, 1.773783, 1.773778, 
    1.77378, 1.773775, 1.773776, 1.773774, 1.773775, 1.773774, 1.773775, 
    1.773773, 1.773772, 1.773772, 1.773771, 1.773775, 1.773774, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773787, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773783, 1.773781, 1.77378, 1.773777, 1.773776, 
    1.773775, 1.773775, 1.773775, 1.773775, 1.773776, 1.773772, 1.773774, 
    1.773771, 1.773772, 1.773773, 1.773772, 1.773784, 1.773785, 1.773786, 
    1.773785, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773776, 1.773774, 1.773775, 1.773775, 
    1.773774, 1.773775, 1.773774, 1.773774, 1.773774, 1.773772, 1.773772, 
    1.773772, 1.773772, 1.773785, 1.773784, 1.773784, 1.773784, 1.773784, 
    1.773782, 1.773781, 1.773779, 1.77378, 1.773778, 1.77378, 1.773779, 
    1.773778, 1.77378, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773774, 1.773773, 1.773772, 1.773771, 1.773771, 1.77377, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.773781, 1.773779, 1.773777, 
    1.773778, 1.773777, 1.773776, 1.773779, 1.773777, 1.773782, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773776, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773768, 1.773766, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773779, 1.773777, 1.773777, 1.773777, 1.773776, 
    1.773775, 1.773776, 1.773775, 1.773781, 1.773778, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773778, 1.773775, 1.773777, 1.77377, 
    1.773773, 1.773765, 1.773767, 1.773782, 1.773782, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773775, 
    1.773774, 1.773777, 1.773776, 1.773779, 1.773779, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.77378, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773776, 
    1.773777, 1.773779, 1.77378, 1.77378, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773776, 1.773776, 1.773775, 1.773778, 
    1.773775, 1.773779, 1.773779, 1.773777, 1.773775, 1.773775, 1.773775, 
    1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 1.773779, 
    1.773779, 1.773778, 1.773776, 1.773775, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773772, 1.773768, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773776, 1.773773, 1.773775, 1.773773, 1.773777, 1.773778, 
    1.773779, 1.77378, 1.773779, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.77377, 1.773768, 1.773766, 1.773765, 
    1.773764, 1.773764 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9694, 249.9697, 249.9697, 249.9699, 249.9697, 249.9699, 249.9695, 
    249.9697, 249.9696, 249.9695, 249.9702, 249.9699, 249.9707, 249.9704, 
    249.9711, 249.9706, 249.9711, 249.9711, 249.9713, 249.9713, 249.9716, 
    249.9714, 249.9718, 249.9716, 249.9716, 249.9714, 249.97, 249.9702, 
    249.9699, 249.97, 249.97, 249.9697, 249.9696, 249.9694, 249.9695, 
    249.9696, 249.97, 249.9699, 249.9702, 249.9702, 249.9705, 249.9704, 
    249.9709, 249.9708, 249.9713, 249.9711, 249.9713, 249.9712, 249.9713, 
    249.9711, 249.9712, 249.971, 249.9704, 249.9706, 249.97, 249.9697, 
    249.9695, 249.9694, 249.9694, 249.9694, 249.9696, 249.9698, 249.97, 
    249.9701, 249.9702, 249.9705, 249.9706, 249.971, 249.9709, 249.971, 
    249.9711, 249.9713, 249.9713, 249.9714, 249.971, 249.9712, 249.9709, 
    249.971, 249.9702, 249.9699, 249.9698, 249.9697, 249.9694, 249.9696, 
    249.9695, 249.9697, 249.9698, 249.9697, 249.9701, 249.9699, 249.9706, 
    249.9703, 249.9711, 249.9709, 249.9712, 249.971, 249.9713, 249.9711, 
    249.9714, 249.9715, 249.9714, 249.9716, 249.9711, 249.9713, 249.9697, 
    249.9697, 249.9698, 249.9696, 249.9696, 249.9694, 249.9696, 249.9696, 
    249.9698, 249.9699, 249.97, 249.9702, 249.9704, 249.9707, 249.9709, 
    249.9711, 249.971, 249.9711, 249.971, 249.9709, 249.9714, 249.9712, 
    249.9716, 249.9715, 249.9714, 249.9715, 249.9698, 249.9697, 249.9695, 
    249.9697, 249.9694, 249.9695, 249.9696, 249.9699, 249.97, 249.9701, 
    249.9702, 249.9704, 249.9707, 249.9709, 249.9711, 249.9711, 249.9711, 
    249.9712, 249.9711, 249.9712, 249.9712, 249.9712, 249.9715, 249.9714, 
    249.9715, 249.9715, 249.9697, 249.9698, 249.9698, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9705, 249.9704, 249.9706, 249.9704, 249.9704, 
    249.9706, 249.9704, 249.9709, 249.9706, 249.9712, 249.9708, 249.9712, 
    249.9711, 249.9712, 249.9713, 249.9715, 249.9717, 249.9716, 249.9718, 
    249.9699, 249.97, 249.97, 249.9702, 249.9702, 249.9704, 249.9707, 
    249.9706, 249.9708, 249.9709, 249.9706, 249.9707, 249.9701, 249.9702, 
    249.9702, 249.9699, 249.9706, 249.9703, 249.9709, 249.9707, 249.9713, 
    249.971, 249.9716, 249.9718, 249.9721, 249.9723, 249.9701, 249.97, 
    249.9702, 249.9704, 249.9705, 249.9708, 249.9708, 249.9708, 249.9709, 
    249.971, 249.9708, 249.9711, 249.9702, 249.9707, 249.97, 249.9702, 
    249.9703, 249.9703, 249.9706, 249.9707, 249.971, 249.9708, 249.9718, 
    249.9714, 249.9725, 249.9722, 249.97, 249.9701, 249.9705, 249.9703, 
    249.9708, 249.9709, 249.971, 249.9711, 249.9711, 249.9712, 249.9711, 
    249.9712, 249.9708, 249.971, 249.9704, 249.9706, 249.9705, 249.9704, 
    249.9706, 249.9708, 249.9709, 249.9709, 249.9711, 249.9708, 249.9718, 
    249.9712, 249.9702, 249.9704, 249.9704, 249.9704, 249.9709, 249.9707, 
    249.9712, 249.9711, 249.9713, 249.9712, 249.9712, 249.971, 249.9709, 
    249.9707, 249.9705, 249.9704, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9711, 249.9713, 249.9707, 249.971, 249.9709, 249.9711, 249.9706, 
    249.971, 249.9705, 249.9706, 249.9707, 249.971, 249.9711, 249.9711, 
    249.9711, 249.9709, 249.9708, 249.9707, 249.9706, 249.9705, 249.9704, 
    249.9705, 249.9706, 249.9709, 249.9711, 249.9713, 249.9714, 249.9717, 
    249.9715, 249.9718, 249.9715, 249.9721, 249.9711, 249.9715, 249.9707, 
    249.9708, 249.9709, 249.9713, 249.9711, 249.9713, 249.9708, 249.9706, 
    249.9705, 249.9704, 249.9705, 249.9705, 249.9706, 249.9706, 249.9709, 
    249.9707, 249.9712, 249.9713, 249.9718, 249.9721, 249.9724, 249.9725, 
    249.9725, 249.9725 ;

 TREFMNAV_R =
  249.9694, 249.9697, 249.9697, 249.9699, 249.9697, 249.9699, 249.9695, 
    249.9697, 249.9696, 249.9695, 249.9702, 249.9699, 249.9707, 249.9704, 
    249.9711, 249.9706, 249.9711, 249.9711, 249.9713, 249.9713, 249.9716, 
    249.9714, 249.9718, 249.9716, 249.9716, 249.9714, 249.97, 249.9702, 
    249.9699, 249.97, 249.97, 249.9697, 249.9696, 249.9694, 249.9695, 
    249.9696, 249.97, 249.9699, 249.9702, 249.9702, 249.9705, 249.9704, 
    249.9709, 249.9708, 249.9713, 249.9711, 249.9713, 249.9712, 249.9713, 
    249.9711, 249.9712, 249.971, 249.9704, 249.9706, 249.97, 249.9697, 
    249.9695, 249.9694, 249.9694, 249.9694, 249.9696, 249.9698, 249.97, 
    249.9701, 249.9702, 249.9705, 249.9706, 249.971, 249.9709, 249.971, 
    249.9711, 249.9713, 249.9713, 249.9714, 249.971, 249.9712, 249.9709, 
    249.971, 249.9702, 249.9699, 249.9698, 249.9697, 249.9694, 249.9696, 
    249.9695, 249.9697, 249.9698, 249.9697, 249.9701, 249.9699, 249.9706, 
    249.9703, 249.9711, 249.9709, 249.9712, 249.971, 249.9713, 249.9711, 
    249.9714, 249.9715, 249.9714, 249.9716, 249.9711, 249.9713, 249.9697, 
    249.9697, 249.9698, 249.9696, 249.9696, 249.9694, 249.9696, 249.9696, 
    249.9698, 249.9699, 249.97, 249.9702, 249.9704, 249.9707, 249.9709, 
    249.9711, 249.971, 249.9711, 249.971, 249.9709, 249.9714, 249.9712, 
    249.9716, 249.9715, 249.9714, 249.9715, 249.9698, 249.9697, 249.9695, 
    249.9697, 249.9694, 249.9695, 249.9696, 249.9699, 249.97, 249.9701, 
    249.9702, 249.9704, 249.9707, 249.9709, 249.9711, 249.9711, 249.9711, 
    249.9712, 249.9711, 249.9712, 249.9712, 249.9712, 249.9715, 249.9714, 
    249.9715, 249.9715, 249.9697, 249.9698, 249.9698, 249.9698, 249.9698, 
    249.97, 249.9701, 249.9705, 249.9704, 249.9706, 249.9704, 249.9704, 
    249.9706, 249.9704, 249.9709, 249.9706, 249.9712, 249.9708, 249.9712, 
    249.9711, 249.9712, 249.9713, 249.9715, 249.9717, 249.9716, 249.9718, 
    249.9699, 249.97, 249.97, 249.9702, 249.9702, 249.9704, 249.9707, 
    249.9706, 249.9708, 249.9709, 249.9706, 249.9707, 249.9701, 249.9702, 
    249.9702, 249.9699, 249.9706, 249.9703, 249.9709, 249.9707, 249.9713, 
    249.971, 249.9716, 249.9718, 249.9721, 249.9723, 249.9701, 249.97, 
    249.9702, 249.9704, 249.9705, 249.9708, 249.9708, 249.9708, 249.9709, 
    249.971, 249.9708, 249.9711, 249.9702, 249.9707, 249.97, 249.9702, 
    249.9703, 249.9703, 249.9706, 249.9707, 249.971, 249.9708, 249.9718, 
    249.9714, 249.9725, 249.9722, 249.97, 249.9701, 249.9705, 249.9703, 
    249.9708, 249.9709, 249.971, 249.9711, 249.9711, 249.9712, 249.9711, 
    249.9712, 249.9708, 249.971, 249.9704, 249.9706, 249.9705, 249.9704, 
    249.9706, 249.9708, 249.9709, 249.9709, 249.9711, 249.9708, 249.9718, 
    249.9712, 249.9702, 249.9704, 249.9704, 249.9704, 249.9709, 249.9707, 
    249.9712, 249.9711, 249.9713, 249.9712, 249.9712, 249.971, 249.9709, 
    249.9707, 249.9705, 249.9704, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9711, 249.9713, 249.9707, 249.971, 249.9709, 249.9711, 249.9706, 
    249.971, 249.9705, 249.9706, 249.9707, 249.971, 249.9711, 249.9711, 
    249.9711, 249.9709, 249.9708, 249.9707, 249.9706, 249.9705, 249.9704, 
    249.9705, 249.9706, 249.9709, 249.9711, 249.9713, 249.9714, 249.9717, 
    249.9715, 249.9718, 249.9715, 249.9721, 249.9711, 249.9715, 249.9707, 
    249.9708, 249.9709, 249.9713, 249.9711, 249.9713, 249.9708, 249.9706, 
    249.9705, 249.9704, 249.9705, 249.9705, 249.9706, 249.9706, 249.9709, 
    249.9707, 249.9712, 249.9713, 249.9718, 249.9721, 249.9724, 249.9725, 
    249.9725, 249.9725 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.516, 258.5164, 258.5163, 258.5167, 258.5165, 258.5167, 258.5161, 
    258.5164, 258.5162, 258.5161, 258.5173, 258.5167, 258.5179, 258.5175, 
    258.5185, 258.5179, 258.5187, 258.5185, 258.519, 258.5189, 258.5194, 
    258.519, 258.5197, 258.5193, 258.5194, 258.519, 258.5168, 258.5172, 
    258.5168, 258.5168, 258.5168, 258.5165, 258.5163, 258.516, 258.5161, 
    258.5163, 258.5169, 258.5167, 258.5172, 258.5172, 258.5177, 258.5175, 
    258.5184, 258.5181, 258.5189, 258.5187, 258.5189, 258.5188, 258.5189, 
    258.5186, 258.5187, 258.5185, 258.5175, 258.5178, 258.5169, 258.5164, 
    258.5161, 258.5159, 258.5159, 258.516, 258.5163, 258.5166, 258.5168, 
    258.517, 258.5172, 258.5176, 258.5179, 258.5184, 258.5183, 258.5185, 
    258.5186, 258.5189, 258.5189, 258.519, 258.5185, 258.5188, 258.5183, 
    258.5184, 258.5172, 258.5167, 258.5165, 258.5164, 258.5159, 258.5162, 
    258.5161, 258.5164, 258.5166, 258.5165, 258.517, 258.5168, 258.5179, 
    258.5174, 258.5186, 258.5183, 258.5187, 258.5185, 258.5188, 258.5186, 
    258.519, 258.5192, 258.5191, 258.5194, 258.5185, 258.5189, 258.5165, 
    258.5165, 258.5165, 258.5163, 258.5162, 258.516, 258.5162, 258.5163, 
    258.5166, 258.5167, 258.5168, 258.5172, 258.5175, 258.518, 258.5184, 
    258.5186, 258.5185, 258.5186, 258.5184, 258.5184, 258.5191, 258.5187, 
    258.5193, 258.5193, 258.519, 258.5193, 258.5165, 258.5164, 258.5161, 
    258.5164, 258.516, 258.5162, 258.5163, 258.5168, 258.5169, 258.517, 
    258.5172, 258.5175, 258.5179, 258.5183, 258.5187, 258.5186, 258.5186, 
    258.5187, 258.5185, 258.5188, 258.5188, 258.5187, 258.5193, 258.5191, 
    258.5193, 258.5192, 258.5164, 258.5166, 258.5165, 258.5166, 258.5165, 
    258.517, 258.5171, 258.5177, 258.5175, 258.5179, 258.5175, 258.5175, 
    258.5179, 258.5175, 258.5183, 258.5178, 258.5187, 258.5182, 258.5188, 
    258.5187, 258.5188, 258.519, 258.5192, 258.5195, 258.5194, 258.5197, 
    258.5168, 258.5169, 258.5169, 258.5171, 258.5172, 258.5175, 258.518, 
    258.5179, 258.5182, 258.5182, 258.5177, 258.518, 258.5171, 258.5172, 
    258.5171, 258.5168, 258.5179, 258.5173, 258.5184, 258.5181, 258.519, 
    258.5185, 258.5194, 258.5197, 258.5201, 258.5205, 258.5171, 258.5169, 
    258.5172, 258.5174, 258.5177, 258.5181, 258.5181, 258.5182, 258.5184, 
    258.5185, 258.5182, 258.5186, 258.5172, 258.5179, 258.5169, 258.5172, 
    258.5174, 258.5173, 258.5178, 258.5179, 258.5184, 258.5182, 258.5197, 
    258.519, 258.5208, 258.5203, 258.5169, 258.5171, 258.5176, 258.5173, 
    258.5181, 258.5183, 258.5184, 258.5186, 258.5186, 258.5188, 258.5186, 
    258.5188, 258.5181, 258.5184, 258.5175, 258.5178, 258.5177, 258.5175, 
    258.5179, 258.5182, 258.5182, 258.5183, 258.5186, 258.5181, 258.5197, 
    258.5187, 258.5172, 258.5175, 258.5176, 258.5175, 258.5183, 258.518, 
    258.5188, 258.5186, 258.5189, 258.5187, 258.5187, 258.5185, 258.5183, 
    258.518, 258.5177, 258.5175, 258.5175, 258.5178, 258.5182, 258.5186, 
    258.5186, 258.5189, 258.518, 258.5184, 258.5182, 258.5186, 258.5179, 
    258.5185, 258.5177, 258.5178, 258.518, 258.5184, 258.5185, 258.5186, 
    258.5186, 258.5182, 258.5182, 258.518, 258.5179, 258.5177, 258.5176, 
    258.5177, 258.5179, 258.5182, 258.5186, 258.519, 258.5191, 258.5195, 
    258.5191, 258.5197, 258.5192, 258.5201, 258.5185, 258.5192, 258.518, 
    258.5181, 258.5183, 258.5189, 258.5186, 258.519, 258.5182, 258.5178, 
    258.5177, 258.5175, 258.5177, 258.5177, 258.5179, 258.5178, 258.5182, 
    258.518, 258.5187, 258.519, 258.5197, 258.5201, 258.5206, 258.5208, 
    258.5208, 258.5209 ;

 TREFMXAV_R =
  258.516, 258.5164, 258.5163, 258.5167, 258.5165, 258.5167, 258.5161, 
    258.5164, 258.5162, 258.5161, 258.5173, 258.5167, 258.5179, 258.5175, 
    258.5185, 258.5179, 258.5187, 258.5185, 258.519, 258.5189, 258.5194, 
    258.519, 258.5197, 258.5193, 258.5194, 258.519, 258.5168, 258.5172, 
    258.5168, 258.5168, 258.5168, 258.5165, 258.5163, 258.516, 258.5161, 
    258.5163, 258.5169, 258.5167, 258.5172, 258.5172, 258.5177, 258.5175, 
    258.5184, 258.5181, 258.5189, 258.5187, 258.5189, 258.5188, 258.5189, 
    258.5186, 258.5187, 258.5185, 258.5175, 258.5178, 258.5169, 258.5164, 
    258.5161, 258.5159, 258.5159, 258.516, 258.5163, 258.5166, 258.5168, 
    258.517, 258.5172, 258.5176, 258.5179, 258.5184, 258.5183, 258.5185, 
    258.5186, 258.5189, 258.5189, 258.519, 258.5185, 258.5188, 258.5183, 
    258.5184, 258.5172, 258.5167, 258.5165, 258.5164, 258.5159, 258.5162, 
    258.5161, 258.5164, 258.5166, 258.5165, 258.517, 258.5168, 258.5179, 
    258.5174, 258.5186, 258.5183, 258.5187, 258.5185, 258.5188, 258.5186, 
    258.519, 258.5192, 258.5191, 258.5194, 258.5185, 258.5189, 258.5165, 
    258.5165, 258.5165, 258.5163, 258.5162, 258.516, 258.5162, 258.5163, 
    258.5166, 258.5167, 258.5168, 258.5172, 258.5175, 258.518, 258.5184, 
    258.5186, 258.5185, 258.5186, 258.5184, 258.5184, 258.5191, 258.5187, 
    258.5193, 258.5193, 258.519, 258.5193, 258.5165, 258.5164, 258.5161, 
    258.5164, 258.516, 258.5162, 258.5163, 258.5168, 258.5169, 258.517, 
    258.5172, 258.5175, 258.5179, 258.5183, 258.5187, 258.5186, 258.5186, 
    258.5187, 258.5185, 258.5188, 258.5188, 258.5187, 258.5193, 258.5191, 
    258.5193, 258.5192, 258.5164, 258.5166, 258.5165, 258.5166, 258.5165, 
    258.517, 258.5171, 258.5177, 258.5175, 258.5179, 258.5175, 258.5175, 
    258.5179, 258.5175, 258.5183, 258.5178, 258.5187, 258.5182, 258.5188, 
    258.5187, 258.5188, 258.519, 258.5192, 258.5195, 258.5194, 258.5197, 
    258.5168, 258.5169, 258.5169, 258.5171, 258.5172, 258.5175, 258.518, 
    258.5179, 258.5182, 258.5182, 258.5177, 258.518, 258.5171, 258.5172, 
    258.5171, 258.5168, 258.5179, 258.5173, 258.5184, 258.5181, 258.519, 
    258.5185, 258.5194, 258.5197, 258.5201, 258.5205, 258.5171, 258.5169, 
    258.5172, 258.5174, 258.5177, 258.5181, 258.5181, 258.5182, 258.5184, 
    258.5185, 258.5182, 258.5186, 258.5172, 258.5179, 258.5169, 258.5172, 
    258.5174, 258.5173, 258.5178, 258.5179, 258.5184, 258.5182, 258.5197, 
    258.519, 258.5208, 258.5203, 258.5169, 258.5171, 258.5176, 258.5173, 
    258.5181, 258.5183, 258.5184, 258.5186, 258.5186, 258.5188, 258.5186, 
    258.5188, 258.5181, 258.5184, 258.5175, 258.5178, 258.5177, 258.5175, 
    258.5179, 258.5182, 258.5182, 258.5183, 258.5186, 258.5181, 258.5197, 
    258.5187, 258.5172, 258.5175, 258.5176, 258.5175, 258.5183, 258.518, 
    258.5188, 258.5186, 258.5189, 258.5187, 258.5187, 258.5185, 258.5183, 
    258.518, 258.5177, 258.5175, 258.5175, 258.5178, 258.5182, 258.5186, 
    258.5186, 258.5189, 258.518, 258.5184, 258.5182, 258.5186, 258.5179, 
    258.5185, 258.5177, 258.5178, 258.518, 258.5184, 258.5185, 258.5186, 
    258.5186, 258.5182, 258.5182, 258.518, 258.5179, 258.5177, 258.5176, 
    258.5177, 258.5179, 258.5182, 258.5186, 258.519, 258.5191, 258.5195, 
    258.5191, 258.5197, 258.5192, 258.5201, 258.5185, 258.5192, 258.518, 
    258.5181, 258.5183, 258.5189, 258.5186, 258.519, 258.5182, 258.5178, 
    258.5177, 258.5175, 258.5177, 258.5177, 258.5179, 258.5178, 258.5182, 
    258.518, 258.5187, 258.519, 258.5197, 258.5201, 258.5206, 258.5208, 
    258.5208, 258.5209 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9562, 253.9564, 253.9563, 253.9565, 253.9564, 253.9565, 253.9562, 
    253.9564, 253.9563, 253.9562, 253.9567, 253.9565, 253.957, 253.9568, 
    253.9573, 253.957, 253.9573, 253.9573, 253.9575, 253.9574, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.9577, 253.9575, 253.9565, 253.9567, 
    253.9565, 253.9565, 253.9565, 253.9564, 253.9563, 253.9562, 253.9562, 
    253.9563, 253.9566, 253.9565, 253.9567, 253.9567, 253.9569, 253.9568, 
    253.9572, 253.9571, 253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 
    253.9573, 253.9574, 253.9572, 253.9568, 253.957, 253.9566, 253.9564, 
    253.9562, 253.9561, 253.9561, 253.9562, 253.9563, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.9569, 253.957, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9574, 253.9575, 253.9573, 253.9574, 253.9572, 
    253.9572, 253.9567, 253.9565, 253.9564, 253.9563, 253.9562, 253.9563, 
    253.9562, 253.9564, 253.9564, 253.9564, 253.9566, 253.9565, 253.957, 
    253.9568, 253.9573, 253.9572, 253.9574, 253.9573, 253.9574, 253.9573, 
    253.9575, 253.9575, 253.9575, 253.9576, 253.9573, 253.9574, 253.9564, 
    253.9564, 253.9564, 253.9563, 253.9563, 253.9562, 253.9563, 253.9563, 
    253.9564, 253.9565, 253.9566, 253.9567, 253.9568, 253.957, 253.9572, 
    253.9573, 253.9572, 253.9573, 253.9572, 253.9572, 253.9575, 253.9574, 
    253.9576, 253.9576, 253.9575, 253.9576, 253.9564, 253.9564, 253.9563, 
    253.9563, 253.9562, 253.9563, 253.9563, 253.9565, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9572, 253.9573, 253.9573, 253.9573, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9576, 253.9575, 
    253.9576, 253.9576, 253.9564, 253.9564, 253.9564, 253.9565, 253.9564, 
    253.9566, 253.9567, 253.9569, 253.9568, 253.957, 253.9568, 253.9569, 
    253.957, 253.9568, 253.9572, 253.9569, 253.9574, 253.9571, 253.9574, 
    253.9573, 253.9574, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9565, 253.9566, 253.9566, 253.9567, 253.9567, 253.9568, 253.9571, 
    253.957, 253.9571, 253.9572, 253.9569, 253.9571, 253.9566, 253.9567, 
    253.9567, 253.9565, 253.957, 253.9568, 253.9572, 253.9571, 253.9575, 
    253.9573, 253.9576, 253.9578, 253.958, 253.9581, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.9569, 253.9571, 253.9571, 253.9571, 253.9572, 
    253.9573, 253.9571, 253.9573, 253.9567, 253.957, 253.9566, 253.9567, 
    253.9568, 253.9568, 253.957, 253.957, 253.9572, 253.9571, 253.9578, 
    253.9575, 253.9583, 253.958, 253.9566, 253.9566, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9572, 253.9573, 253.9573, 253.9574, 253.9573, 
    253.9574, 253.9571, 253.9572, 253.9568, 253.9569, 253.9569, 253.9568, 
    253.957, 253.9571, 253.9571, 253.9572, 253.9573, 253.9571, 253.9578, 
    253.9574, 253.9567, 253.9568, 253.9569, 253.9568, 253.9572, 253.957, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.957, 253.9569, 253.9568, 253.9568, 253.957, 253.9571, 253.9573, 
    253.9573, 253.9574, 253.9571, 253.9572, 253.9572, 253.9573, 253.957, 
    253.9572, 253.9569, 253.9569, 253.957, 253.9572, 253.9573, 253.9573, 
    253.9573, 253.9572, 253.9571, 253.957, 253.957, 253.9569, 253.9569, 
    253.9569, 253.957, 253.9572, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.957, 
    253.9571, 253.9572, 253.9574, 253.9573, 253.9575, 253.9571, 253.957, 
    253.9569, 253.9568, 253.9569, 253.9569, 253.957, 253.957, 253.9572, 
    253.957, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9562, 253.9564, 253.9563, 253.9565, 253.9564, 253.9565, 253.9562, 
    253.9564, 253.9563, 253.9562, 253.9567, 253.9565, 253.957, 253.9568, 
    253.9573, 253.957, 253.9573, 253.9573, 253.9575, 253.9574, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.9577, 253.9575, 253.9565, 253.9567, 
    253.9565, 253.9565, 253.9565, 253.9564, 253.9563, 253.9562, 253.9562, 
    253.9563, 253.9566, 253.9565, 253.9567, 253.9567, 253.9569, 253.9568, 
    253.9572, 253.9571, 253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 
    253.9573, 253.9574, 253.9572, 253.9568, 253.957, 253.9566, 253.9564, 
    253.9562, 253.9561, 253.9561, 253.9562, 253.9563, 253.9565, 253.9565, 
    253.9566, 253.9567, 253.9569, 253.957, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9574, 253.9575, 253.9573, 253.9574, 253.9572, 
    253.9572, 253.9567, 253.9565, 253.9564, 253.9563, 253.9562, 253.9563, 
    253.9562, 253.9564, 253.9564, 253.9564, 253.9566, 253.9565, 253.957, 
    253.9568, 253.9573, 253.9572, 253.9574, 253.9573, 253.9574, 253.9573, 
    253.9575, 253.9575, 253.9575, 253.9576, 253.9573, 253.9574, 253.9564, 
    253.9564, 253.9564, 253.9563, 253.9563, 253.9562, 253.9563, 253.9563, 
    253.9564, 253.9565, 253.9566, 253.9567, 253.9568, 253.957, 253.9572, 
    253.9573, 253.9572, 253.9573, 253.9572, 253.9572, 253.9575, 253.9574, 
    253.9576, 253.9576, 253.9575, 253.9576, 253.9564, 253.9564, 253.9563, 
    253.9563, 253.9562, 253.9563, 253.9563, 253.9565, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9572, 253.9573, 253.9573, 253.9573, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9576, 253.9575, 
    253.9576, 253.9576, 253.9564, 253.9564, 253.9564, 253.9565, 253.9564, 
    253.9566, 253.9567, 253.9569, 253.9568, 253.957, 253.9568, 253.9569, 
    253.957, 253.9568, 253.9572, 253.9569, 253.9574, 253.9571, 253.9574, 
    253.9573, 253.9574, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9565, 253.9566, 253.9566, 253.9567, 253.9567, 253.9568, 253.9571, 
    253.957, 253.9571, 253.9572, 253.9569, 253.9571, 253.9566, 253.9567, 
    253.9567, 253.9565, 253.957, 253.9568, 253.9572, 253.9571, 253.9575, 
    253.9573, 253.9576, 253.9578, 253.958, 253.9581, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.9569, 253.9571, 253.9571, 253.9571, 253.9572, 
    253.9573, 253.9571, 253.9573, 253.9567, 253.957, 253.9566, 253.9567, 
    253.9568, 253.9568, 253.957, 253.957, 253.9572, 253.9571, 253.9578, 
    253.9575, 253.9583, 253.958, 253.9566, 253.9566, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9572, 253.9573, 253.9573, 253.9574, 253.9573, 
    253.9574, 253.9571, 253.9572, 253.9568, 253.9569, 253.9569, 253.9568, 
    253.957, 253.9571, 253.9571, 253.9572, 253.9573, 253.9571, 253.9578, 
    253.9574, 253.9567, 253.9568, 253.9569, 253.9568, 253.9572, 253.957, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.957, 253.9569, 253.9568, 253.9568, 253.957, 253.9571, 253.9573, 
    253.9573, 253.9574, 253.9571, 253.9572, 253.9572, 253.9573, 253.957, 
    253.9572, 253.9569, 253.9569, 253.957, 253.9572, 253.9573, 253.9573, 
    253.9573, 253.9572, 253.9571, 253.957, 253.957, 253.9569, 253.9569, 
    253.9569, 253.957, 253.9572, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.957, 
    253.9571, 253.9572, 253.9574, 253.9573, 253.9575, 253.9571, 253.957, 
    253.9569, 253.9568, 253.9569, 253.9569, 253.957, 253.957, 253.9572, 
    253.957, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.3909, 254.3923, 254.392, 254.3932, 254.3926, 254.3933, 254.3912, 
    254.3924, 254.3916, 254.391, 254.3954, 254.3932, 254.3977, 254.3963, 
    254.3999, 254.3975, 254.4003, 254.3998, 254.4015, 254.401, 254.4031, 
    254.4017, 254.4042, 254.4028, 254.403, 254.4016, 254.3937, 254.3951, 
    254.3936, 254.3938, 254.3937, 254.3926, 254.392, 254.3908, 254.391, 
    254.3919, 254.3939, 254.3932, 254.395, 254.3949, 254.3969, 254.396, 
    254.3993, 254.3983, 254.401, 254.4003, 254.401, 254.4008, 254.401, 254.4, 
    254.4004, 254.3996, 254.3961, 254.3971, 254.3942, 254.3924, 254.3912, 
    254.3904, 254.3905, 254.3907, 254.3919, 254.393, 254.3938, 254.3944, 
    254.3949, 254.3965, 254.3974, 254.3994, 254.3991, 254.3997, 254.4003, 
    254.4012, 254.4011, 254.4015, 254.3997, 254.4009, 254.3989, 254.3994, 
    254.395, 254.3934, 254.3927, 254.3921, 254.3906, 254.3916, 254.3912, 
    254.3922, 254.3928, 254.3925, 254.3944, 254.3937, 254.3975, 254.3958, 
    254.4002, 254.3992, 254.4005, 254.3998, 254.4009, 254.3999, 254.4017, 
    254.4021, 254.4018, 254.4028, 254.3999, 254.401, 254.3925, 254.3926, 
    254.3928, 254.3918, 254.3917, 254.3908, 254.3916, 254.392, 254.3929, 
    254.3934, 254.3939, 254.395, 254.3962, 254.398, 254.3992, 254.4001, 
    254.3996, 254.4, 254.3995, 254.3993, 254.4019, 254.4004, 254.4027, 
    254.4026, 254.4015, 254.4026, 254.3926, 254.3923, 254.3913, 254.3921, 
    254.3907, 254.3915, 254.3919, 254.3937, 254.3941, 254.3944, 254.3951, 
    254.396, 254.3976, 254.399, 254.4003, 254.4002, 254.4003, 254.4005, 
    254.3998, 254.4007, 254.4008, 254.4004, 254.4025, 254.4019, 254.4025, 
    254.4022, 254.3924, 254.3929, 254.3926, 254.3931, 254.3928, 254.3943, 
    254.3947, 254.3969, 254.396, 254.3974, 254.3962, 254.3964, 254.3974, 
    254.3962, 254.3989, 254.3971, 254.4005, 254.3986, 254.4007, 254.4003, 
    254.4009, 254.4014, 254.4021, 254.4033, 254.403, 254.4041, 254.3936, 
    254.3942, 254.3942, 254.3948, 254.3953, 254.3963, 254.398, 254.3974, 
    254.3986, 254.3988, 254.397, 254.3981, 254.3946, 254.3952, 254.3949, 
    254.3936, 254.3975, 254.3955, 254.3992, 254.3982, 254.4014, 254.3997, 
    254.4029, 254.4042, 254.4055, 254.4069, 254.3946, 254.3941, 254.3949, 
    254.3959, 254.3969, 254.3982, 254.3984, 254.3986, 254.3992, 254.3998, 
    254.3987, 254.3999, 254.3952, 254.3977, 254.394, 254.3951, 254.3959, 
    254.3955, 254.3973, 254.3978, 254.3995, 254.3986, 254.4038, 254.4015, 
    254.4081, 254.4062, 254.394, 254.3946, 254.3965, 254.3956, 254.3983, 
    254.399, 254.3995, 254.4002, 254.4003, 254.4007, 254.4, 254.4007, 
    254.3982, 254.3993, 254.3963, 254.397, 254.3967, 254.3963, 254.3975, 
    254.3987, 254.3987, 254.3991, 254.4001, 254.3983, 254.4041, 254.4005, 
    254.3952, 254.3962, 254.3964, 254.396, 254.3989, 254.3979, 254.4007, 
    254.3999, 254.4012, 254.4006, 254.4005, 254.3997, 254.3992, 254.3979, 
    254.3969, 254.3961, 254.3963, 254.3971, 254.3988, 254.4003, 254.4, 
    254.4011, 254.3981, 254.3994, 254.3989, 254.4001, 254.3974, 254.3996, 
    254.3968, 254.397, 254.3978, 254.3994, 254.3998, 254.4002, 254.4, 
    254.3988, 254.3986, 254.3978, 254.3976, 254.397, 254.3965, 254.3969, 
    254.3974, 254.3988, 254.4001, 254.4014, 254.4018, 254.4033, 254.402, 
    254.4041, 254.4023, 254.4055, 254.3998, 254.4023, 254.3979, 254.3984, 
    254.3992, 254.4012, 254.4001, 254.4014, 254.3986, 254.3972, 254.3968, 
    254.3961, 254.3968, 254.3968, 254.3975, 254.3972, 254.3989, 254.398, 
    254.4005, 254.4014, 254.404, 254.4055, 254.4072, 254.4079, 254.4081, 
    254.4082,
  255.5029, 255.5043, 255.5041, 255.5052, 255.5046, 255.5054, 255.5032, 
    255.5044, 255.5036, 255.503, 255.5075, 255.5053, 255.5099, 255.5085, 
    255.5121, 255.5097, 255.5126, 255.5121, 255.5138, 255.5133, 255.5155, 
    255.5141, 255.5166, 255.5152, 255.5154, 255.514, 255.5058, 255.5072, 
    255.5057, 255.5059, 255.5058, 255.5046, 255.504, 255.5028, 255.503, 
    255.5039, 255.506, 255.5053, 255.5071, 255.507, 255.509, 255.5081, 
    255.5115, 255.5106, 255.5134, 255.5126, 255.5133, 255.5131, 255.5133, 
    255.5123, 255.5127, 255.5118, 255.5083, 255.5093, 255.5063, 255.5044, 
    255.5032, 255.5024, 255.5025, 255.5027, 255.5039, 255.505, 255.5059, 
    255.5065, 255.507, 255.5087, 255.5096, 255.5117, 255.5113, 255.5119, 
    255.5126, 255.5136, 255.5134, 255.5139, 255.512, 255.5132, 255.5111, 
    255.5117, 255.5071, 255.5055, 255.5047, 255.5041, 255.5026, 255.5036, 
    255.5032, 255.5042, 255.5049, 255.5045, 255.5065, 255.5057, 255.5097, 
    255.508, 255.5125, 255.5114, 255.5128, 255.5121, 255.5132, 255.5122, 
    255.514, 255.5144, 255.5141, 255.5152, 255.5121, 255.5133, 255.5045, 
    255.5046, 255.5048, 255.5038, 255.5037, 255.5028, 255.5036, 255.504, 
    255.5049, 255.5054, 255.506, 255.5071, 255.5084, 255.5102, 255.5115, 
    255.5124, 255.5118, 255.5123, 255.5118, 255.5115, 255.5143, 255.5127, 
    255.5151, 255.5149, 255.5139, 255.515, 255.5046, 255.5043, 255.5033, 
    255.5041, 255.5027, 255.5034, 255.5039, 255.5057, 255.5061, 255.5065, 
    255.5072, 255.5082, 255.5098, 255.5113, 255.5126, 255.5125, 255.5125, 
    255.5128, 255.5121, 255.513, 255.5131, 255.5127, 255.5149, 255.5143, 
    255.5149, 255.5145, 255.5044, 255.5049, 255.5047, 255.5051, 255.5048, 
    255.5063, 255.5068, 255.509, 255.5081, 255.5096, 255.5083, 255.5085, 
    255.5096, 255.5084, 255.5112, 255.5092, 255.5128, 255.5109, 255.513, 
    255.5126, 255.5132, 255.5138, 255.5145, 255.5157, 255.5154, 255.5165, 
    255.5057, 255.5063, 255.5062, 255.5069, 255.5074, 255.5085, 255.5102, 
    255.5096, 255.5108, 255.511, 255.5092, 255.5103, 255.5067, 255.5073, 
    255.507, 255.5057, 255.5097, 255.5076, 255.5115, 255.5104, 255.5137, 
    255.512, 255.5153, 255.5166, 255.518, 255.5195, 255.5067, 255.5062, 
    255.507, 255.5081, 255.5091, 255.5104, 255.5106, 255.5108, 255.5115, 
    255.5121, 255.5109, 255.5122, 255.5074, 255.5099, 255.506, 255.5072, 
    255.508, 255.5077, 255.5095, 255.51, 255.5117, 255.5108, 255.5163, 
    255.5139, 255.5207, 255.5188, 255.5061, 255.5067, 255.5087, 255.5077, 
    255.5105, 255.5112, 255.5118, 255.5125, 255.5126, 255.513, 255.5123, 
    255.513, 255.5104, 255.5116, 255.5085, 255.5092, 255.5089, 255.5085, 
    255.5097, 255.5109, 255.511, 255.5114, 255.5124, 255.5106, 255.5166, 
    255.5128, 255.5073, 255.5084, 255.5086, 255.5082, 255.5112, 255.5101, 
    255.513, 255.5122, 255.5135, 255.5129, 255.5128, 255.5119, 255.5114, 
    255.5101, 255.509, 255.5082, 255.5084, 255.5093, 255.511, 255.5126, 
    255.5122, 255.5134, 255.5103, 255.5116, 255.5111, 255.5124, 255.5096, 
    255.5119, 255.509, 255.5092, 255.51, 255.5117, 255.5121, 255.5125, 
    255.5122, 255.511, 255.5109, 255.51, 255.5098, 255.5092, 255.5086, 
    255.5091, 255.5096, 255.511, 255.5123, 255.5138, 255.5141, 255.5157, 
    255.5144, 255.5166, 255.5146, 255.518, 255.5121, 255.5146, 255.5101, 
    255.5106, 255.5115, 255.5135, 255.5124, 255.5137, 255.5108, 255.5093, 
    255.509, 255.5083, 255.509, 255.5089, 255.5096, 255.5094, 255.5111, 
    255.5102, 255.5128, 255.5137, 255.5164, 255.5181, 255.5198, 255.5205, 
    255.5208, 255.5208,
  257.1093, 257.1106, 257.1104, 257.1115, 257.1108, 257.1115, 257.1096, 
    257.1107, 257.11, 257.1094, 257.1135, 257.1115, 257.1157, 257.1144, 
    257.1178, 257.1155, 257.1182, 257.1177, 257.1193, 257.1189, 257.1208, 
    257.1195, 257.1219, 257.1205, 257.1207, 257.1195, 257.1119, 257.1133, 
    257.1118, 257.112, 257.1119, 257.1109, 257.1103, 257.1092, 257.1094, 
    257.1102, 257.1121, 257.1115, 257.1131, 257.1131, 257.1149, 257.1141, 
    257.1172, 257.1163, 257.1189, 257.1182, 257.1188, 257.1187, 257.1188, 
    257.1179, 257.1183, 257.1175, 257.1142, 257.1152, 257.1124, 257.1107, 
    257.1096, 257.1088, 257.1089, 257.1092, 257.1102, 257.1113, 257.112, 
    257.1125, 257.1131, 257.1146, 257.1154, 257.1173, 257.117, 257.1176, 
    257.1182, 257.1191, 257.1189, 257.1194, 257.1176, 257.1187, 257.1168, 
    257.1173, 257.1131, 257.1117, 257.111, 257.1104, 257.109, 257.11, 
    257.1096, 257.1105, 257.1111, 257.1108, 257.1126, 257.1119, 257.1155, 
    257.1139, 257.1181, 257.1171, 257.1183, 257.1177, 257.1188, 257.1178, 
    257.1195, 257.1199, 257.1196, 257.1206, 257.1178, 257.1188, 257.1108, 
    257.1108, 257.1111, 257.1101, 257.11, 257.1092, 257.11, 257.1103, 
    257.1111, 257.1116, 257.1121, 257.1131, 257.1143, 257.1159, 257.1172, 
    257.118, 257.1175, 257.1179, 257.1174, 257.1172, 257.1197, 257.1183, 
    257.1205, 257.1203, 257.1194, 257.1204, 257.1109, 257.1106, 257.1097, 
    257.1104, 257.1091, 257.1098, 257.1102, 257.1119, 257.1123, 257.1126, 
    257.1133, 257.1141, 257.1156, 257.1169, 257.1182, 257.1181, 257.1181, 
    257.1184, 257.1177, 257.1185, 257.1187, 257.1183, 257.1203, 257.1198, 
    257.1203, 257.12, 257.1107, 257.1111, 257.1109, 257.1114, 257.111, 
    257.1125, 257.1129, 257.1149, 257.1141, 257.1154, 257.1142, 257.1144, 
    257.1154, 257.1143, 257.1169, 257.1151, 257.1184, 257.1166, 257.1185, 
    257.1182, 257.1187, 257.1193, 257.1199, 257.1211, 257.1208, 257.1218, 
    257.1118, 257.1124, 257.1124, 257.113, 257.1134, 257.1144, 257.116, 
    257.1154, 257.1165, 257.1168, 257.1151, 257.1161, 257.1128, 257.1133, 
    257.113, 257.1118, 257.1155, 257.1136, 257.1172, 257.1161, 257.1192, 
    257.1176, 257.1207, 257.1219, 257.1232, 257.1246, 257.1127, 257.1123, 
    257.113, 257.114, 257.115, 257.1162, 257.1163, 257.1165, 257.1172, 
    257.1177, 257.1166, 257.1178, 257.1134, 257.1157, 257.1122, 257.1132, 
    257.114, 257.1136, 257.1154, 257.1158, 257.1174, 257.1165, 257.1216, 
    257.1193, 257.1257, 257.1239, 257.1122, 257.1127, 257.1146, 257.1137, 
    257.1163, 257.1169, 257.1175, 257.1181, 257.1182, 257.1186, 257.1179, 
    257.1186, 257.1162, 257.1172, 257.1144, 257.1151, 257.1148, 257.1144, 
    257.1155, 257.1166, 257.1167, 257.117, 257.118, 257.1163, 257.1218, 
    257.1183, 257.1133, 257.1143, 257.1145, 257.1141, 257.1169, 257.1158, 
    257.1186, 257.1178, 257.119, 257.1184, 257.1183, 257.1176, 257.1171, 
    257.1159, 257.1149, 257.1142, 257.1143, 257.1152, 257.1167, 257.1182, 
    257.1179, 257.119, 257.1161, 257.1173, 257.1168, 257.118, 257.1154, 
    257.1176, 257.1148, 257.1151, 257.1158, 257.1173, 257.1177, 257.1181, 
    257.1179, 257.1168, 257.1166, 257.1158, 257.1156, 257.115, 257.1145, 
    257.115, 257.1154, 257.1168, 257.118, 257.1193, 257.1196, 257.1211, 
    257.1198, 257.1219, 257.1201, 257.1232, 257.1177, 257.1201, 257.1159, 
    257.1163, 257.1171, 257.119, 257.118, 257.1192, 257.1166, 257.1152, 
    257.1149, 257.1142, 257.1149, 257.1148, 257.1155, 257.1153, 257.1168, 
    257.116, 257.1183, 257.1192, 257.1217, 257.1232, 257.1248, 257.1255, 
    257.1257, 257.1258,
  259.2229, 259.2238, 259.2236, 259.2244, 259.224, 259.2245, 259.2231, 
    259.2238, 259.2234, 259.223, 259.2259, 259.2245, 259.2275, 259.2266, 
    259.229, 259.2274, 259.2294, 259.229, 259.2302, 259.2299, 259.2313, 
    259.2303, 259.2321, 259.2311, 259.2313, 259.2303, 259.2248, 259.2257, 
    259.2247, 259.2249, 259.2248, 259.224, 259.2236, 259.2228, 259.2229, 
    259.2235, 259.2249, 259.2245, 259.2256, 259.2256, 259.2269, 259.2263, 
    259.2286, 259.228, 259.2299, 259.2294, 259.2298, 259.2297, 259.2298, 
    259.2291, 259.2294, 259.2288, 259.2264, 259.2271, 259.2251, 259.2238, 
    259.2231, 259.2225, 259.2226, 259.2228, 259.2235, 259.2243, 259.2249, 
    259.2252, 259.2256, 259.2267, 259.2274, 259.2287, 259.2285, 259.2289, 
    259.2293, 259.23, 259.2299, 259.2302, 259.2289, 259.2298, 259.2284, 
    259.2287, 259.2256, 259.2246, 259.2241, 259.2237, 259.2227, 259.2234, 
    259.2231, 259.2238, 259.2242, 259.224, 259.2253, 259.2247, 259.2274, 
    259.2262, 259.2293, 259.2285, 259.2295, 259.229, 259.2298, 259.2291, 
    259.2303, 259.2306, 259.2304, 259.2311, 259.229, 259.2298, 259.2239, 
    259.224, 259.2242, 259.2234, 259.2234, 259.2228, 259.2234, 259.2236, 
    259.2242, 259.2245, 259.2249, 259.2256, 259.2265, 259.2277, 259.2286, 
    259.2292, 259.2288, 259.2292, 259.2288, 259.2286, 259.2305, 259.2294, 
    259.231, 259.231, 259.2302, 259.231, 259.224, 259.2238, 259.2231, 
    259.2237, 259.2227, 259.2232, 259.2235, 259.2247, 259.225, 259.2253, 
    259.2257, 259.2264, 259.2275, 259.2285, 259.2294, 259.2293, 259.2293, 
    259.2295, 259.229, 259.2296, 259.2297, 259.2294, 259.2309, 259.2305, 
    259.231, 259.2307, 259.2239, 259.2242, 259.224, 259.2244, 259.2241, 
    259.2252, 259.2255, 259.227, 259.2263, 259.2273, 259.2264, 259.2266, 
    259.2273, 259.2265, 259.2284, 259.2271, 259.2295, 259.2282, 259.2296, 
    259.2294, 259.2298, 259.2301, 259.2306, 259.2315, 259.2313, 259.2321, 
    259.2247, 259.2251, 259.2251, 259.2255, 259.2259, 259.2266, 259.2278, 
    259.2273, 259.2281, 259.2283, 259.2271, 259.2278, 259.2254, 259.2258, 
    259.2256, 259.2247, 259.2274, 259.226, 259.2286, 259.2278, 259.2301, 
    259.2289, 259.2312, 259.2321, 259.2331, 259.2341, 259.2253, 259.2251, 
    259.2256, 259.2263, 259.227, 259.2279, 259.228, 259.2281, 259.2286, 
    259.229, 259.2282, 259.2291, 259.2258, 259.2275, 259.2249, 259.2257, 
    259.2263, 259.226, 259.2273, 259.2276, 259.2288, 259.2281, 259.2319, 
    259.2302, 259.235, 259.2336, 259.225, 259.2253, 259.2267, 259.2261, 
    259.228, 259.2284, 259.2288, 259.2293, 259.2293, 259.2296, 259.2292, 
    259.2296, 259.2279, 259.2287, 259.2266, 259.2271, 259.2268, 259.2266, 
    259.2274, 259.2282, 259.2282, 259.2285, 259.2292, 259.228, 259.2321, 
    259.2295, 259.2258, 259.2265, 259.2267, 259.2263, 259.2284, 259.2276, 
    259.2296, 259.2291, 259.23, 259.2296, 259.2295, 259.2289, 259.2285, 
    259.2277, 259.227, 259.2264, 259.2265, 259.2271, 259.2283, 259.2293, 
    259.2291, 259.2299, 259.2278, 259.2287, 259.2283, 259.2292, 259.2273, 
    259.2289, 259.2269, 259.2271, 259.2276, 259.2287, 259.229, 259.2293, 
    259.2291, 259.2283, 259.2282, 259.2276, 259.2274, 259.227, 259.2267, 
    259.227, 259.2273, 259.2283, 259.2292, 259.2302, 259.2304, 259.2315, 
    259.2306, 259.2321, 259.2308, 259.2331, 259.229, 259.2308, 259.2277, 
    259.228, 259.2286, 259.23, 259.2292, 259.2301, 259.2281, 259.2271, 
    259.2269, 259.2264, 259.2269, 259.2269, 259.2274, 259.2272, 259.2283, 
    259.2277, 259.2295, 259.2301, 259.232, 259.2331, 259.2343, 259.2348, 
    259.235, 259.2351,
  261.4069, 261.4073, 261.4072, 261.4076, 261.4074, 261.4076, 261.407, 
    261.4073, 261.4071, 261.4069, 261.4083, 261.4076, 261.4091, 261.4086, 
    261.4098, 261.409, 261.41, 261.4098, 261.4104, 261.4102, 261.4109, 
    261.4105, 261.4113, 261.4108, 261.4109, 261.4104, 261.4077, 261.4082, 
    261.4077, 261.4078, 261.4077, 261.4074, 261.4072, 261.4068, 261.4069, 
    261.4072, 261.4078, 261.4076, 261.4082, 261.4081, 261.4088, 261.4085, 
    261.4096, 261.4093, 261.4102, 261.41, 261.4102, 261.4101, 261.4102, 
    261.4099, 261.41, 261.4097, 261.4085, 261.4089, 261.4079, 261.4073, 
    261.407, 261.4067, 261.4067, 261.4068, 261.4072, 261.4075, 261.4078, 
    261.408, 261.4081, 261.4087, 261.409, 261.4097, 261.4095, 261.4098, 
    261.4099, 261.4103, 261.4102, 261.4104, 261.4098, 261.4102, 261.4095, 
    261.4097, 261.4082, 261.4077, 261.4074, 261.4072, 261.4068, 261.4071, 
    261.407, 261.4073, 261.4075, 261.4074, 261.408, 261.4077, 261.409, 
    261.4084, 261.4099, 261.4096, 261.41, 261.4098, 261.4102, 261.4098, 
    261.4104, 261.4106, 261.4105, 261.4109, 261.4098, 261.4102, 261.4074, 
    261.4074, 261.4075, 261.4071, 261.4071, 261.4068, 261.4071, 261.4072, 
    261.4075, 261.4077, 261.4078, 261.4082, 261.4086, 261.4091, 261.4096, 
    261.4099, 261.4097, 261.4099, 261.4097, 261.4096, 261.4105, 261.41, 
    261.4108, 261.4107, 261.4104, 261.4108, 261.4074, 261.4073, 261.407, 
    261.4072, 261.4068, 261.407, 261.4072, 261.4077, 261.4079, 261.408, 
    261.4082, 261.4085, 261.4091, 261.4095, 261.41, 261.4099, 261.4099, 
    261.41, 261.4098, 261.4101, 261.4101, 261.41, 261.4107, 261.4105, 
    261.4107, 261.4106, 261.4073, 261.4075, 261.4074, 261.4076, 261.4074, 
    261.4079, 261.4081, 261.4088, 261.4085, 261.409, 261.4085, 261.4086, 
    261.409, 261.4086, 261.4095, 261.4088, 261.41, 261.4094, 261.4101, 
    261.41, 261.4102, 261.4103, 261.4106, 261.411, 261.4109, 261.4113, 
    261.4077, 261.4079, 261.4079, 261.4081, 261.4083, 261.4086, 261.4092, 
    261.409, 261.4094, 261.4095, 261.4088, 261.4092, 261.4081, 261.4082, 
    261.4081, 261.4077, 261.409, 261.4083, 261.4096, 261.4092, 261.4103, 
    261.4098, 261.4109, 261.4113, 261.4118, 261.4124, 261.408, 261.4079, 
    261.4081, 261.4085, 261.4088, 261.4092, 261.4093, 261.4094, 261.4096, 
    261.4098, 261.4094, 261.4098, 261.4083, 261.4091, 261.4078, 261.4082, 
    261.4084, 261.4084, 261.4089, 261.4091, 261.4097, 261.4094, 261.4112, 
    261.4104, 261.4128, 261.4121, 261.4078, 261.408, 261.4087, 261.4084, 
    261.4093, 261.4095, 261.4097, 261.4099, 261.41, 261.4101, 261.4099, 
    261.4101, 261.4092, 261.4096, 261.4086, 261.4088, 261.4088, 261.4086, 
    261.409, 261.4094, 261.4094, 261.4095, 261.4099, 261.4093, 261.4113, 
    261.41, 261.4082, 261.4086, 261.4086, 261.4085, 261.4095, 261.4091, 
    261.4101, 261.4098, 261.4103, 261.4101, 261.41, 261.4097, 261.4096, 
    261.4091, 261.4088, 261.4085, 261.4086, 261.4089, 261.4094, 261.41, 
    261.4099, 261.4102, 261.4092, 261.4096, 261.4095, 261.4099, 261.409, 
    261.4097, 261.4088, 261.4088, 261.4091, 261.4097, 261.4098, 261.4099, 
    261.4099, 261.4095, 261.4094, 261.4091, 261.409, 261.4088, 261.4087, 
    261.4088, 261.409, 261.4095, 261.4099, 261.4103, 261.4105, 261.411, 
    261.4106, 261.4113, 261.4106, 261.4118, 261.4098, 261.4106, 261.4091, 
    261.4093, 261.4096, 261.4103, 261.4099, 261.4103, 261.4094, 261.4089, 
    261.4088, 261.4085, 261.4088, 261.4088, 261.409, 261.4089, 261.4095, 
    261.4092, 261.41, 261.4103, 261.4113, 261.4118, 261.4124, 261.4127, 
    261.4128, 261.4128,
  262.7627, 262.7628, 262.7628, 262.7629, 262.7628, 262.7629, 262.7628, 
    262.7628, 262.7628, 262.7627, 262.7631, 262.7629, 262.7632, 262.7631, 
    262.7634, 262.7632, 262.7635, 262.7634, 262.7635, 262.7635, 262.7637, 
    262.7636, 262.7638, 262.7637, 262.7637, 262.7636, 262.7629, 262.763, 
    262.7629, 262.7629, 262.7629, 262.7628, 262.7628, 262.7627, 262.7627, 
    262.7628, 262.7629, 262.7629, 262.763, 262.763, 262.7632, 262.7631, 
    262.7634, 262.7633, 262.7635, 262.7635, 262.7635, 262.7635, 262.7635, 
    262.7634, 262.7635, 262.7634, 262.7631, 262.7632, 262.763, 262.7628, 
    262.7628, 262.7627, 262.7627, 262.7627, 262.7628, 262.7629, 262.7629, 
    262.763, 262.763, 262.7631, 262.7632, 262.7634, 262.7633, 262.7634, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7634, 262.7635, 262.7633, 
    262.7634, 262.763, 262.7629, 262.7628, 262.7628, 262.7627, 262.7628, 
    262.7628, 262.7628, 262.7628, 262.7628, 262.763, 262.7629, 262.7632, 
    262.7631, 262.7634, 262.7633, 262.7635, 262.7634, 262.7635, 262.7634, 
    262.7636, 262.7636, 262.7636, 262.7637, 262.7634, 262.7635, 262.7628, 
    262.7628, 262.7628, 262.7628, 262.7628, 262.7627, 262.7628, 262.7628, 
    262.7628, 262.7629, 262.7629, 262.763, 262.7631, 262.7632, 262.7634, 
    262.7634, 262.7634, 262.7634, 262.7634, 262.7634, 262.7636, 262.7635, 
    262.7637, 262.7636, 262.7635, 262.7636, 262.7628, 262.7628, 262.7628, 
    262.7628, 262.7627, 262.7628, 262.7628, 262.7629, 262.7629, 262.763, 
    262.763, 262.7631, 262.7632, 262.7633, 262.7635, 262.7634, 262.7635, 
    262.7635, 262.7634, 262.7635, 262.7635, 262.7635, 262.7636, 262.7636, 
    262.7636, 262.7636, 262.7628, 262.7628, 262.7628, 262.7629, 262.7628, 
    262.763, 262.763, 262.7632, 262.7631, 262.7632, 262.7631, 262.7631, 
    262.7632, 262.7631, 262.7633, 262.7632, 262.7635, 262.7633, 262.7635, 
    262.7635, 262.7635, 262.7635, 262.7636, 262.7637, 262.7637, 262.7638, 
    262.7629, 262.763, 262.763, 262.763, 262.763, 262.7631, 262.7632, 
    262.7632, 262.7633, 262.7633, 262.7632, 262.7633, 262.763, 262.763, 
    262.763, 262.7629, 262.7632, 262.7631, 262.7634, 262.7633, 262.7635, 
    262.7634, 262.7637, 262.7638, 262.7639, 262.7641, 262.763, 262.7629, 
    262.763, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 
    262.7634, 262.7633, 262.7634, 262.763, 262.7632, 262.7629, 262.763, 
    262.7631, 262.7631, 262.7632, 262.7632, 262.7634, 262.7633, 262.7638, 
    262.7635, 262.7642, 262.764, 262.7629, 262.763, 262.7631, 262.7631, 
    262.7633, 262.7633, 262.7634, 262.7634, 262.7635, 262.7635, 262.7634, 
    262.7635, 262.7633, 262.7634, 262.7631, 262.7632, 262.7632, 262.7631, 
    262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 262.7633, 262.7638, 
    262.7635, 262.763, 262.7631, 262.7631, 262.7631, 262.7633, 262.7632, 
    262.7635, 262.7634, 262.7635, 262.7635, 262.7635, 262.7634, 262.7634, 
    262.7632, 262.7632, 262.7631, 262.7631, 262.7632, 262.7633, 262.7635, 
    262.7634, 262.7635, 262.7633, 262.7634, 262.7633, 262.7634, 262.7632, 
    262.7634, 262.7632, 262.7632, 262.7632, 262.7634, 262.7634, 262.7634, 
    262.7634, 262.7633, 262.7633, 262.7632, 262.7632, 262.7632, 262.7631, 
    262.7632, 262.7632, 262.7633, 262.7634, 262.7635, 262.7636, 262.7637, 
    262.7636, 262.7638, 262.7636, 262.7639, 262.7634, 262.7636, 262.7632, 
    262.7633, 262.7634, 262.7635, 262.7634, 262.7635, 262.7633, 262.7632, 
    262.7632, 262.7631, 262.7632, 262.7632, 262.7632, 262.7632, 262.7633, 
    262.7632, 262.7635, 262.7635, 262.7638, 262.7639, 262.7641, 262.7642, 
    262.7642, 262.7642,
  263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1178, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 263.1177, 263.1177, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 263.1179, 
    263.1179, 263.1179,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1013, 263.1153, 263.1126, 263.1238, 263.1176, 263.1249, 263.1042, 
    263.1159, 263.1084, 263.1026, 263.1453, 263.1243, 263.167, 263.1537, 
    263.1872, 263.1649, 263.1917, 263.1866, 263.2019, 263.1975, 263.2171, 
    263.2039, 263.2272, 263.214, 263.216, 263.2035, 263.1286, 263.1426, 
    263.1277, 263.1297, 263.1288, 263.1178, 263.1121, 263.1003, 263.1024, 
    263.1111, 263.1306, 263.1241, 263.1406, 263.1403, 263.1586, 263.1504, 
    263.1812, 263.1725, 263.1977, 263.1914, 263.1974, 263.1956, 263.1974, 
    263.1881, 263.1921, 263.1839, 263.1519, 263.1613, 263.1332, 263.1161, 
    263.1047, 263.0966, 263.0977, 263.0999, 263.1112, 263.1217, 263.1297, 
    263.135, 263.1402, 263.1559, 263.1643, 263.183, 263.1796, 263.1853, 
    263.1907, 263.1998, 263.1983, 263.2024, 263.1852, 263.1966, 263.1777, 
    263.1829, 263.1415, 263.1259, 263.1191, 263.1131, 263.0986, 263.1086, 
    263.1047, 263.1141, 263.1201, 263.1171, 263.1351, 263.1281, 263.1648, 
    263.149, 263.1901, 263.1803, 263.1924, 263.1862, 263.1969, 263.1873, 
    263.2039, 263.2074, 263.205, 263.2144, 263.1868, 263.1974, 263.117, 
    263.1175, 263.1198, 263.1099, 263.1093, 263.1002, 263.1083, 263.1117, 
    263.1204, 263.1255, 263.1303, 263.1409, 263.1526, 263.1691, 263.1809, 
    263.1888, 263.184, 263.1883, 263.1835, 263.1812, 263.2061, 263.1921, 
    263.2131, 263.2119, 263.2025, 263.212, 263.1179, 263.1151, 263.1054, 
    263.113, 263.0992, 263.1069, 263.1114, 263.1283, 263.132, 263.1354, 
    263.1422, 263.1508, 263.1659, 263.179, 263.191, 263.1902, 263.1905, 
    263.1931, 263.1865, 263.1942, 263.1955, 263.1921, 263.2118, 263.2062, 
    263.2119, 263.2083, 263.116, 263.1206, 263.1181, 263.1228, 263.1195, 
    263.1342, 263.1385, 263.159, 263.1506, 263.1639, 263.1519, 263.1541, 
    263.1643, 263.1526, 263.1783, 263.1609, 263.1933, 263.1758, 263.1943, 
    263.191, 263.1965, 263.2015, 263.2077, 263.2192, 263.2166, 263.2261, 
    263.1275, 263.1335, 263.1329, 263.1392, 263.1438, 263.1537, 263.1697, 
    263.1637, 263.1747, 263.1769, 263.1602, 263.1704, 263.1374, 263.1428, 
    263.1396, 263.128, 263.165, 263.146, 263.1811, 263.1708, 263.2008, 
    263.1859, 263.2151, 263.2275, 263.2392, 263.2527, 263.1367, 263.1327, 
    263.1399, 263.1499, 263.1591, 263.1715, 263.1727, 263.175, 263.181, 
    263.186, 263.1758, 263.1873, 263.144, 263.1667, 263.1311, 263.1418, 
    263.1493, 263.146, 263.163, 263.167, 263.1832, 263.1748, 263.2244, 
    263.2025, 263.2631, 263.2462, 263.1313, 263.1367, 263.1556, 263.1466, 
    263.1723, 263.1786, 263.1837, 263.1903, 263.191, 263.1949, 263.1885, 
    263.1946, 263.1715, 263.1818, 263.1534, 263.1604, 263.1572, 263.1537, 
    263.1645, 263.1759, 263.1762, 263.1798, 263.1901, 263.1724, 263.2272, 
    263.1934, 263.1426, 263.153, 263.1546, 263.1505, 263.178, 263.168, 
    263.1948, 263.1876, 263.1994, 263.1935, 263.1926, 263.1851, 263.1804, 
    263.1685, 263.1588, 263.1511, 263.1529, 263.1613, 263.1766, 263.191, 
    263.1879, 263.1985, 263.1704, 263.1822, 263.1776, 263.1895, 263.1635, 
    263.1856, 263.1579, 263.1603, 263.1678, 263.183, 263.1864, 263.1899, 
    263.1877, 263.177, 263.1753, 263.1677, 263.1656, 263.1598, 263.155, 
    263.1593, 263.1639, 263.177, 263.1888, 263.2016, 263.2047, 263.2195, 
    263.2074, 263.2274, 263.2104, 263.2398, 263.1869, 263.2099, 263.1682, 
    263.1727, 263.1808, 263.1995, 263.1895, 263.2012, 263.1752, 263.1616, 
    263.1581, 263.1516, 263.1583, 263.1577, 263.1642, 263.1621, 263.1775, 
    263.1692, 263.1926, 263.2011, 263.2251, 263.2397, 263.2547, 263.2612, 
    263.2632, 263.2641 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9048, 253.9056, 253.9054, 253.9061, 253.9057, 253.9062, 253.9049, 
    253.9056, 253.9052, 253.9048, 253.9074, 253.9061, 253.9088, 253.908, 
    253.91, 253.9086, 253.9103, 253.91, 253.911, 253.9107, 253.9119, 
    253.9111, 253.9126, 253.9117, 253.9118, 253.9111, 253.9064, 253.9072, 
    253.9064, 253.9065, 253.9064, 253.9057, 253.9054, 253.9047, 253.9048, 
    253.9053, 253.9065, 253.9061, 253.9072, 253.9071, 253.9083, 253.9078, 
    253.9097, 253.9091, 253.9107, 253.9103, 253.9107, 253.9106, 253.9107, 
    253.9101, 253.9104, 253.9099, 253.9079, 253.9084, 253.9067, 253.9056, 
    253.905, 253.9045, 253.9045, 253.9047, 253.9053, 253.906, 253.9065, 
    253.9068, 253.9071, 253.9081, 253.9086, 253.9098, 253.9096, 253.9099, 
    253.9103, 253.9108, 253.9108, 253.911, 253.9099, 253.9106, 253.9095, 
    253.9098, 253.9072, 253.9062, 253.9058, 253.9055, 253.9046, 253.9052, 
    253.905, 253.9055, 253.9059, 253.9057, 253.9068, 253.9064, 253.9086, 
    253.9077, 253.9102, 253.9096, 253.9104, 253.91, 253.9106, 253.9101, 
    253.9111, 253.9113, 253.9112, 253.9118, 253.91, 253.9107, 253.9057, 
    253.9057, 253.9059, 253.9053, 253.9052, 253.9047, 253.9052, 253.9054, 
    253.9059, 253.9062, 253.9065, 253.9072, 253.9079, 253.9089, 253.9097, 
    253.9102, 253.9099, 253.9101, 253.9098, 253.9097, 253.9112, 253.9104, 
    253.9117, 253.9116, 253.911, 253.9116, 253.9058, 253.9056, 253.905, 
    253.9055, 253.9046, 253.9051, 253.9053, 253.9064, 253.9066, 253.9068, 
    253.9073, 253.9078, 253.9087, 253.9095, 253.9103, 253.9102, 253.9103, 
    253.9104, 253.91, 253.9105, 253.9106, 253.9104, 253.9116, 253.9112, 
    253.9116, 253.9114, 253.9056, 253.9059, 253.9058, 253.9061, 253.9059, 
    253.9067, 253.907, 253.9083, 253.9078, 253.9086, 253.9079, 253.908, 
    253.9086, 253.9079, 253.9095, 253.9084, 253.9104, 253.9093, 253.9105, 
    253.9103, 253.9106, 253.9109, 253.9113, 253.912, 253.9119, 253.9125, 
    253.9063, 253.9067, 253.9067, 253.9071, 253.9073, 253.908, 253.909, 
    253.9086, 253.9093, 253.9094, 253.9084, 253.909, 253.907, 253.9073, 
    253.9071, 253.9064, 253.9087, 253.9075, 253.9097, 253.909, 253.9109, 
    253.91, 253.9118, 253.9126, 253.9133, 253.9142, 253.9069, 253.9067, 
    253.9071, 253.9077, 253.9083, 253.9091, 253.9091, 253.9093, 253.9097, 
    253.91, 253.9093, 253.9101, 253.9073, 253.9088, 253.9066, 253.9072, 
    253.9077, 253.9075, 253.9085, 253.9088, 253.9098, 253.9093, 253.9124, 
    253.911, 253.9148, 253.9138, 253.9066, 253.9069, 253.9081, 253.9075, 
    253.9091, 253.9095, 253.9098, 253.9102, 253.9103, 253.9105, 253.9101, 
    253.9105, 253.9091, 253.9097, 253.908, 253.9084, 253.9082, 253.908, 
    253.9086, 253.9093, 253.9094, 253.9096, 253.9102, 253.9091, 253.9125, 
    253.9104, 253.9073, 253.9079, 253.908, 253.9078, 253.9095, 253.9089, 
    253.9105, 253.9101, 253.9108, 253.9104, 253.9104, 253.9099, 253.9096, 
    253.9089, 253.9083, 253.9078, 253.9079, 253.9084, 253.9094, 253.9103, 
    253.9101, 253.9108, 253.909, 253.9097, 253.9094, 253.9102, 253.9086, 
    253.9099, 253.9082, 253.9084, 253.9088, 253.9098, 253.91, 253.9102, 
    253.9101, 253.9094, 253.9093, 253.9088, 253.9087, 253.9083, 253.9081, 
    253.9083, 253.9086, 253.9094, 253.9101, 253.9109, 253.9111, 253.912, 
    253.9113, 253.9125, 253.9114, 253.9133, 253.91, 253.9114, 253.9089, 
    253.9091, 253.9096, 253.9108, 253.9102, 253.9109, 253.9093, 253.9084, 
    253.9082, 253.9078, 253.9082, 253.9082, 253.9086, 253.9085, 253.9094, 
    253.9089, 253.9104, 253.9109, 253.9124, 253.9133, 253.9143, 253.9147, 
    253.9149, 253.9149 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1399992, 0.1400071, 0.1400056, 0.1400118, 0.1400084, 0.1400125, 
    0.1400009, 0.1400073, 0.1400033, 0.14, 0.1400238, 0.1400121, 0.1400367, 
    0.1400291, 0.1400484, 0.1400354, 0.1400511, 0.1400482, 0.1400573, 
    0.1400547, 0.140066, 0.1400585, 0.1400721, 0.1400643, 0.1400655, 
    0.1400582, 0.1400146, 0.1400223, 0.1400142, 0.1400153, 0.1400148, 
    0.1400084, 0.1400052, 0.1399987, 0.1399999, 0.1400047, 0.1400158, 
    0.1400121, 0.1400216, 0.1400214, 0.140032, 0.1400272, 0.1400451, 0.14004, 
    0.1400548, 0.1400511, 0.1400546, 0.1400536, 0.1400546, 0.1400491, 
    0.1400515, 0.1400467, 0.1400281, 0.1400335, 0.1400173, 0.1400073, 
    0.1400011, 0.1399966, 0.1399973, 0.1399985, 0.1400047, 0.1400108, 
    0.1400153, 0.1400184, 0.1400214, 0.1400301, 0.1400351, 0.140046, 
    0.1400442, 0.1400474, 0.1400507, 0.140056, 0.1400552, 0.1400575, 
    0.1400474, 0.1400541, 0.1400431, 0.1400461, 0.1400217, 0.1400131, 
    0.140009, 0.1400059, 0.1399978, 0.1400033, 0.1400011, 0.1400065, 
    0.1400098, 0.1400082, 0.1400185, 0.1400144, 0.1400354, 0.1400264, 
    0.1400503, 0.1400446, 0.1400517, 0.1400481, 0.1400543, 0.1400487, 
    0.1400584, 0.1400605, 0.140059, 0.1400647, 0.1400484, 0.1400546, 
    0.1400081, 0.1400084, 0.1400097, 0.140004, 0.1400037, 0.1399987, 
    0.1400032, 0.1400051, 0.1400101, 0.1400129, 0.1400157, 0.1400217, 
    0.1400284, 0.140038, 0.140045, 0.1400496, 0.1400468, 0.1400493, 
    0.1400465, 0.1400452, 0.1400596, 0.1400515, 0.1400639, 0.1400632, 
    0.1400575, 0.1400633, 0.1400086, 0.140007, 0.1400016, 0.1400059, 
    0.1399981, 0.1400024, 0.1400048, 0.1400144, 0.1400167, 0.1400186, 
    0.1400225, 0.1400274, 0.1400361, 0.1400438, 0.1400509, 0.1400504, 
    0.1400506, 0.1400521, 0.1400483, 0.1400528, 0.1400535, 0.1400515, 
    0.1400631, 0.1400598, 0.1400632, 0.140061, 0.1400076, 0.1400101, 
    0.1400087, 0.1400114, 0.1400095, 0.1400177, 0.1400202, 0.140032, 
    0.1400273, 0.140035, 0.1400281, 0.1400293, 0.140035, 0.1400286, 
    0.1400433, 0.1400331, 0.1400522, 0.1400417, 0.1400528, 0.1400509, 
    0.1400542, 0.140057, 0.1400607, 0.1400674, 0.1400659, 0.1400716, 
    0.1400141, 0.1400174, 0.1400172, 0.1400208, 0.1400234, 0.1400292, 
    0.1400384, 0.1400349, 0.1400414, 0.1400426, 0.1400329, 0.1400388, 
    0.1400197, 0.1400227, 0.140021, 0.1400143, 0.1400356, 0.1400246, 
    0.1400451, 0.1400391, 0.1400566, 0.1400478, 0.140065, 0.1400721, 
    0.1400794, 0.1400873, 0.1400193, 0.1400171, 0.1400212, 0.1400268, 
    0.1400323, 0.1400394, 0.1400402, 0.1400415, 0.140045, 0.140048, 
    0.1400418, 0.1400487, 0.1400232, 0.1400366, 0.1400161, 0.1400221, 
    0.1400265, 0.1400247, 0.1400346, 0.1400369, 0.1400462, 0.1400414, 
    0.1400703, 0.1400575, 0.1400936, 0.1400834, 0.1400162, 0.1400194, 
    0.1400301, 0.140025, 0.14004, 0.1400436, 0.1400467, 0.1400504, 0.1400509, 
    0.1400531, 0.1400494, 0.140053, 0.1400394, 0.1400455, 0.140029, 0.140033, 
    0.1400312, 0.1400292, 0.1400354, 0.1400419, 0.1400422, 0.1400443, 
    0.1400498, 0.14004, 0.1400716, 0.1400518, 0.1400228, 0.1400286, 
    0.1400296, 0.1400273, 0.1400432, 0.1400374, 0.1400531, 0.1400489, 
    0.1400558, 0.1400523, 0.1400518, 0.1400474, 0.1400446, 0.1400377, 
    0.1400321, 0.1400277, 0.1400287, 0.1400335, 0.1400423, 0.1400508, 
    0.140049, 0.1400553, 0.1400389, 0.1400456, 0.140043, 0.14005, 0.1400348, 
    0.1400472, 0.1400316, 0.140033, 0.1400373, 0.140046, 0.1400482, 
    0.1400502, 0.140049, 0.1400426, 0.1400416, 0.1400373, 0.140036, 
    0.1400327, 0.1400299, 0.1400324, 0.140035, 0.1400427, 0.1400495, 
    0.140057, 0.1400589, 0.1400673, 0.1400603, 0.1400717, 0.1400616, 
    0.1400793, 0.1400482, 0.1400617, 0.1400376, 0.1400402, 0.1400448, 
    0.1400557, 0.14005, 0.1400567, 0.1400416, 0.1400336, 0.1400317, 
    0.1400279, 0.1400318, 0.1400315, 0.1400352, 0.140034, 0.1400429, 
    0.1400382, 0.1400518, 0.1400567, 0.1400709, 0.1400795, 0.1400886, 
    0.1400926, 0.1400938, 0.1400943,
  0.1463938, 0.1464025, 0.1464009, 0.1464078, 0.146404, 0.1464086, 0.1463957, 
    0.1464028, 0.1463983, 0.1463947, 0.1464212, 0.1464082, 0.1464355, 
    0.146427, 0.1464486, 0.1464341, 0.1464516, 0.1464484, 0.1464585, 
    0.1464556, 0.1464682, 0.1464598, 0.1464751, 0.1464663, 0.1464676, 
    0.1464595, 0.1464109, 0.1464195, 0.1464104, 0.1464116, 0.1464111, 
    0.1464041, 0.1464004, 0.1463933, 0.1463946, 0.1463999, 0.1464122, 
    0.1464081, 0.1464187, 0.1464185, 0.1464302, 0.1464249, 0.1464449, 
    0.1464392, 0.1464557, 0.1464515, 0.1464555, 0.1464543, 0.1464555, 
    0.1464494, 0.146452, 0.1464466, 0.1464259, 0.1464319, 0.1464139, 
    0.1464028, 0.146396, 0.1463909, 0.1463916, 0.146393, 0.1463999, 
    0.1464066, 0.1464117, 0.1464151, 0.1464184, 0.1464282, 0.1464337, 
    0.1464459, 0.1464439, 0.1464474, 0.1464511, 0.1464571, 0.1464561, 
    0.1464587, 0.1464475, 0.1464549, 0.1464427, 0.146446, 0.1464188, 
    0.1464092, 0.1464047, 0.1464012, 0.1463922, 0.1463984, 0.1463959, 
    0.1464019, 0.1464056, 0.1464038, 0.1464152, 0.1464107, 0.1464341, 
    0.146424, 0.1464507, 0.1464443, 0.1464522, 0.1464482, 0.1464551, 
    0.1464489, 0.1464597, 0.146462, 0.1464604, 0.1464667, 0.1464485, 
    0.1464554, 0.1464037, 0.146404, 0.1464054, 0.1463991, 0.1463988, 
    0.1463932, 0.1463982, 0.1464003, 0.1464058, 0.146409, 0.1464121, 
    0.1464188, 0.1464263, 0.1464369, 0.1464447, 0.1464499, 0.1464467, 
    0.1464495, 0.1464464, 0.1464449, 0.1464611, 0.146452, 0.1464658, 
    0.146465, 0.1464587, 0.1464651, 0.1464042, 0.1464025, 0.1463964, 
    0.1464012, 0.1463926, 0.1463973, 0.1464, 0.1464107, 0.1464132, 0.1464153, 
    0.1464197, 0.1464252, 0.1464349, 0.1464434, 0.1464513, 0.1464508, 
    0.146451, 0.1464527, 0.1464484, 0.1464534, 0.1464542, 0.146452, 
    0.1464649, 0.1464612, 0.146465, 0.1464626, 0.1464031, 0.146406, 
    0.1464044, 0.1464073, 0.1464052, 0.1464144, 0.1464172, 0.1464303, 
    0.146425, 0.1464336, 0.1464259, 0.1464273, 0.1464336, 0.1464264, 
    0.1464428, 0.1464315, 0.1464528, 0.1464411, 0.1464535, 0.1464513, 
    0.1464549, 0.1464581, 0.1464623, 0.1464698, 0.1464681, 0.1464744, 
    0.1464103, 0.146414, 0.1464138, 0.1464178, 0.1464207, 0.1464271, 
    0.1464373, 0.1464335, 0.1464407, 0.1464421, 0.1464313, 0.1464378, 
    0.1464166, 0.1464199, 0.146418, 0.1464105, 0.1464343, 0.146422, 
    0.1464448, 0.1464381, 0.1464577, 0.1464478, 0.1464671, 0.1464751, 
    0.1464832, 0.146492, 0.1464161, 0.1464136, 0.1464182, 0.1464245, 
    0.1464306, 0.1464385, 0.1464394, 0.1464409, 0.1464448, 0.146448, 
    0.1464412, 0.1464489, 0.1464204, 0.1464354, 0.1464126, 0.1464193, 
    0.1464242, 0.1464221, 0.1464331, 0.1464357, 0.1464461, 0.1464408, 
    0.146473, 0.1464587, 0.1464992, 0.1464877, 0.1464127, 0.1464162, 
    0.1464282, 0.1464225, 0.1464391, 0.1464432, 0.1464466, 0.1464508, 
    0.1464513, 0.1464538, 0.1464497, 0.1464537, 0.1464385, 0.1464453, 
    0.1464269, 0.1464313, 0.1464294, 0.1464271, 0.1464341, 0.1464413, 
    0.1464416, 0.1464439, 0.1464501, 0.1464392, 0.1464746, 0.1464524, 
    0.14642, 0.1464265, 0.1464276, 0.1464251, 0.1464428, 0.1464363, 
    0.1464538, 0.1464491, 0.1464568, 0.1464529, 0.1464524, 0.1464474, 
    0.1464444, 0.1464366, 0.1464303, 0.1464255, 0.1464266, 0.146432, 
    0.1464418, 0.1464513, 0.1464492, 0.1464562, 0.1464379, 0.1464455, 
    0.1464425, 0.1464503, 0.1464334, 0.1464473, 0.1464298, 0.1464314, 
    0.1464362, 0.1464459, 0.1464483, 0.1464505, 0.1464492, 0.1464421, 
    0.146441, 0.1464361, 0.1464347, 0.146431, 0.1464279, 0.1464307, 
    0.1464336, 0.1464421, 0.1464498, 0.1464582, 0.1464603, 0.1464697, 
    0.1464618, 0.1464747, 0.1464634, 0.1464831, 0.1464483, 0.1464634, 
    0.1464365, 0.1464394, 0.1464445, 0.1464567, 0.1464503, 0.1464578, 
    0.146441, 0.146432, 0.14643, 0.1464257, 0.1464301, 0.1464297, 0.1464339, 
    0.1464325, 0.1464424, 0.1464371, 0.1464523, 0.1464578, 0.1464737, 
    0.1464834, 0.1464936, 0.146498, 0.1464993, 0.1464999,
  0.1561807, 0.1561891, 0.1561875, 0.1561942, 0.1561905, 0.1561949, 
    0.1561824, 0.1561894, 0.156185, 0.1561815, 0.1562072, 0.1561945, 
    0.1562211, 0.1562128, 0.1562339, 0.1562197, 0.1562368, 0.1562337, 
    0.1562436, 0.1562407, 0.1562532, 0.1562449, 0.1562599, 0.1562513, 
    0.1562526, 0.1562446, 0.1561972, 0.1562056, 0.1561967, 0.1561979, 
    0.1561974, 0.1561906, 0.156187, 0.1561801, 0.1561814, 0.1561865, 
    0.1561984, 0.1561945, 0.1562048, 0.1562045, 0.156216, 0.1562108, 
    0.1562302, 0.1562247, 0.1562409, 0.1562368, 0.1562406, 0.1562395, 
    0.1562407, 0.1562347, 0.1562372, 0.156232, 0.1562117, 0.1562176, 
    0.1562001, 0.1561894, 0.1561827, 0.1561779, 0.1561786, 0.1561798, 
    0.1561866, 0.156193, 0.156198, 0.1562012, 0.1562045, 0.156214, 0.1562194, 
    0.1562313, 0.1562293, 0.1562328, 0.1562364, 0.1562422, 0.1562413, 
    0.1562438, 0.1562328, 0.15624, 0.1562281, 0.1562313, 0.1562049, 
    0.1561956, 0.1561912, 0.1561878, 0.1561791, 0.156185, 0.1561827, 
    0.1561884, 0.156192, 0.1561903, 0.1562013, 0.156197, 0.1562197, 
    0.1562099, 0.1562359, 0.1562297, 0.1562375, 0.1562335, 0.1562403, 
    0.1562342, 0.1562448, 0.156247, 0.1562455, 0.1562517, 0.1562338, 
    0.1562406, 0.1561902, 0.1561905, 0.1561918, 0.1561858, 0.1561854, 
    0.1561801, 0.1561849, 0.1561869, 0.1561923, 0.1561953, 0.1561983, 
    0.1562049, 0.1562121, 0.1562225, 0.1562301, 0.1562352, 0.1562321, 
    0.1562348, 0.1562317, 0.1562303, 0.1562462, 0.1562372, 0.1562508, 
    0.15625, 0.1562438, 0.1562501, 0.1561907, 0.156189, 0.1561832, 0.1561878, 
    0.1561795, 0.156184, 0.1561866, 0.156197, 0.1561994, 0.1562015, 
    0.1562057, 0.156211, 0.1562205, 0.1562288, 0.1562366, 0.156236, 
    0.1562362, 0.1562379, 0.1562337, 0.1562386, 0.1562394, 0.1562373, 
    0.1562499, 0.1562463, 0.15625, 0.1562477, 0.1561896, 0.1561924, 
    0.1561909, 0.1561937, 0.1561916, 0.1562006, 0.1562033, 0.156216, 
    0.1562109, 0.1562192, 0.1562118, 0.1562131, 0.1562193, 0.1562122, 
    0.1562283, 0.1562172, 0.156238, 0.1562266, 0.1562387, 0.1562366, 
    0.1562401, 0.1562433, 0.1562473, 0.1562547, 0.156253, 0.1562593, 
    0.1561966, 0.1562002, 0.1562, 0.1562038, 0.1562066, 0.1562129, 0.1562229, 
    0.1562192, 0.1562261, 0.1562275, 0.156217, 0.1562233, 0.1562027, 
    0.1562059, 0.1562041, 0.1561968, 0.1562199, 0.1562079, 0.1562302, 
    0.1562237, 0.1562428, 0.1562332, 0.1562521, 0.15626, 0.1562679, 
    0.1562767, 0.1562023, 0.1561998, 0.1562043, 0.1562104, 0.1562163, 
    0.1562241, 0.1562249, 0.1562263, 0.1562302, 0.1562334, 0.1562267, 
    0.1562342, 0.1562065, 0.156221, 0.1561988, 0.1562053, 0.15621, 0.1562081, 
    0.1562188, 0.1562213, 0.1562314, 0.1562262, 0.1562579, 0.1562438, 
    0.1562838, 0.1562724, 0.1561989, 0.1562023, 0.156214, 0.1562084, 
    0.1562246, 0.1562286, 0.1562319, 0.156236, 0.1562365, 0.156239, 0.156235, 
    0.1562389, 0.1562241, 0.1562307, 0.1562128, 0.156217, 0.1562151, 
    0.1562129, 0.1562197, 0.1562268, 0.1562271, 0.1562293, 0.1562354, 
    0.1562247, 0.1562594, 0.1562376, 0.156206, 0.1562123, 0.1562134, 
    0.1562109, 0.1562282, 0.1562219, 0.1562389, 0.1562344, 0.1562419, 
    0.1562381, 0.1562376, 0.1562328, 0.1562297, 0.1562221, 0.156216, 
    0.1562113, 0.1562124, 0.1562176, 0.1562272, 0.1562365, 0.1562345, 
    0.1562414, 0.1562234, 0.1562308, 0.1562279, 0.1562356, 0.156219, 
    0.1562326, 0.1562155, 0.1562171, 0.1562218, 0.1562312, 0.1562336, 
    0.1562358, 0.1562345, 0.1562275, 0.1562265, 0.1562217, 0.1562203, 
    0.1562167, 0.1562137, 0.1562164, 0.1562193, 0.1562276, 0.1562351, 
    0.1562433, 0.1562454, 0.1562547, 0.1562469, 0.1562596, 0.1562485, 
    0.1562679, 0.1562337, 0.1562484, 0.156222, 0.1562249, 0.1562299, 
    0.1562418, 0.1562355, 0.156243, 0.1562264, 0.1562177, 0.1562157, 
    0.1562116, 0.1562158, 0.1562155, 0.1562195, 0.1562182, 0.1562279, 
    0.1562227, 0.1562375, 0.1562429, 0.1562586, 0.1562681, 0.1562782, 
    0.1562825, 0.1562839, 0.1562845,
  0.169923, 0.1699295, 0.1699283, 0.1699335, 0.1699306, 0.169934, 0.1699243, 
    0.1699297, 0.1699263, 0.1699236, 0.1699436, 0.1699337, 0.1699545, 
    0.169948, 0.1699646, 0.1699534, 0.1699669, 0.1699644, 0.1699723, 0.16997, 
    0.1699799, 0.1699733, 0.1699853, 0.1699784, 0.1699794, 0.1699731, 
    0.1699358, 0.1699423, 0.1699354, 0.1699363, 0.1699359, 0.1699306, 
    0.1699279, 0.1699226, 0.1699236, 0.1699275, 0.1699367, 0.1699337, 
    0.1699417, 0.1699415, 0.1699504, 0.1699464, 0.1699617, 0.1699573, 
    0.1699701, 0.1699668, 0.1699699, 0.169969, 0.1699699, 0.1699652, 
    0.1699672, 0.1699631, 0.1699471, 0.1699517, 0.169938, 0.1699297, 
    0.1699246, 0.1699208, 0.1699214, 0.1699223, 0.1699275, 0.1699325, 
    0.1699364, 0.1699389, 0.1699415, 0.1699489, 0.1699531, 0.1699625, 
    0.1699609, 0.1699637, 0.1699665, 0.1699712, 0.1699704, 0.1699724, 
    0.1699637, 0.1699695, 0.16996, 0.1699625, 0.1699418, 0.1699345, 
    0.1699311, 0.1699285, 0.1699218, 0.1699264, 0.1699245, 0.169929, 
    0.1699318, 0.1699304, 0.169939, 0.1699356, 0.1699534, 0.1699457, 
    0.1699662, 0.1699612, 0.1699674, 0.1699643, 0.1699696, 0.1699648, 
    0.1699732, 0.169975, 0.1699738, 0.1699787, 0.1699645, 0.1699699, 
    0.1699303, 0.1699306, 0.1699316, 0.1699269, 0.1699267, 0.1699225, 
    0.1699262, 0.1699278, 0.1699319, 0.1699343, 0.1699366, 0.1699417, 
    0.1699474, 0.1699556, 0.1699616, 0.1699656, 0.1699631, 0.1699653, 
    0.1699629, 0.1699618, 0.1699743, 0.1699672, 0.169978, 0.1699774, 
    0.1699725, 0.1699775, 0.1699307, 0.1699294, 0.1699249, 0.1699285, 
    0.1699221, 0.1699256, 0.1699276, 0.1699356, 0.1699375, 0.1699391, 
    0.1699424, 0.1699466, 0.169954, 0.1699606, 0.1699667, 0.1699663, 
    0.1699664, 0.1699677, 0.1699644, 0.1699683, 0.1699689, 0.1699672, 
    0.1699773, 0.1699744, 0.1699774, 0.1699755, 0.1699299, 0.169932, 
    0.1699309, 0.1699331, 0.1699315, 0.1699384, 0.1699405, 0.1699505, 
    0.1699465, 0.169953, 0.1699472, 0.1699482, 0.169953, 0.1699475, 
    0.1699601, 0.1699514, 0.1699678, 0.1699588, 0.1699684, 0.1699667, 
    0.1699695, 0.169972, 0.1699752, 0.1699811, 0.1699798, 0.1699848, 
    0.1699353, 0.1699381, 0.1699379, 0.1699409, 0.1699431, 0.169948, 
    0.1699559, 0.169953, 0.1699584, 0.1699595, 0.1699512, 0.1699562, 
    0.1699401, 0.1699426, 0.1699411, 0.1699355, 0.1699535, 0.1699442, 
    0.1699616, 0.1699565, 0.1699716, 0.169964, 0.169979, 0.1699853, 
    0.1699917, 0.1699988, 0.1699397, 0.1699378, 0.1699413, 0.169946, 
    0.1699507, 0.1699568, 0.1699575, 0.1699586, 0.1699616, 0.1699641, 
    0.1699589, 0.1699648, 0.169943, 0.1699544, 0.169937, 0.1699421, 
    0.1699458, 0.1699442, 0.1699526, 0.1699546, 0.1699626, 0.1699585, 
    0.1699837, 0.1699724, 0.1700045, 0.1699954, 0.1699371, 0.1699398, 
    0.1699489, 0.1699445, 0.1699573, 0.1699604, 0.169963, 0.1699663, 
    0.1699667, 0.1699686, 0.1699654, 0.1699685, 0.1699568, 0.169962, 
    0.1699479, 0.1699513, 0.1699498, 0.169948, 0.1699534, 0.1699589, 
    0.1699592, 0.169961, 0.1699658, 0.1699573, 0.169985, 0.1699675, 
    0.1699426, 0.1699476, 0.1699484, 0.1699465, 0.1699601, 0.1699551, 
    0.1699686, 0.1699649, 0.1699709, 0.1699679, 0.1699675, 0.1699637, 
    0.1699613, 0.1699553, 0.1699505, 0.1699468, 0.1699477, 0.1699518, 
    0.1699593, 0.1699666, 0.169965, 0.1699705, 0.1699563, 0.1699622, 
    0.1699599, 0.1699659, 0.1699529, 0.1699636, 0.1699501, 0.1699513, 
    0.169955, 0.1699625, 0.1699643, 0.1699661, 0.169965, 0.1699595, 
    0.1699587, 0.1699549, 0.1699538, 0.169951, 0.1699487, 0.1699508, 
    0.169953, 0.1699596, 0.1699655, 0.169972, 0.1699737, 0.1699811, 
    0.1699749, 0.169985, 0.1699762, 0.1699917, 0.1699644, 0.1699761, 
    0.1699552, 0.1699575, 0.1699614, 0.1699709, 0.1699659, 0.1699718, 
    0.1699587, 0.1699518, 0.1699502, 0.169947, 0.1699503, 0.16995, 0.1699532, 
    0.1699522, 0.1699598, 0.1699557, 0.1699674, 0.1699717, 0.1699842, 
    0.1699919, 0.17, 0.1700035, 0.1700046, 0.1700051,
  0.1852191, 0.1852224, 0.1852218, 0.1852244, 0.185223, 0.1852247, 0.1852198, 
    0.1852225, 0.1852208, 0.1852195, 0.1852296, 0.1852246, 0.1852353, 
    0.1852319, 0.1852407, 0.1852348, 0.1852419, 0.1852406, 0.1852448, 
    0.1852436, 0.1852489, 0.1852453, 0.1852518, 0.1852481, 0.1852486, 
    0.1852452, 0.1852256, 0.185229, 0.1852254, 0.1852259, 0.1852257, 
    0.185223, 0.1852216, 0.1852189, 0.1852194, 0.1852214, 0.1852261, 
    0.1852245, 0.1852286, 0.1852286, 0.1852332, 0.1852311, 0.1852391, 
    0.1852368, 0.1852436, 0.1852419, 0.1852435, 0.185243, 0.1852435, 
    0.185241, 0.1852421, 0.1852399, 0.1852315, 0.1852339, 0.1852268, 
    0.1852225, 0.1852199, 0.1852181, 0.1852183, 0.1852188, 0.1852214, 
    0.185224, 0.1852259, 0.1852272, 0.1852285, 0.1852324, 0.1852346, 
    0.1852396, 0.1852387, 0.1852402, 0.1852417, 0.1852442, 0.1852438, 
    0.1852449, 0.1852402, 0.1852433, 0.1852382, 0.1852396, 0.1852287, 
    0.185225, 0.1852232, 0.1852219, 0.1852185, 0.1852208, 0.1852199, 
    0.1852221, 0.1852236, 0.1852229, 0.1852273, 0.1852255, 0.1852347, 
    0.1852307, 0.1852415, 0.1852389, 0.1852422, 0.1852405, 0.1852434, 
    0.1852408, 0.1852453, 0.1852463, 0.1852456, 0.1852482, 0.1852406, 
    0.1852435, 0.1852228, 0.185223, 0.1852235, 0.1852211, 0.185221, 
    0.1852189, 0.1852208, 0.1852216, 0.1852237, 0.1852249, 0.1852261, 
    0.1852287, 0.1852316, 0.1852359, 0.1852391, 0.1852412, 0.1852399, 
    0.185241, 0.1852397, 0.1852392, 0.1852459, 0.1852421, 0.1852479, 
    0.1852475, 0.1852449, 0.1852476, 0.185223, 0.1852224, 0.1852201, 
    0.1852219, 0.1852187, 0.1852204, 0.1852214, 0.1852255, 0.1852265, 
    0.1852273, 0.185229, 0.1852312, 0.1852351, 0.1852385, 0.1852418, 
    0.1852416, 0.1852416, 0.1852424, 0.1852406, 0.1852427, 0.185243, 
    0.1852421, 0.1852475, 0.1852459, 0.1852475, 0.1852465, 0.1852226, 
    0.1852237, 0.1852231, 0.1852242, 0.1852234, 0.185227, 0.185228, 
    0.1852332, 0.1852311, 0.1852345, 0.1852315, 0.185232, 0.1852346, 
    0.1852317, 0.1852383, 0.1852337, 0.1852424, 0.1852376, 0.1852427, 
    0.1852418, 0.1852433, 0.1852446, 0.1852464, 0.1852496, 0.1852488, 
    0.1852515, 0.1852254, 0.1852268, 0.1852267, 0.1852283, 0.1852294, 
    0.185232, 0.1852361, 0.1852345, 0.1852374, 0.185238, 0.1852336, 
    0.1852362, 0.1852278, 0.1852291, 0.1852284, 0.1852255, 0.1852348, 
    0.1852299, 0.1852391, 0.1852364, 0.1852444, 0.1852404, 0.1852484, 
    0.1852518, 0.1852553, 0.1852592, 0.1852276, 0.1852267, 0.1852285, 
    0.1852309, 0.1852333, 0.1852365, 0.1852369, 0.1852375, 0.1852391, 
    0.1852404, 0.1852376, 0.1852408, 0.1852293, 0.1852353, 0.1852263, 
    0.1852289, 0.1852308, 0.18523, 0.1852344, 0.1852354, 0.1852396, 
    0.1852375, 0.185251, 0.1852449, 0.1852624, 0.1852573, 0.1852263, 
    0.1852277, 0.1852324, 0.1852301, 0.1852368, 0.1852384, 0.1852398, 
    0.1852416, 0.1852418, 0.1852428, 0.1852411, 0.1852428, 0.1852366, 
    0.1852393, 0.1852319, 0.1852337, 0.1852328, 0.185232, 0.1852347, 
    0.1852377, 0.1852378, 0.1852387, 0.1852413, 0.1852368, 0.1852516, 
    0.1852422, 0.1852292, 0.1852317, 0.1852322, 0.1852311, 0.1852383, 
    0.1852356, 0.1852428, 0.1852408, 0.1852441, 0.1852425, 0.1852422, 
    0.1852402, 0.1852389, 0.1852358, 0.1852332, 0.1852313, 0.1852318, 
    0.1852339, 0.1852379, 0.1852418, 0.1852409, 0.1852438, 0.1852363, 
    0.1852394, 0.1852382, 0.1852414, 0.1852345, 0.1852401, 0.185233, 
    0.1852337, 0.1852356, 0.1852395, 0.1852405, 0.1852415, 0.1852409, 
    0.185238, 0.1852375, 0.1852356, 0.185235, 0.1852335, 0.1852323, 
    0.1852334, 0.1852346, 0.185238, 0.1852411, 0.1852446, 0.1852455, 
    0.1852495, 0.1852462, 0.1852517, 0.1852469, 0.1852553, 0.1852406, 
    0.1852468, 0.1852357, 0.1852369, 0.185239, 0.185244, 0.1852414, 
    0.1852445, 0.1852375, 0.1852339, 0.1852331, 0.1852314, 0.1852331, 
    0.185233, 0.1852347, 0.1852341, 0.1852381, 0.185236, 0.1852422, 
    0.1852445, 0.1852512, 0.1852554, 0.1852599, 0.1852619, 0.1852625, 
    0.1852627,
  0.195451, 0.1954518, 0.1954516, 0.1954522, 0.1954519, 0.1954523, 0.1954511, 
    0.1954518, 0.1954514, 0.195451, 0.1954535, 0.1954523, 0.195455, 
    0.1954541, 0.1954564, 0.1954548, 0.1954567, 0.1954563, 0.1954575, 
    0.1954571, 0.1954586, 0.1954576, 0.1954594, 0.1954584, 0.1954585, 
    0.1954576, 0.1954525, 0.1954534, 0.1954525, 0.1954526, 0.1954525, 
    0.1954519, 0.1954516, 0.1954509, 0.195451, 0.1954515, 0.1954526, 
    0.1954523, 0.1954533, 0.1954533, 0.1954544, 0.1954539, 0.195456, 
    0.1954554, 0.1954571, 0.1954567, 0.1954571, 0.195457, 0.1954571, 
    0.1954564, 0.1954567, 0.1954562, 0.195454, 0.1954546, 0.1954528, 
    0.1954518, 0.1954512, 0.1954507, 0.1954508, 0.1954509, 0.1954515, 
    0.1954521, 0.1954526, 0.1954529, 0.1954533, 0.1954542, 0.1954548, 
    0.1954561, 0.1954558, 0.1954562, 0.1954566, 0.1954573, 0.1954572, 
    0.1954575, 0.1954563, 0.1954571, 0.1954557, 0.1954561, 0.1954533, 
    0.1954524, 0.1954519, 0.1954516, 0.1954508, 0.1954514, 0.1954512, 
    0.1954517, 0.195452, 0.1954519, 0.1954529, 0.1954525, 0.1954548, 
    0.1954538, 0.1954566, 0.1954559, 0.1954568, 0.1954563, 0.1954571, 
    0.1954564, 0.1954576, 0.1954579, 0.1954577, 0.1954584, 0.1954564, 
    0.1954571, 0.1954519, 0.1954519, 0.195452, 0.1954514, 0.1954514, 
    0.1954509, 0.1954513, 0.1954515, 0.195452, 0.1954523, 0.1954526, 
    0.1954533, 0.195454, 0.1954551, 0.1954559, 0.1954565, 0.1954562, 
    0.1954565, 0.1954561, 0.195456, 0.1954578, 0.1954567, 0.1954583, 
    0.1954582, 0.1954575, 0.1954582, 0.1954519, 0.1954518, 0.1954512, 
    0.1954516, 0.1954509, 0.1954513, 0.1954515, 0.1954525, 0.1954527, 
    0.1954529, 0.1954534, 0.1954539, 0.1954549, 0.1954558, 0.1954567, 
    0.1954566, 0.1954566, 0.1954568, 0.1954563, 0.1954569, 0.195457, 
    0.1954567, 0.1954582, 0.1954578, 0.1954582, 0.1954579, 0.1954518, 
    0.1954521, 0.1954519, 0.1954522, 0.195452, 0.1954529, 0.1954531, 
    0.1954544, 0.1954539, 0.1954548, 0.195454, 0.1954541, 0.1954548, 
    0.195454, 0.1954557, 0.1954546, 0.1954568, 0.1954556, 0.1954569, 
    0.1954567, 0.1954571, 0.1954574, 0.1954579, 0.1954588, 0.1954586, 
    0.1954593, 0.1954525, 0.1954528, 0.1954528, 0.1954532, 0.1954535, 
    0.1954541, 0.1954552, 0.1954548, 0.1954555, 0.1954557, 0.1954545, 
    0.1954552, 0.1954531, 0.1954534, 0.1954532, 0.1954525, 0.1954548, 
    0.1954536, 0.195456, 0.1954553, 0.1954574, 0.1954563, 0.1954584, 
    0.1954594, 0.1954603, 0.1954615, 0.195453, 0.1954528, 0.1954532, 
    0.1954539, 0.1954545, 0.1954553, 0.1954554, 0.1954555, 0.195456, 
    0.1954563, 0.1954556, 0.1954564, 0.1954535, 0.195455, 0.1954527, 
    0.1954533, 0.1954538, 0.1954536, 0.1954547, 0.195455, 0.1954561, 
    0.1954555, 0.1954591, 0.1954575, 0.1954623, 0.1954609, 0.1954527, 
    0.195453, 0.1954542, 0.1954537, 0.1954554, 0.1954558, 0.1954561, 
    0.1954566, 0.1954567, 0.1954569, 0.1954565, 0.1954569, 0.1954553, 
    0.195456, 0.1954541, 0.1954545, 0.1954543, 0.1954541, 0.1954548, 
    0.1954556, 0.1954556, 0.1954559, 0.1954565, 0.1954554, 0.1954593, 
    0.1954568, 0.1954534, 0.195454, 0.1954542, 0.1954539, 0.1954557, 
    0.1954551, 0.1954569, 0.1954564, 0.1954573, 0.1954568, 0.1954568, 
    0.1954562, 0.1954559, 0.1954551, 0.1954544, 0.1954539, 0.1954541, 
    0.1954546, 0.1954556, 0.1954567, 0.1954564, 0.1954572, 0.1954552, 
    0.195456, 0.1954557, 0.1954565, 0.1954548, 0.1954562, 0.1954544, 
    0.1954545, 0.195455, 0.1954561, 0.1954563, 0.1954566, 0.1954564, 
    0.1954557, 0.1954556, 0.195455, 0.1954549, 0.1954545, 0.1954542, 
    0.1954545, 0.1954548, 0.1954557, 0.1954565, 0.1954574, 0.1954577, 
    0.1954588, 0.1954578, 0.1954593, 0.195458, 0.1954603, 0.1954563, 
    0.195458, 0.1954551, 0.1954554, 0.1954559, 0.1954572, 0.1954565, 
    0.1954574, 0.1954556, 0.1954546, 0.1954544, 0.195454, 0.1954544, 
    0.1954544, 0.1954548, 0.1954547, 0.1954557, 0.1954551, 0.1954568, 
    0.1954574, 0.1954592, 0.1954604, 0.1954616, 0.1954622, 0.1954624, 
    0.1954624,
  0.1982629, 0.198263, 0.198263, 0.1982631, 0.198263, 0.1982631, 0.1982629, 
    0.198263, 0.198263, 0.1982629, 0.1982632, 0.1982631, 0.1982634, 
    0.1982633, 0.1982636, 0.1982634, 0.1982636, 0.1982636, 0.1982637, 
    0.1982637, 0.1982639, 0.1982637, 0.198264, 0.1982638, 0.1982639, 
    0.1982637, 0.1982631, 0.1982632, 0.1982631, 0.1982631, 0.1982631, 
    0.198263, 0.198263, 0.1982629, 0.1982629, 0.198263, 0.1982631, 0.1982631, 
    0.1982632, 0.1982632, 0.1982633, 0.1982633, 0.1982635, 0.1982634, 
    0.1982637, 0.1982636, 0.1982637, 0.1982636, 0.1982637, 0.1982636, 
    0.1982636, 0.1982635, 0.1982633, 0.1982633, 0.1982631, 0.198263, 
    0.1982629, 0.1982629, 0.1982629, 0.1982629, 0.198263, 0.198263, 
    0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982636, 0.1982637, 0.1982637, 0.1982637, 
    0.1982636, 0.1982637, 0.1982635, 0.1982635, 0.1982632, 0.1982631, 
    0.198263, 0.198263, 0.1982629, 0.198263, 0.1982629, 0.198263, 0.198263, 
    0.198263, 0.1982632, 0.1982631, 0.1982634, 0.1982633, 0.1982636, 
    0.1982635, 0.1982636, 0.1982636, 0.1982637, 0.1982636, 0.1982637, 
    0.1982638, 0.1982637, 0.1982638, 0.1982636, 0.1982637, 0.198263, 
    0.198263, 0.198263, 0.198263, 0.198263, 0.1982629, 0.198263, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982635, 0.1982636, 0.1982635, 0.1982635, 
    0.1982637, 0.1982636, 0.1982638, 0.1982638, 0.1982637, 0.1982638, 
    0.198263, 0.198263, 0.1982629, 0.198263, 0.1982629, 0.1982629, 0.198263, 
    0.1982631, 0.1982631, 0.1982632, 0.1982632, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 
    0.1982636, 0.1982636, 0.1982636, 0.1982638, 0.1982637, 0.1982638, 
    0.1982638, 0.198263, 0.198263, 0.198263, 0.1982631, 0.198263, 0.1982631, 
    0.1982632, 0.1982633, 0.1982633, 0.1982634, 0.1982633, 0.1982633, 
    0.1982634, 0.1982633, 0.1982635, 0.1982633, 0.1982636, 0.1982635, 
    0.1982636, 0.1982636, 0.1982637, 0.1982637, 0.1982638, 0.1982639, 
    0.1982639, 0.198264, 0.1982631, 0.1982631, 0.1982631, 0.1982632, 
    0.1982632, 0.1982633, 0.1982634, 0.1982634, 0.1982635, 0.1982635, 
    0.1982633, 0.1982634, 0.1982632, 0.1982632, 0.1982632, 0.1982631, 
    0.1982634, 0.1982632, 0.1982635, 0.1982634, 0.1982637, 0.1982636, 
    0.1982638, 0.198264, 0.1982641, 0.1982642, 0.1982632, 0.1982631, 
    0.1982632, 0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982635, 
    0.1982635, 0.1982636, 0.1982635, 0.1982636, 0.1982632, 0.1982634, 
    0.1982631, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982634, 
    0.1982635, 0.1982635, 0.1982639, 0.1982637, 0.1982644, 0.1982642, 
    0.1982631, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 
    0.1982634, 0.1982635, 0.1982633, 0.1982633, 0.1982633, 0.1982633, 
    0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982636, 0.1982634, 
    0.198264, 0.1982636, 0.1982632, 0.1982633, 0.1982633, 0.1982633, 
    0.1982635, 0.1982634, 0.1982636, 0.1982636, 0.1982637, 0.1982636, 
    0.1982636, 0.1982636, 0.1982635, 0.1982634, 0.1982633, 0.1982633, 
    0.1982633, 0.1982633, 0.1982635, 0.1982636, 0.1982636, 0.1982637, 
    0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982634, 0.1982636, 
    0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982636, 0.1982636, 
    0.1982636, 0.1982635, 0.1982635, 0.1982634, 0.1982634, 0.1982633, 
    0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982636, 0.1982637, 
    0.1982637, 0.1982639, 0.1982638, 0.198264, 0.1982638, 0.1982641, 
    0.1982636, 0.1982638, 0.1982634, 0.1982635, 0.1982635, 0.1982637, 
    0.1982636, 0.1982637, 0.1982635, 0.1982633, 0.1982633, 0.1982633, 
    0.1982633, 0.1982633, 0.1982634, 0.1982634, 0.1982635, 0.1982634, 
    0.1982636, 0.1982637, 0.1982639, 0.1982641, 0.1982643, 0.1982643, 
    0.1982644, 0.1982644,
  0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.601478, 8.601528, 8.601519, 8.60156, 8.601538, 8.601563, 8.601488, 
    8.60153, 8.601503, 8.601482, 8.601637, 8.601562, 8.60172, 8.601671, 
    8.601795, 8.601711, 8.601812, 8.601793, 8.601851, 8.601835, 8.601907, 
    8.601859, 8.601946, 8.601896, 8.601904, 8.601857, 8.601578, 8.601627, 
    8.601575, 8.601582, 8.601579, 8.601538, 8.601516, 8.601475, 8.601482, 
    8.601513, 8.601584, 8.601562, 8.601623, 8.601622, 8.601689, 8.601659, 
    8.601773, 8.601741, 8.601836, 8.601811, 8.601834, 8.601828, 8.601834, 
    8.6018, 8.601814, 8.601784, 8.601665, 8.601699, 8.601595, 8.60153, 
    8.60149, 8.60146, 8.601465, 8.601473, 8.601513, 8.601553, 8.601583, 
    8.601602, 8.601622, 8.601677, 8.601709, 8.60178, 8.601768, 8.601789, 
    8.60181, 8.601844, 8.601838, 8.601853, 8.601789, 8.601831, 8.601761, 
    8.60178, 8.601623, 8.601567, 8.601542, 8.601521, 8.601468, 8.601504, 
    8.60149, 8.601524, 8.601546, 8.601536, 8.601603, 8.601576, 8.601711, 
    8.601653, 8.601807, 8.60177, 8.601816, 8.601793, 8.601832, 8.601797, 
    8.601859, 8.601871, 8.601863, 8.601898, 8.601795, 8.601834, 8.601536, 
    8.601537, 8.601545, 8.601509, 8.601506, 8.601474, 8.601503, 8.601516, 
    8.601548, 8.601566, 8.601584, 8.601624, 8.601666, 8.601728, 8.601772, 
    8.601803, 8.601785, 8.6018, 8.601783, 8.601774, 8.601867, 8.601814, 
    8.601893, 8.60189, 8.601853, 8.60189, 8.601539, 8.601528, 8.601493, 
    8.601521, 8.601471, 8.601499, 8.601514, 8.601576, 8.60159, 8.601603, 
    8.601628, 8.60166, 8.601716, 8.601766, 8.60181, 8.601808, 8.601809, 
    8.601819, 8.601794, 8.601823, 8.601828, 8.601815, 8.601889, 8.601868, 
    8.601889, 8.601875, 8.601532, 8.601548, 8.60154, 8.601557, 8.601544, 
    8.601598, 8.601614, 8.601689, 8.60166, 8.601708, 8.601665, 8.601672, 
    8.601708, 8.601667, 8.601762, 8.601696, 8.601819, 8.601752, 8.601823, 
    8.60181, 8.601831, 8.60185, 8.601873, 8.601916, 8.601907, 8.601943, 
    8.601574, 8.601596, 8.601594, 8.601617, 8.601634, 8.601671, 8.60173, 
    8.601708, 8.601749, 8.601758, 8.601695, 8.601733, 8.60161, 8.601629, 
    8.601619, 8.601575, 8.601712, 8.601642, 8.601773, 8.601735, 8.601847, 
    8.60179, 8.601901, 8.601946, 8.601993, 8.602042, 8.601608, 8.601593, 
    8.60162, 8.601656, 8.601691, 8.601737, 8.601743, 8.60175, 8.601773, 
    8.601792, 8.601752, 8.601797, 8.601632, 8.601719, 8.601587, 8.601625, 
    8.601654, 8.601643, 8.601707, 8.601721, 8.601781, 8.60175, 8.601934, 
    8.601852, 8.602083, 8.602018, 8.601588, 8.601608, 8.601678, 8.601645, 
    8.601741, 8.601764, 8.601784, 8.601808, 8.60181, 8.601825, 8.601801, 
    8.601824, 8.601737, 8.601776, 8.60167, 8.601696, 8.601685, 8.601671, 
    8.601711, 8.601753, 8.601755, 8.601768, 8.601804, 8.601741, 8.601943, 
    8.601816, 8.60163, 8.601667, 8.601674, 8.60166, 8.601762, 8.601725, 
    8.601825, 8.601798, 8.601842, 8.60182, 8.601817, 8.601789, 8.60177, 
    8.601726, 8.60169, 8.601662, 8.601668, 8.601699, 8.601756, 8.60181, 
    8.601798, 8.601839, 8.601733, 8.601777, 8.60176, 8.601805, 8.601707, 
    8.601788, 8.601686, 8.601696, 8.601724, 8.601779, 8.601793, 8.601807, 
    8.601798, 8.601758, 8.601751, 8.601724, 8.601715, 8.601694, 8.601676, 
    8.601692, 8.601709, 8.601758, 8.601802, 8.60185, 8.601862, 8.601915, 
    8.601871, 8.601943, 8.601879, 8.601992, 8.601793, 8.601879, 8.601726, 
    8.601742, 8.601771, 8.601841, 8.601805, 8.601848, 8.601751, 8.6017, 
    8.601687, 8.601664, 8.601688, 8.601686, 8.60171, 8.601703, 8.60176, 
    8.601729, 8.601816, 8.601848, 8.601938, 8.601994, 8.602051, 8.602076, 
    8.602084, 8.602087 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.955336e-15, 3.95574e-15, 3.955663e-15, 3.955985e-15, 3.955809e-15, 
    3.956018e-15, 3.955421e-15, 3.955753e-15, 3.955543e-15, 3.955377e-15, 
    3.9566e-15, 3.956e-15, 3.957258e-15, 3.956869e-15, 3.957858e-15, 
    3.957193e-15, 3.957994e-15, 3.957847e-15, 3.958309e-15, 3.958177e-15, 
    3.958753e-15, 3.95837e-15, 3.959065e-15, 3.958666e-15, 3.958725e-15, 
    3.958356e-15, 3.956128e-15, 3.956523e-15, 3.956103e-15, 3.95616e-15, 
    3.956136e-15, 3.95581e-15, 3.95564e-15, 3.95531e-15, 3.955372e-15, 
    3.955617e-15, 3.956186e-15, 3.955997e-15, 3.956487e-15, 3.956476e-15, 
    3.957016e-15, 3.956772e-15, 3.957687e-15, 3.957428e-15, 3.958183e-15, 
    3.957992e-15, 3.958173e-15, 3.958119e-15, 3.958173e-15, 3.957893e-15, 
    3.958013e-15, 3.957769e-15, 3.956816e-15, 3.957093e-15, 3.956263e-15, 
    3.955753e-15, 3.955434e-15, 3.955203e-15, 3.955235e-15, 3.955296e-15, 
    3.955618e-15, 3.955929e-15, 3.956164e-15, 3.956319e-15, 3.956474e-15, 
    3.956922e-15, 3.957177e-15, 3.957735e-15, 3.957641e-15, 3.957806e-15, 
    3.957973e-15, 3.958245e-15, 3.958201e-15, 3.958319e-15, 3.957806e-15, 
    3.958145e-15, 3.957586e-15, 3.957738e-15, 3.956489e-15, 3.95605e-15, 
    3.95584e-15, 3.955676e-15, 3.95526e-15, 3.955546e-15, 3.955433e-15, 
    3.955709e-15, 3.95588e-15, 3.955796e-15, 3.956324e-15, 3.956117e-15, 
    3.957192e-15, 3.956729e-15, 3.957954e-15, 3.957661e-15, 3.958025e-15, 
    3.95784e-15, 3.958154e-15, 3.957872e-15, 3.958365e-15, 3.95847e-15, 
    3.958398e-15, 3.958684e-15, 3.957855e-15, 3.95817e-15, 3.955793e-15, 
    3.955806e-15, 3.955872e-15, 3.955582e-15, 3.955565e-15, 3.955307e-15, 
    3.955539e-15, 3.955636e-15, 3.955892e-15, 3.956039e-15, 3.95618e-15, 
    3.956491e-15, 3.956835e-15, 3.957324e-15, 3.95768e-15, 3.957917e-15, 
    3.957773e-15, 3.9579e-15, 3.957757e-15, 3.957692e-15, 3.958429e-15, 
    3.958012e-15, 3.958643e-15, 3.958609e-15, 3.958321e-15, 3.958613e-15, 
    3.955816e-15, 3.955737e-15, 3.955457e-15, 3.955676e-15, 3.95528e-15, 
    3.955498e-15, 3.955622e-15, 3.956116e-15, 3.956231e-15, 3.956329e-15, 
    3.95653e-15, 3.956784e-15, 3.957229e-15, 3.957621e-15, 3.957984e-15, 
    3.957958e-15, 3.957967e-15, 3.958045e-15, 3.957847e-15, 3.958078e-15, 
    3.958114e-15, 3.958016e-15, 3.958604e-15, 3.958436e-15, 3.958608e-15, 
    3.958499e-15, 3.955764e-15, 3.955897e-15, 3.955825e-15, 3.95596e-15, 
    3.955862e-15, 3.956287e-15, 3.956415e-15, 3.957019e-15, 3.956778e-15, 
    3.95717e-15, 3.95682e-15, 3.95688e-15, 3.957171e-15, 3.95684e-15, 
    3.957595e-15, 3.957073e-15, 3.958048e-15, 3.957515e-15, 3.958081e-15, 
    3.957982e-15, 3.958148e-15, 3.958294e-15, 3.958483e-15, 3.958824e-15, 
    3.958746e-15, 3.959035e-15, 3.956099e-15, 3.956269e-15, 3.95626e-15, 
    3.956442e-15, 3.956576e-15, 3.956872e-15, 3.957343e-15, 3.957168e-15, 
    3.957495e-15, 3.957559e-15, 3.957065e-15, 3.957364e-15, 3.956388e-15, 
    3.95654e-15, 3.956453e-15, 3.956109e-15, 3.957201e-15, 3.956637e-15, 
    3.957684e-15, 3.957379e-15, 3.958273e-15, 3.957823e-15, 3.958702e-15, 
    3.959065e-15, 3.959432e-15, 3.959833e-15, 3.956369e-15, 3.956252e-15, 
    3.956465e-15, 3.956751e-15, 3.957032e-15, 3.957397e-15, 3.957437e-15, 
    3.957504e-15, 3.957684e-15, 3.957833e-15, 3.95752e-15, 3.957871e-15, 
    3.956565e-15, 3.957252e-15, 3.956203e-15, 3.956512e-15, 3.956737e-15, 
    3.956643e-15, 3.957149e-15, 3.957266e-15, 3.957743e-15, 3.9575e-15, 
    3.958971e-15, 3.958318e-15, 3.960156e-15, 3.959638e-15, 3.95621e-15, 
    3.95637e-15, 3.956923e-15, 3.956661e-15, 3.957424e-15, 3.95761e-15, 
    3.957766e-15, 3.957957e-15, 3.957981e-15, 3.958095e-15, 3.957908e-15, 
    3.95809e-15, 3.957398e-15, 3.957708e-15, 3.956866e-15, 3.957067e-15, 
    3.956976e-15, 3.956872e-15, 3.957192e-15, 3.957524e-15, 3.95754e-15, 
    3.957645e-15, 3.957927e-15, 3.957427e-15, 3.95904e-15, 3.958028e-15, 
    3.956545e-15, 3.956844e-15, 3.956896e-15, 3.956779e-15, 3.957591e-15, 
    3.957296e-15, 3.958093e-15, 3.957879e-15, 3.958233e-15, 3.958056e-15, 
    3.95803e-15, 3.957805e-15, 3.957664e-15, 3.957307e-15, 3.95702e-15, 
    3.956797e-15, 3.95685e-15, 3.957095e-15, 3.957546e-15, 3.95798e-15, 
    3.957884e-15, 3.958206e-15, 3.957368e-15, 3.957715e-15, 3.957578e-15, 
    3.957936e-15, 3.957161e-15, 3.957796e-15, 3.956996e-15, 3.957068e-15, 
    3.95729e-15, 3.957733e-15, 3.957843e-15, 3.957947e-15, 3.957884e-15, 
    3.957559e-15, 3.95751e-15, 3.957286e-15, 3.957221e-15, 3.957053e-15, 
    3.956911e-15, 3.957039e-15, 3.957171e-15, 3.957563e-15, 3.957911e-15, 
    3.958295e-15, 3.958392e-15, 3.958821e-15, 3.958461e-15, 3.959044e-15, 
    3.958531e-15, 3.959429e-15, 3.957845e-15, 3.958532e-15, 3.957302e-15, 
    3.957437e-15, 3.957671e-15, 3.958226e-15, 3.957935e-15, 3.958279e-15, 
    3.957509e-15, 3.957099e-15, 3.957004e-15, 3.956809e-15, 3.957008e-15, 
    3.956992e-15, 3.957183e-15, 3.957122e-15, 3.957576e-15, 3.957332e-15, 
    3.958027e-15, 3.958279e-15, 3.959002e-15, 3.959441e-15, 3.959902e-15, 
    3.960102e-15, 3.960164e-15, 3.960189e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.791278, 9.839125, 9.82981, 9.868475, 9.847019, 9.872292, 9.800964, 
    9.841029, 9.815439, 9.795576, 9.942685, 9.870175, 10.01833, 9.971833, 
    10.08889, 10.01109, 10.10462, 10.08664, 10.14082, 10.12528, 10.19479, 
    10.148, 10.23093, 10.1836, 10.191, 10.14646, 9.884735, 9.933641, 
    9.881844, 9.888807, 9.885681, 9.847465, 9.828105, 9.787623, 9.794964, 
    9.824698, 9.891939, 9.869296, 9.926414, 9.925121, 9.988953, 9.96014, 
    10.06781, 10.03713, 10.12593, 10.10355, 10.12488, 10.11841, 10.12496, 
    10.09216, 10.1062, 10.07736, 9.965533, 9.998322, 9.900737, 9.841975, 
    9.80272, 9.774928, 9.778853, 9.786342, 9.824873, 9.861181, 9.888589, 
    9.906887, 9.924935, 9.979709, 10.00876, 10.07402, 10.06222, 10.08221, 
    10.10133, 10.13348, 10.12818, 10.14236, 10.08168, 10.12199, 10.0555, 
    10.07366, 9.929865, 9.875401, 9.852093, 9.831601, 9.781874, 9.816198, 
    9.802659, 9.834886, 9.855401, 9.84525, 9.907387, 9.883331, 10.01049, 
    9.955591, 10.0991, 10.06464, 10.10736, 10.08555, 10.12295, 10.08928, 
    10.14764, 10.16038, 10.15167, 10.18513, 10.08742, 10.12488, 9.844967, 
    9.846622, 9.854333, 9.820466, 9.818396, 9.787423, 9.814978, 9.826728, 
    9.856589, 9.874181, 9.890765, 9.927289, 9.968184, 10.02554, 10.06687, 
    10.09463, 10.0776, 10.09264, 10.07583, 10.06796, 10.15561, 10.10634, 
    10.18031, 10.17621, 10.1427, 10.17667, 9.847784, 9.838262, 9.805252, 
    9.831079, 9.784053, 9.810361, 9.825509, 9.883838, 9.896539, 9.908332, 
    9.931643, 9.961614, 10.01433, 10.06033, 10.10244, 10.09935, 10.10044, 
    10.10986, 10.08653, 10.11369, 10.11826, 10.10633, 10.17566, 10.15582, 
    10.17612, 10.1632, 9.841356, 9.857384, 9.848722, 9.865016, 9.853536, 
    9.904096, 9.919223, 9.990195, 9.961024, 10.00747, 9.965734, 9.973124, 
    10.009, 9.967986, 10.05779, 9.99686, 10.11023, 10.04919, 10.11406, 
    10.10226, 10.1218, 10.13933, 10.1614, 10.2022, 10.19274, 10.22692, 
    9.8811, 9.901634, 9.899822, 9.921335, 9.937264, 9.971843, 10.02746, 
    10.00652, 10.04498, 10.05271, 9.994293, 10.03014, 9.915389, 9.933877, 
    9.922864, 9.882721, 10.01135, 9.94521, 10.06755, 10.03156, 10.13683, 
    10.0844, 10.18754, 10.23184, 10.27362, 10.3226, 9.912848, 9.898884, 
    9.923894, 9.95857, 9.990801, 10.03376, 10.03816, 10.04622, 10.06712, 
    10.08472, 10.04877, 10.08913, 9.938175, 10.0171, 9.89361, 9.9307, 
    9.956522, 9.945186, 10.00413, 10.01806, 10.07477, 10.04543, 10.2209, 
    10.14303, 10.35997, 10.29907, 9.894008, 9.912799, 9.978378, 9.947141, 
    10.03663, 10.05873, 10.07672, 10.09975, 10.10224, 10.1159, 10.09352, 
    10.11501, 10.03385, 10.07007, 9.970864, 9.994956, 9.983867, 9.971715, 
    10.00925, 10.04934, 10.05019, 10.06307, 10.09943, 10.03699, 10.23099, 
    10.11092, 9.933315, 9.969628, 9.974814, 9.960734, 10.05651, 10.02174, 
    10.11557, 10.09015, 10.13181, 10.1111, 10.10805, 10.08149, 10.06498, 
    10.02334, 9.989533, 9.962775, 9.968992, 9.998401, 10.0518, 10.10247, 
    10.09135, 10.12864, 10.03012, 10.07136, 10.05541, 10.09703, 10.00597, 
    10.0835, 9.986213, 9.994718, 10.02106, 10.07417, 10.08593, 10.09852, 
    10.09075, 10.05315, 10.047, 10.02041, 10.01308, 9.992865, 9.976148, 
    9.991423, 10.00748, 10.05316, 10.09445, 10.13958, 10.15064, 10.20357, 
    10.16047, 10.23166, 10.17113, 10.27604, 10.088, 10.16934, 10.02225, 
    10.03803, 10.06662, 10.13237, 10.09684, 10.1384, 10.04676, 9.999419, 
    9.987186, 9.964402, 9.987708, 9.985811, 10.00814, 10.00096, 10.05468, 
    10.0258, 10.10798, 10.13807, 10.22334, 10.27583, 10.32943, 10.35314, 
    10.36037, 10.36339 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  1.751983e-09, 1.731532e-09, 1.735468e-09, 1.71926e-09, 1.728211e-09, 
    1.717655e-09, 1.747796e-09, 1.730731e-09, 1.741584e-09, 1.750121e-09, 
    1.688698e-09, 1.718544e-09, 1.658823e-09, 1.677032e-09, 1.632061e-09, 
    1.66163e-09, 1.626231e-09, 1.632899e-09, 1.613001e-09, 1.61865e-09, 
    1.593744e-09, 1.610408e-09, 1.581144e-09, 1.597691e-09, 1.595079e-09, 
    1.610964e-09, 1.712448e-09, 1.692354e-09, 1.713655e-09, 1.710754e-09, 
    1.712054e-09, 1.728026e-09, 1.736194e-09, 1.753567e-09, 1.750386e-09, 
    1.737639e-09, 1.709454e-09, 1.718912e-09, 1.695281e-09, 1.695807e-09, 
    1.670273e-09, 1.681685e-09, 1.63995e-09, 1.65159e-09, 1.618413e-09, 
    1.626626e-09, 1.618797e-09, 1.621162e-09, 1.618766e-09, 1.630846e-09, 
    1.625647e-09, 1.636361e-09, 1.679536e-09, 1.666602e-09, 1.70581e-09, 
    1.730335e-09, 1.74704e-09, 1.759102e-09, 1.757386e-09, 1.754125e-09, 
    1.737565e-09, 1.722293e-09, 1.710843e-09, 1.703273e-09, 1.695883e-09, 
    1.673919e-09, 1.662533e-09, 1.637617e-09, 1.642056e-09, 1.634551e-09, 
    1.627447e-09, 1.615665e-09, 1.617592e-09, 1.612444e-09, 1.634748e-09, 
    1.619854e-09, 1.644595e-09, 1.63775e-09, 1.693887e-09, 1.71635e-09, 
    1.72609e-09, 1.73471e-09, 1.75607e-09, 1.74126e-09, 1.747067e-09, 
    1.73332e-09, 1.724703e-09, 1.728953e-09, 1.703067e-09, 1.713033e-09, 
    1.661863e-09, 1.683506e-09, 1.628272e-09, 1.641143e-09, 1.625219e-09, 
    1.633304e-09, 1.619501e-09, 1.631912e-09, 1.610537e-09, 1.60596e-09, 
    1.609085e-09, 1.597148e-09, 1.632606e-09, 1.618797e-09, 1.729073e-09, 
    1.728378e-09, 1.725148e-09, 1.73944e-09, 1.740322e-09, 1.753655e-09, 
    1.741781e-09, 1.736776e-09, 1.724206e-09, 1.716861e-09, 1.709939e-09, 
    1.694926e-09, 1.678482e-09, 1.656041e-09, 1.640302e-09, 1.629925e-09, 
    1.636272e-09, 1.630666e-09, 1.636935e-09, 1.639891e-09, 1.607672e-09, 
    1.625599e-09, 1.598854e-09, 1.60031e-09, 1.612322e-09, 1.600145e-09, 
    1.72789e-09, 1.731894e-09, 1.74595e-09, 1.73493e-09, 1.75512e-09, 
    1.743758e-09, 1.737295e-09, 1.712824e-09, 1.707544e-09, 1.70268e-09, 
    1.693156e-09, 1.681097e-09, 1.660372e-09, 1.642769e-09, 1.627036e-09, 
    1.628178e-09, 1.627776e-09, 1.624301e-09, 1.632937e-09, 1.622892e-09, 
    1.621218e-09, 1.625601e-09, 1.600505e-09, 1.607592e-09, 1.600341e-09, 
    1.604947e-09, 1.730591e-09, 1.723875e-09, 1.727497e-09, 1.720699e-09, 
    1.725483e-09, 1.704426e-09, 1.698217e-09, 1.669787e-09, 1.681333e-09, 
    1.663035e-09, 1.679455e-09, 1.676521e-09, 1.662445e-09, 1.678559e-09, 
    1.64373e-09, 1.667176e-09, 1.624166e-09, 1.646997e-09, 1.622757e-09, 
    1.627103e-09, 1.61992e-09, 1.613543e-09, 1.605594e-09, 1.591138e-09, 
    1.594461e-09, 1.582526e-09, 1.713965e-09, 1.70544e-09, 1.706186e-09, 
    1.697352e-09, 1.690879e-09, 1.677027e-09, 1.6553e-09, 1.663401e-09, 
    1.648592e-09, 1.645652e-09, 1.668176e-09, 1.654271e-09, 1.699784e-09, 
    1.692254e-09, 1.696728e-09, 1.713289e-09, 1.661527e-09, 1.687675e-09, 
    1.640044e-09, 1.653724e-09, 1.614449e-09, 1.633736e-09, 1.596297e-09, 
    1.58083e-09, 1.566554e-09, 1.550205e-09, 1.700824e-09, 1.706574e-09, 
    1.696307e-09, 1.682315e-09, 1.669547e-09, 1.652883e-09, 1.651197e-09, 
    1.648121e-09, 1.640207e-09, 1.633614e-09, 1.647151e-09, 1.631969e-09, 
    1.690518e-09, 1.659297e-09, 1.708759e-09, 1.693542e-09, 1.683133e-09, 
    1.687683e-09, 1.664332e-09, 1.658927e-09, 1.637335e-09, 1.648423e-09, 
    1.584619e-09, 1.612203e-09, 1.537991e-09, 1.55801e-09, 1.708593e-09, 
    1.700844e-09, 1.674441e-09, 1.686895e-09, 1.651783e-09, 1.643373e-09, 
    1.636602e-09, 1.62803e-09, 1.62711e-09, 1.622082e-09, 1.630339e-09, 
    1.622406e-09, 1.652848e-09, 1.639098e-09, 1.677415e-09, 1.667918e-09, 
    1.672273e-09, 1.677078e-09, 1.662341e-09, 1.646936e-09, 1.64661e-09, 
    1.641735e-09, 1.628159e-09, 1.651643e-09, 1.58113e-09, 1.623918e-09, 
    1.692478e-09, 1.67791e-09, 1.67585e-09, 1.681447e-09, 1.644212e-09, 
    1.657503e-09, 1.622204e-09, 1.631589e-09, 1.61627e-09, 1.623845e-09, 
    1.624965e-09, 1.634817e-09, 1.641013e-09, 1.656889e-09, 1.670044e-09, 
    1.680633e-09, 1.678158e-09, 1.66657e-09, 1.646003e-09, 1.627027e-09, 
    1.631145e-09, 1.617424e-09, 1.654277e-09, 1.638613e-09, 1.644631e-09, 
    1.629036e-09, 1.663618e-09, 1.634075e-09, 1.671349e-09, 1.66801e-09, 
    1.657769e-09, 1.637562e-09, 1.63316e-09, 1.628488e-09, 1.631368e-09, 
    1.645488e-09, 1.647825e-09, 1.658016e-09, 1.660853e-09, 1.668736e-09, 
    1.675321e-09, 1.669302e-09, 1.66303e-09, 1.645482e-09, 1.629995e-09, 
    1.613453e-09, 1.609457e-09, 1.590663e-09, 1.605928e-09, 1.580898e-09, 
    1.602126e-09, 1.565744e-09, 1.632396e-09, 1.602759e-09, 1.657306e-09, 
    1.651244e-09, 1.640397e-09, 1.616069e-09, 1.629108e-09, 1.61388e-09, 
    1.647917e-09, 1.666174e-09, 1.670966e-09, 1.679985e-09, 1.670761e-09, 
    1.671507e-09, 1.662771e-09, 1.665568e-09, 1.644906e-09, 1.655937e-09, 
    1.624994e-09, 1.613999e-09, 1.583768e-09, 1.565809e-09, 1.547955e-09, 
    1.540206e-09, 1.537863e-09, 1.536886e-09 ;

 W_SCALAR =
  0.6202525, 0.6219193, 0.6215954, 0.6229389, 0.6221938, 0.6230733, 
    0.6205905, 0.6219854, 0.6210951, 0.6204026, 0.6255435, 0.6229988, 
    0.6281826, 0.6265627, 0.6306291, 0.6279306, 0.6311727, 0.6305513, 
    0.6324207, 0.6318853, 0.6342741, 0.6326677, 0.6355109, 0.6338906, 
    0.6341442, 0.6326147, 0.6235112, 0.6252269, 0.6234095, 0.6236542, 
    0.6235444, 0.6222091, 0.6215359, 0.620125, 0.6203812, 0.6214174, 
    0.6237643, 0.622968, 0.6249742, 0.6249289, 0.6271598, 0.6261543, 
    0.6298996, 0.628836, 0.6319077, 0.6311357, 0.6318714, 0.6316484, 
    0.6318743, 0.630742, 0.6312273, 0.6302305, 0.6263427, 0.6274862, 
    0.6240734, 0.6220182, 0.6206517, 0.6196815, 0.6198187, 0.6200802, 
    0.6214235, 0.6226856, 0.6236467, 0.6242894, 0.6249224, 0.6268372, 
    0.6278497, 0.6301146, 0.6297061, 0.6303981, 0.6310589, 0.6321678, 
    0.6319853, 0.6324736, 0.6303799, 0.6317717, 0.6294733, 0.6301023, 
    0.6250946, 0.6231828, 0.6223698, 0.6216577, 0.6199241, 0.6211215, 
    0.6206496, 0.621772, 0.6224849, 0.6221323, 0.624307, 0.6234618, 
    0.6279097, 0.6259952, 0.6309819, 0.6297899, 0.6312674, 0.6305137, 
    0.6318049, 0.6306428, 0.6326554, 0.6330933, 0.632794, 0.6339431, 
    0.6305784, 0.6318715, 0.6221224, 0.6221799, 0.6224478, 0.6212701, 
    0.621198, 0.620118, 0.621079, 0.6214881, 0.6225262, 0.6231399, 0.6237231, 
    0.6250048, 0.6264352, 0.6284332, 0.6298673, 0.6308278, 0.6302388, 
    0.6307588, 0.6301776, 0.629905, 0.6329292, 0.6312318, 0.6337779, 
    0.6336371, 0.6324853, 0.633653, 0.6222203, 0.6218894, 0.6207401, 
    0.6216395, 0.6200003, 0.6209181, 0.6214456, 0.6234795, 0.623926, 
    0.6243401, 0.6251574, 0.6262058, 0.6280434, 0.6296406, 0.6310973, 
    0.6309906, 0.6310282, 0.6313535, 0.6305477, 0.6314858, 0.6316431, 
    0.6312316, 0.6336183, 0.6329368, 0.6336342, 0.6331905, 0.6219969, 
    0.6225537, 0.6222529, 0.6228185, 0.6224201, 0.6241913, 0.6247219, 
    0.627203, 0.6261852, 0.6278048, 0.6263497, 0.6266077, 0.6278576, 
    0.6264284, 0.6295527, 0.6274352, 0.6313661, 0.629254, 0.6314984, 
    0.6310911, 0.6317654, 0.6323692, 0.6331283, 0.6345283, 0.6342042, 
    0.6353742, 0.6233833, 0.6241049, 0.6240414, 0.6247962, 0.6253542, 
    0.626563, 0.6285001, 0.6277719, 0.6291085, 0.6293766, 0.627346, 
    0.6285931, 0.6245877, 0.6252354, 0.6248497, 0.6234403, 0.6279398, 
    0.6256321, 0.6298909, 0.6286426, 0.6322831, 0.6304737, 0.6340258, 
    0.6355419, 0.6369673, 0.6386315, 0.6244985, 0.6240084, 0.6248859, 
    0.6260993, 0.6272243, 0.6287188, 0.6288716, 0.6291514, 0.629876, 
    0.6304849, 0.6292399, 0.6306375, 0.6253857, 0.62814, 0.6238231, 
    0.6251242, 0.6260278, 0.6256315, 0.6276887, 0.6281732, 0.6301407, 
    0.6291239, 0.6351679, 0.6324967, 0.6398973, 0.6378328, 0.6238372, 
    0.6244969, 0.626791, 0.6256998, 0.6288185, 0.6295853, 0.6302083, 
    0.6310045, 0.6310904, 0.6315619, 0.6307892, 0.6315314, 0.628722, 
    0.629978, 0.6265289, 0.627369, 0.6269826, 0.6265586, 0.6278669, 
    0.6292595, 0.6292892, 0.6297355, 0.6309927, 0.6288311, 0.6355124, 
    0.6313896, 0.6252159, 0.6264855, 0.6266667, 0.6261751, 0.6295084, 
    0.6283014, 0.6315504, 0.6306729, 0.6321104, 0.6313962, 0.6312912, 
    0.6303734, 0.6298018, 0.6283568, 0.6271801, 0.6262464, 0.6264636, 
    0.627489, 0.6293446, 0.6310982, 0.6307142, 0.6320012, 0.6285926, 
    0.6300228, 0.6294701, 0.6309106, 0.6277526, 0.6304424, 0.6270644, 
    0.6273608, 0.6282774, 0.6301197, 0.630527, 0.6309618, 0.6306935, 
    0.6293917, 0.6291783, 0.6282551, 0.6280002, 0.6272963, 0.6267133, 
    0.627246, 0.6278052, 0.6293923, 0.6308212, 0.6323777, 0.6327584, 
    0.6345748, 0.6330964, 0.6355354, 0.6334621, 0.6370491, 0.6305981, 
    0.633401, 0.6283191, 0.6288673, 0.6298586, 0.6321295, 0.6309038, 
    0.6323372, 0.62917, 0.6275244, 0.6270983, 0.6263032, 0.6271165, 
    0.6270504, 0.6278283, 0.6275784, 0.629445, 0.6284425, 0.6312885, 
    0.6323259, 0.6352516, 0.6370425, 0.6388631, 0.6396663, 0.6399106, 
    0.6400128,
  0.5451502, 0.5471774, 0.5467834, 0.5484173, 0.547511, 0.5485807, 0.5455613, 
    0.5472579, 0.5461749, 0.5453327, 0.5515841, 0.5484901, 0.5547913, 
    0.5528225, 0.5577639, 0.5544852, 0.5584242, 0.5576693, 0.5599402, 
    0.5592899, 0.5621916, 0.5602402, 0.5636935, 0.5617257, 0.5620338, 
    0.5601758, 0.549113, 0.5511992, 0.5489894, 0.549287, 0.5491534, 
    0.5475299, 0.5467113, 0.5449951, 0.5453067, 0.5465671, 0.5494208, 
    0.5484525, 0.5508916, 0.5508366, 0.5535483, 0.5523261, 0.5568776, 
    0.5555851, 0.5593171, 0.5583793, 0.559273, 0.559002, 0.5592766, 0.557901, 
    0.5584905, 0.5572796, 0.5525551, 0.553945, 0.5497966, 0.5472978, 
    0.5456358, 0.5444556, 0.5446225, 0.5449407, 0.5465745, 0.5481091, 
    0.5492778, 0.5500591, 0.5508286, 0.5531564, 0.5543867, 0.5571389, 
    0.5566424, 0.5574833, 0.558286, 0.559633, 0.5594113, 0.5600046, 0.557461, 
    0.5591519, 0.5563595, 0.5571237, 0.5510384, 0.5487137, 0.5477253, 
    0.5468592, 0.5447508, 0.5462071, 0.5456332, 0.5469981, 0.547865, 
    0.5474364, 0.5500805, 0.549053, 0.5544596, 0.5521328, 0.5581924, 
    0.5567443, 0.5585393, 0.5576235, 0.5591923, 0.5577804, 0.5602253, 
    0.5607573, 0.5603938, 0.5617895, 0.5577022, 0.5592731, 0.5474244, 
    0.5474943, 0.54782, 0.5463879, 0.5463002, 0.5449865, 0.5461554, 0.546653, 
    0.5479152, 0.5486616, 0.5493707, 0.5509289, 0.5526676, 0.5550959, 
    0.5568382, 0.5580051, 0.5572896, 0.5579214, 0.5572152, 0.5568841, 
    0.560558, 0.5584961, 0.5615888, 0.5614178, 0.5600188, 0.5614371, 
    0.5475434, 0.547141, 0.5457432, 0.5468372, 0.5448434, 0.5459598, 
    0.5466014, 0.5490746, 0.5496174, 0.5501208, 0.5511143, 0.5523887, 
    0.5546221, 0.5565629, 0.5583326, 0.558203, 0.5582486, 0.5586438, 
    0.5576649, 0.5588045, 0.5589957, 0.5584958, 0.5613949, 0.5605671, 
    0.5614141, 0.5608752, 0.5472717, 0.5479488, 0.547583, 0.5482708, 
    0.5477863, 0.5499399, 0.5505852, 0.5536008, 0.5523636, 0.5543321, 
    0.5525637, 0.5528772, 0.5543966, 0.5526592, 0.5564561, 0.5538831, 
    0.5586592, 0.5560933, 0.5588199, 0.558325, 0.5591442, 0.5598776, 
    0.5607998, 0.5625002, 0.5621065, 0.5635274, 0.5489576, 0.5498349, 
    0.5497576, 0.5506752, 0.5513536, 0.5528229, 0.555177, 0.5542921, 
    0.5559162, 0.5562421, 0.5537745, 0.5552901, 0.5504218, 0.5512093, 
    0.5507404, 0.5490268, 0.5544962, 0.5516915, 0.5568669, 0.5553502, 
    0.5597731, 0.557575, 0.5618898, 0.5637314, 0.565462, 0.5674829, 
    0.5503134, 0.5497175, 0.5507843, 0.5522594, 0.5536266, 0.5554428, 
    0.5556284, 0.5559684, 0.5568488, 0.5575886, 0.556076, 0.557774, 
    0.5513922, 0.5547394, 0.5494923, 0.5510741, 0.5521724, 0.5516906, 
    0.5541909, 0.5547797, 0.5571705, 0.555935, 0.5632771, 0.5600327, 
    0.5690195, 0.5665131, 0.5495093, 0.5503113, 0.5531, 0.5517737, 0.5555639, 
    0.5564956, 0.5572525, 0.5582199, 0.5583242, 0.558897, 0.5579582, 
    0.5588599, 0.5554466, 0.5569727, 0.5527813, 0.5538025, 0.5533328, 
    0.5528175, 0.5544074, 0.5560999, 0.5561358, 0.5566782, 0.558206, 
    0.5555792, 0.5636958, 0.5586881, 0.5511855, 0.5527288, 0.552949, 
    0.5523514, 0.5564022, 0.5549356, 0.558883, 0.557817, 0.5595633, 
    0.5586957, 0.5585681, 0.5574532, 0.5567587, 0.5550029, 0.5535729, 
    0.552438, 0.552702, 0.5539483, 0.5562033, 0.5583338, 0.5578673, 
    0.5594306, 0.5552893, 0.5570272, 0.5563558, 0.5581058, 0.5542686, 
    0.5575374, 0.5534322, 0.5537925, 0.5549064, 0.5571451, 0.5576397, 
    0.558168, 0.557842, 0.5562605, 0.5560012, 0.5548793, 0.5545695, 0.553714, 
    0.5530055, 0.5536529, 0.5543326, 0.5562611, 0.5579973, 0.5598881, 
    0.5603505, 0.5625569, 0.5607613, 0.5637237, 0.5612058, 0.5655618, 
    0.5577263, 0.5611313, 0.554957, 0.5556232, 0.5568277, 0.5595868, 
    0.5580976, 0.559839, 0.555991, 0.5539914, 0.5534735, 0.5525071, 
    0.5534956, 0.5534152, 0.5543606, 0.5540568, 0.5563251, 0.5551071, 
    0.558565, 0.5598251, 0.5633786, 0.5655534, 0.5677639, 0.568739, 
    0.5690356, 0.5691596,
  0.5138803, 0.5161285, 0.5156915, 0.5175039, 0.5164986, 0.5176852, 
    0.5143362, 0.5162178, 0.5150167, 0.5140826, 0.5210179, 0.5175847, 
    0.5245786, 0.5223925, 0.5278802, 0.5242386, 0.5286138, 0.527775, 
    0.5302982, 0.5295756, 0.5328008, 0.5306317, 0.5344706, 0.5322828, 
    0.5326253, 0.5305601, 0.5182757, 0.5205908, 0.5181385, 0.5184688, 
    0.5183206, 0.5165194, 0.5156115, 0.5137082, 0.5140538, 0.5154516, 
    0.5186173, 0.5175429, 0.5202493, 0.5201882, 0.5231983, 0.5218415, 
    0.5268955, 0.52546, 0.5296058, 0.5285639, 0.5295569, 0.5292557, 
    0.5295608, 0.5280325, 0.5286874, 0.5273421, 0.5220957, 0.5236388, 
    0.5190342, 0.5162621, 0.5144187, 0.5131101, 0.5132952, 0.5136479, 
    0.5154597, 0.5171619, 0.5184585, 0.5193255, 0.5201795, 0.5227633, 
    0.5241293, 0.5271858, 0.5266343, 0.5275684, 0.5284601, 0.5299569, 
    0.5297106, 0.5303699, 0.5275436, 0.5294223, 0.5263201, 0.527169, 
    0.5204124, 0.5178328, 0.5167363, 0.5157755, 0.5134374, 0.5150523, 
    0.5144159, 0.5159296, 0.5168912, 0.5164157, 0.5193492, 0.5182091, 
    0.5242103, 0.521627, 0.5283561, 0.5267475, 0.5287415, 0.5277241, 
    0.5294672, 0.5278986, 0.5306152, 0.5312064, 0.5308024, 0.5323536, 
    0.5278116, 0.529557, 0.5164024, 0.51648, 0.5168412, 0.5152528, 0.5151556, 
    0.5136988, 0.514995, 0.5155469, 0.5169469, 0.5177749, 0.5185617, 
    0.5202907, 0.5222206, 0.5249166, 0.5268518, 0.5281481, 0.5273532, 
    0.528055, 0.5272706, 0.5269027, 0.5309849, 0.5286936, 0.5321306, 
    0.5319405, 0.5303856, 0.5319619, 0.5165344, 0.516088, 0.5145378, 
    0.5157511, 0.5135401, 0.514778, 0.5154896, 0.5182331, 0.5188354, 
    0.5193939, 0.5204965, 0.521911, 0.5243906, 0.526546, 0.528512, 0.528368, 
    0.5284187, 0.5288578, 0.5277701, 0.5290363, 0.5292488, 0.5286932, 
    0.5319151, 0.530995, 0.5319365, 0.5313374, 0.5162331, 0.5169841, 
    0.5165783, 0.5173414, 0.5168039, 0.5191933, 0.5199093, 0.5232567, 
    0.5218832, 0.5240686, 0.5221052, 0.5224532, 0.5241402, 0.5222113, 
    0.5264274, 0.5235701, 0.5288748, 0.5260245, 0.5290533, 0.5285035, 
    0.5294138, 0.5302288, 0.5312536, 0.5331438, 0.5327061, 0.5342859, 
    0.5181032, 0.5190767, 0.5189909, 0.5200092, 0.5207621, 0.522393, 
    0.5250068, 0.5240242, 0.5258277, 0.5261897, 0.5234494, 0.5251324, 
    0.5197279, 0.520602, 0.5200815, 0.5181801, 0.5242509, 0.5211372, 
    0.5268838, 0.5251991, 0.5301126, 0.5276704, 0.5324653, 0.5345126, 
    0.5364373, 0.5386853, 0.5196077, 0.5189464, 0.5201302, 0.5217674, 
    0.5232852, 0.5253019, 0.5255081, 0.5258858, 0.5268635, 0.5276854, 
    0.5260053, 0.5278914, 0.520805, 0.5245209, 0.5186965, 0.5204519, 
    0.5216709, 0.521136, 0.5239118, 0.5245656, 0.5272209, 0.5258486, 
    0.5340076, 0.5304011, 0.5403951, 0.5376064, 0.5187154, 0.5196053, 
    0.5227007, 0.5212284, 0.5254364, 0.5264713, 0.527312, 0.5283867, 
    0.5285026, 0.5291391, 0.528096, 0.5290979, 0.5253062, 0.5270013, 
    0.5223469, 0.5234806, 0.5229591, 0.522387, 0.5241522, 0.5260318, 
    0.5260717, 0.5266741, 0.5283715, 0.5254534, 0.5344732, 0.5289071, 
    0.5205755, 0.5222886, 0.5225329, 0.5218695, 0.5263675, 0.5247387, 
    0.5291235, 0.5279391, 0.5298794, 0.5289155, 0.5287736, 0.5275349, 
    0.5267635, 0.5248134, 0.5232256, 0.5219657, 0.5222587, 0.5236425, 
    0.5261467, 0.5285132, 0.527995, 0.529732, 0.5251315, 0.5270617, 
    0.5263159, 0.52826, 0.5239981, 0.5276286, 0.5230694, 0.5234694, 
    0.5247063, 0.5271928, 0.5277421, 0.5283291, 0.5279669, 0.5262101, 
    0.5259221, 0.5246762, 0.5243322, 0.5233823, 0.5225957, 0.5233145, 
    0.5240691, 0.5262108, 0.5281394, 0.5302404, 0.5307542, 0.5332069, 
    0.5312108, 0.5345042, 0.531705, 0.5365483, 0.5278384, 0.5316222, 
    0.5247625, 0.5255023, 0.5268402, 0.5299056, 0.5282509, 0.5301858, 
    0.5259108, 0.5236903, 0.5231152, 0.5220424, 0.5231398, 0.5230505, 
    0.5241002, 0.5237629, 0.5262818, 0.5249291, 0.5287701, 0.5301704, 
    0.5341204, 0.536539, 0.5389979, 0.5400829, 0.540413, 0.540551,
  0.5071225, 0.5095131, 0.5090484, 0.5109763, 0.5099068, 0.5111692, 
    0.5076072, 0.5096081, 0.5083308, 0.5073376, 0.5147167, 0.5110623, 
    0.5185099, 0.5161807, 0.5220301, 0.5181476, 0.5228127, 0.5219179, 
    0.5246101, 0.5238389, 0.5272818, 0.524966, 0.5290655, 0.5267287, 
    0.5270944, 0.5248896, 0.5117975, 0.5142619, 0.5116516, 0.5120031, 
    0.5118453, 0.509929, 0.5089633, 0.5069396, 0.507307, 0.5087932, 
    0.5121611, 0.5110178, 0.5138983, 0.5138332, 0.5170391, 0.5155938, 
    0.5209799, 0.5194494, 0.5238711, 0.5227594, 0.5238189, 0.5234976, 
    0.5238231, 0.5221925, 0.5228912, 0.5214562, 0.5158646, 0.5175084, 
    0.5126048, 0.5096552, 0.507695, 0.5063038, 0.5065005, 0.5068755, 
    0.5088019, 0.5106125, 0.5119921, 0.5129148, 0.5138239, 0.5165756, 
    0.5180311, 0.5212895, 0.5207013, 0.5216975, 0.5226488, 0.5242458, 
    0.5239829, 0.5246865, 0.5216711, 0.5236754, 0.5203664, 0.5212716, 
    0.5140719, 0.5113262, 0.5101597, 0.5091377, 0.5066518, 0.5083687, 
    0.5076919, 0.5093017, 0.5103245, 0.5098186, 0.51294, 0.5117267, 
    0.5181174, 0.5153653, 0.5225378, 0.520822, 0.522949, 0.5218637, 
    0.5237232, 0.5220497, 0.5249483, 0.5255795, 0.5251482, 0.5268044, 
    0.5219569, 0.523819, 0.5098045, 0.509887, 0.5102713, 0.5085818, 
    0.5084784, 0.5069296, 0.5083077, 0.5088945, 0.5103837, 0.5112646, 
    0.5121019, 0.5139424, 0.5159975, 0.5188702, 0.5209333, 0.5223159, 
    0.521468, 0.5222166, 0.5213798, 0.5209876, 0.525343, 0.5228978, 
    0.5265662, 0.5263632, 0.5247033, 0.5263861, 0.5099449, 0.5094701, 
    0.5078216, 0.5091117, 0.5067609, 0.508077, 0.5088336, 0.5117522, 
    0.5123932, 0.5129877, 0.5141615, 0.5156678, 0.5183095, 0.5206072, 
    0.5227041, 0.5225504, 0.5226045, 0.523073, 0.5219127, 0.5232634, 
    0.5234901, 0.5228974, 0.526336, 0.5253538, 0.5263589, 0.5257193, 
    0.5096244, 0.5104233, 0.5099916, 0.5108034, 0.5102316, 0.5127741, 
    0.5135363, 0.5171013, 0.5156382, 0.5179664, 0.5158746, 0.5162454, 
    0.5180427, 0.5159876, 0.5204808, 0.5174352, 0.5230911, 0.5200512, 
    0.5232816, 0.522695, 0.5236661, 0.524536, 0.5256299, 0.5276482, 
    0.5271808, 0.5288682, 0.5116141, 0.5126501, 0.5125587, 0.5136427, 
    0.5144442, 0.5161812, 0.5189663, 0.5179191, 0.5198414, 0.5202273, 
    0.5173066, 0.5191002, 0.5133432, 0.5142738, 0.5137196, 0.5116959, 
    0.5181606, 0.5148436, 0.5209674, 0.5191713, 0.524412, 0.5218063, 
    0.5269235, 0.5291105, 0.5311673, 0.5335712, 0.5132152, 0.5125114, 
    0.5137715, 0.5155149, 0.5171317, 0.5192809, 0.5195007, 0.5199032, 
    0.5209458, 0.5218223, 0.5200307, 0.522042, 0.5144899, 0.5184484, 
    0.5122454, 0.514114, 0.5154121, 0.5148425, 0.5177993, 0.5184961, 
    0.521327, 0.5198636, 0.528571, 0.5247199, 0.5354004, 0.5324174, 
    0.5122655, 0.5132127, 0.5165089, 0.5149407, 0.5194243, 0.5205275, 
    0.5214242, 0.5225704, 0.5226941, 0.5233731, 0.5222604, 0.5233291, 
    0.5192854, 0.5210927, 0.5161321, 0.5173398, 0.5167842, 0.5161747, 
    0.5180555, 0.520059, 0.5201015, 0.5207438, 0.5225541, 0.5194424, 
    0.5290684, 0.5231255, 0.5142456, 0.51607, 0.5163302, 0.5156236, 
    0.5204169, 0.5186805, 0.5233565, 0.522093, 0.5241631, 0.5231345, 
    0.5229832, 0.5216618, 0.5208392, 0.5187602, 0.5170682, 0.5157261, 
    0.5160382, 0.5175124, 0.5201814, 0.5227054, 0.5221526, 0.5240058, 
    0.5190992, 0.5211571, 0.520362, 0.5224352, 0.5178913, 0.5217617, 
    0.5169017, 0.5173279, 0.5186461, 0.5212969, 0.5218829, 0.5225089, 
    0.5221226, 0.5202491, 0.519942, 0.5186139, 0.5182474, 0.5172351, 
    0.5163971, 0.5171629, 0.517967, 0.5202498, 0.5223066, 0.5245484, 
    0.5250968, 0.5277156, 0.5255842, 0.5291015, 0.5261118, 0.5312861, 
    0.5219855, 0.5260233, 0.5187059, 0.5194945, 0.5209209, 0.524191, 
    0.5224255, 0.5244901, 0.51993, 0.5175633, 0.5169506, 0.5158077, 
    0.5169767, 0.5168816, 0.5180001, 0.5176407, 0.5203256, 0.5188835, 
    0.5229794, 0.5244737, 0.5286915, 0.5312761, 0.5339056, 0.5350664, 
    0.5354196, 0.5355672,
  0.5311408, 0.5336102, 0.5331299, 0.5351226, 0.534017, 0.5353221, 0.5316412, 
    0.5337083, 0.5323886, 0.531363, 0.5389929, 0.5352115, 0.5429235, 
    0.5405092, 0.5465765, 0.5425478, 0.5473893, 0.5464599, 0.549257, 
    0.5484555, 0.5520359, 0.549627, 0.5538929, 0.5514604, 0.5518409, 
    0.5495476, 0.5359719, 0.5385219, 0.535821, 0.5361845, 0.5360213, 0.53404, 
    0.533042, 0.530952, 0.5313313, 0.5328663, 0.5363479, 0.5351655, 
    0.5381456, 0.5380782, 0.5413987, 0.5399013, 0.5454862, 0.5438979, 
    0.5484889, 0.5473339, 0.5484347, 0.5481008, 0.5484391, 0.5467452, 
    0.5474708, 0.5459806, 0.5401817, 0.5418851, 0.536807, 0.5337571, 
    0.5317319, 0.5302957, 0.5304987, 0.5308858, 0.5328753, 0.5347465, 
    0.5361732, 0.5371278, 0.5380686, 0.5409184, 0.542427, 0.5458075, 
    0.545197, 0.5462311, 0.547219, 0.5488784, 0.5486052, 0.5493365, 
    0.5462037, 0.5482855, 0.5448493, 0.5457889, 0.5383253, 0.5354845, 
    0.5342784, 0.5332223, 0.5306548, 0.5324277, 0.5317287, 0.5333917, 
    0.5344488, 0.5339259, 0.5371539, 0.5358987, 0.5425165, 0.5396646, 
    0.5471038, 0.5453222, 0.5475308, 0.5464036, 0.5483353, 0.5465968, 
    0.5496086, 0.5502649, 0.5498164, 0.5515391, 0.5465004, 0.5484348, 
    0.5339113, 0.5339966, 0.5343938, 0.532648, 0.5325411, 0.5309416, 
    0.5323647, 0.532971, 0.53451, 0.5354208, 0.5362867, 0.5381913, 0.5403195, 
    0.5432972, 0.5454377, 0.5468733, 0.5459929, 0.5467702, 0.5459013, 
    0.5454941, 0.5500191, 0.5474777, 0.5512913, 0.5510802, 0.549354, 
    0.5511039, 0.5340564, 0.5335657, 0.5318627, 0.5331954, 0.5307675, 
    0.5321264, 0.5329081, 0.5359251, 0.536588, 0.5372031, 0.5384181, 
    0.5399778, 0.5427157, 0.5450993, 0.5472764, 0.5471168, 0.547173, 
    0.5476596, 0.5464545, 0.5478575, 0.5480931, 0.5474772, 0.5510519, 
    0.5500303, 0.5510756, 0.5504104, 0.5337252, 0.5345509, 0.5341047, 
    0.5349439, 0.5343527, 0.5369822, 0.5377709, 0.5414632, 0.5399472, 
    0.5423599, 0.5401922, 0.5405762, 0.542439, 0.5403092, 0.544968, 
    0.5418092, 0.5476785, 0.5445223, 0.5478764, 0.547267, 0.5482759, 0.54918, 
    0.5503173, 0.5524172, 0.5519308, 0.5536874, 0.5357822, 0.5368538, 
    0.5367593, 0.537881, 0.5387108, 0.5405097, 0.5433968, 0.5423108, 
    0.5443046, 0.544705, 0.541676, 0.5435357, 0.5375711, 0.5385343, 
    0.5379606, 0.5358668, 0.5425613, 0.5391243, 0.5454732, 0.5436094, 
    0.5490511, 0.546344, 0.5516631, 0.5539397, 0.5560828, 0.5585898, 
    0.5374387, 0.5367104, 0.5380144, 0.5398195, 0.5414947, 0.5437231, 
    0.5439511, 0.5443688, 0.5454507, 0.5463607, 0.544501, 0.5465888, 
    0.5387581, 0.5428597, 0.5364352, 0.5383689, 0.539713, 0.5391232, 
    0.5421867, 0.5429091, 0.5458464, 0.5443276, 0.5533779, 0.5493712, 
    0.5604993, 0.5573862, 0.536456, 0.5374361, 0.5408493, 0.5392249, 
    0.5438718, 0.5450166, 0.5459473, 0.5471376, 0.547266, 0.5479715, 
    0.5468156, 0.5479257, 0.5437279, 0.5456032, 0.5404589, 0.5417104, 
    0.5411345, 0.5405031, 0.5424523, 0.5445303, 0.5445745, 0.5452411, 
    0.5471207, 0.5438907, 0.5538958, 0.5477143, 0.5385051, 0.5403945, 
    0.5406641, 0.5399321, 0.5449018, 0.5431004, 0.5479542, 0.5466418, 
    0.5487924, 0.5477236, 0.5475664, 0.5461941, 0.54534, 0.543183, 0.5414289, 
    0.5400383, 0.5403615, 0.5418893, 0.5446574, 0.5472778, 0.5467036, 
    0.5486289, 0.5435347, 0.5456702, 0.5448447, 0.5469972, 0.542282, 
    0.5462978, 0.5412564, 0.541698, 0.5430647, 0.5458152, 0.5464236, 
    0.5470738, 0.5466725, 0.5447277, 0.544409, 0.5430314, 0.5426512, 
    0.5416019, 0.5407335, 0.541527, 0.5423605, 0.5447284, 0.5468636, 
    0.5491928, 0.549763, 0.5524874, 0.5502698, 0.5539303, 0.5508186, 
    0.5562065, 0.5465302, 0.5507265, 0.5431268, 0.5439447, 0.5454249, 
    0.5488214, 0.5469871, 0.5491322, 0.5443965, 0.5419421, 0.541307, 
    0.5401229, 0.541334, 0.5412355, 0.5423949, 0.5420222, 0.544807, 
    0.5433109, 0.5475625, 0.5491152, 0.5535034, 0.5561962, 0.5589388, 
    0.5601504, 0.5605193, 0.5606735,
  0.5352592, 0.5381025, 0.5375492, 0.5398464, 0.5385714, 0.5400766, 0.535835, 
    0.5382156, 0.5366953, 0.5355148, 0.5443175, 0.539949, 0.5488714, 
    0.5460728, 0.5531155, 0.5484356, 0.5540615, 0.5529799, 0.5562374, 
    0.5553032, 0.5594807, 0.5566688, 0.5616519, 0.5588083, 0.5592528, 
    0.5565763, 0.5408266, 0.5437729, 0.5406523, 0.5410719, 0.5408835, 
    0.5385979, 0.5374479, 0.535042, 0.5354784, 0.5372455, 0.5412607, 
    0.539896, 0.5433377, 0.5432599, 0.5471033, 0.5453688, 0.5518475, 
    0.5500024, 0.5553422, 0.553997, 0.555279, 0.5548901, 0.5552841, 
    0.5533118, 0.5541564, 0.5524224, 0.5456935, 0.5476671, 0.5417908, 
    0.5382718, 0.5359394, 0.5342872, 0.5345206, 0.5349658, 0.5372558, 
    0.5394126, 0.5410588, 0.5421613, 0.5432487, 0.5465468, 0.5482955, 
    0.5522211, 0.5515114, 0.5527138, 0.5538632, 0.555796, 0.5554776, 
    0.5563301, 0.5526819, 0.5551053, 0.5511074, 0.5521995, 0.5435454, 
    0.540264, 0.5388727, 0.5376555, 0.5347002, 0.5367404, 0.5359357, 
    0.5378507, 0.5390692, 0.5384664, 0.5421915, 0.540742, 0.5483992, 
    0.5450948, 0.5537291, 0.551657, 0.5542263, 0.5529145, 0.5551631, 
    0.5531392, 0.5566474, 0.5574129, 0.5568898, 0.5589003, 0.5530271, 
    0.5552791, 0.5384495, 0.5385479, 0.5390058, 0.536994, 0.536871, 
    0.5350301, 0.5366679, 0.537366, 0.5391398, 0.5401905, 0.5411899, 
    0.5433905, 0.5458531, 0.549305, 0.5517913, 0.5534609, 0.5524367, 
    0.5533409, 0.5523302, 0.5518568, 0.5571261, 0.5541644, 0.5586109, 
    0.5583644, 0.5563504, 0.5583922, 0.5386168, 0.5380512, 0.5360899, 
    0.5376245, 0.5348297, 0.5363935, 0.5372936, 0.5407724, 0.5415379, 
    0.5422484, 0.5436527, 0.5454575, 0.5486304, 0.5513979, 0.5539301, 
    0.5537444, 0.5538098, 0.5543762, 0.5529737, 0.5546067, 0.554881, 
    0.5541639, 0.5583314, 0.5571392, 0.5583591, 0.5575827, 0.5382351, 
    0.539187, 0.5386725, 0.5396402, 0.5389585, 0.5419931, 0.5429045, 
    0.547178, 0.545422, 0.5482177, 0.5457056, 0.5461504, 0.5483094, 
    0.5458412, 0.5512454, 0.5475791, 0.5543982, 0.5507275, 0.5546287, 
    0.5539191, 0.5550941, 0.5561476, 0.5574741, 0.5599262, 0.5593578, 
    0.5614114, 0.5406075, 0.5418449, 0.5417357, 0.5430318, 0.5439913, 
    0.5460733, 0.5494207, 0.5481607, 0.5504746, 0.5509398, 0.5474247, 
    0.5495818, 0.5426736, 0.5437872, 0.5431239, 0.5407051, 0.5484512, 
    0.5444697, 0.5518324, 0.5496675, 0.5559973, 0.5528452, 0.5590451, 
    0.5617067, 0.5642166, 0.5671582, 0.5425206, 0.5416791, 0.5431859, 
    0.5452742, 0.5472145, 0.5497994, 0.5500641, 0.5505492, 0.5518063, 
    0.5528646, 0.5507028, 0.5531299, 0.544046, 0.5487974, 0.5413614, 
    0.5435959, 0.5451509, 0.5444683, 0.5480168, 0.5488548, 0.5522664, 
    0.5505014, 0.5610493, 0.5563705, 0.5694026, 0.5657451, 0.5413854, 
    0.5425175, 0.5464667, 0.5445861, 0.5499721, 0.5513018, 0.5523837, 
    0.5537685, 0.553918, 0.5547394, 0.5533937, 0.5546861, 0.5498049, 
    0.5519837, 0.5460144, 0.5474645, 0.5467972, 0.5460657, 0.5483248, 
    0.5507368, 0.5507881, 0.5515627, 0.5537488, 0.5499939, 0.5616553, 
    0.5544398, 0.5437534, 0.54594, 0.5462523, 0.5454046, 0.5511684, 
    0.5490767, 0.5547193, 0.5531915, 0.5556958, 0.5544507, 0.5542676, 
    0.5526707, 0.5516776, 0.5491726, 0.5471383, 0.5455275, 0.5459018, 
    0.5476719, 0.5508845, 0.5539317, 0.5532635, 0.5555053, 0.5495807, 
    0.5520614, 0.5511021, 0.5536051, 0.5481274, 0.5527913, 0.5469384, 
    0.5474502, 0.5490352, 0.5522301, 0.5529376, 0.5536942, 0.5532272, 
    0.5509661, 0.5505959, 0.5489966, 0.5485556, 0.5473388, 0.5463325, 
    0.5472519, 0.5482184, 0.5509669, 0.5534497, 0.5561626, 0.5568274, 
    0.5600082, 0.5574186, 0.5616957, 0.558059, 0.5643616, 0.5530617, 
    0.5579516, 0.5491073, 0.5500568, 0.5517763, 0.5557296, 0.5535933, 
    0.556092, 0.5505814, 0.5477332, 0.546997, 0.5456254, 0.5470284, 
    0.5469142, 0.5482582, 0.5478261, 0.5510583, 0.5493209, 0.5542631, 
    0.5560721, 0.5611962, 0.5643494, 0.5675681, 0.5689924, 0.5694262, 
    0.5696076,
  0.5840976, 0.5875086, 0.5868437, 0.5896073, 0.5880724, 0.5898846, 
    0.5847872, 0.5876446, 0.5858188, 0.5844036, 0.5950114, 0.5897309, 
    0.6005509, 0.5971422, 0.6057471, 0.6000192, 0.6069097, 0.6055806, 
    0.6095905, 0.6084385, 0.613603, 0.610123, 0.6163005, 0.6127695, 
    0.6133204, 0.6100087, 0.5907891, 0.5943512, 0.5905789, 0.5910851, 
    0.5908578, 0.5881042, 0.5867221, 0.5838375, 0.58436, 0.586479, 0.5913129, 
    0.589667, 0.5938241, 0.5937299, 0.5983957, 0.596287, 0.6041912, 
    0.6019324, 0.6084865, 0.6068304, 0.6084087, 0.6079295, 0.6084149, 
    0.6059882, 0.6070265, 0.6048962, 0.5966813, 0.5990824, 0.5919532, 
    0.5877121, 0.5849124, 0.5829344, 0.5832136, 0.5837463, 0.5864915, 
    0.5890847, 0.5910693, 0.5924011, 0.5937164, 0.5977185, 0.5998483, 
    0.6046493, 0.6037793, 0.6052538, 0.6066659, 0.609046, 0.6086534, 
    0.6097049, 0.6052146, 0.6081945, 0.6032844, 0.6046228, 0.5940757, 
    0.5901105, 0.5884349, 0.5869715, 0.5834284, 0.5858728, 0.5849079, 
    0.587206, 0.5886714, 0.5879461, 0.5924375, 0.590687, 0.5999748, 
    0.5959544, 0.606501, 0.6039577, 0.6071125, 0.6055002, 0.6082659, 
    0.6057761, 0.6100966, 0.6110424, 0.6103959, 0.6128834, 0.6056384, 
    0.6084088, 0.5879259, 0.588044, 0.5885951, 0.5861772, 0.5860295, 
    0.5838232, 0.5857859, 0.5866238, 0.5887564, 0.5900219, 0.5912276, 
    0.593888, 0.5968752, 0.6010803, 0.6041222, 0.6061714, 0.6049138, 
    0.6060239, 0.6047831, 0.6042026, 0.6106879, 0.6070363, 0.6125249, 
    0.6122196, 0.6097299, 0.612254, 0.5881271, 0.587447, 0.5850927, 
    0.5869343, 0.5835835, 0.5854568, 0.5865368, 0.5907238, 0.5916477, 
    0.5925063, 0.5942057, 0.5963947, 0.6002568, 0.6036403, 0.6067482, 
    0.6065198, 0.6066002, 0.6072969, 0.6055729, 0.6075805, 0.6079184, 
    0.6070357, 0.6121787, 0.6107041, 0.6122131, 0.6112524, 0.5876679, 
    0.5888132, 0.5881941, 0.5893589, 0.5885381, 0.5921977, 0.5932998, 
    0.5984868, 0.5963516, 0.5997534, 0.596696, 0.5972366, 0.5998653, 
    0.5968608, 0.6034534, 0.5989752, 0.6073241, 0.6028193, 0.6076077, 
    0.6067347, 0.6081808, 0.6094796, 0.6111181, 0.6141557, 0.6134506, 
    0.6160014, 0.5905248, 0.5920186, 0.5918867, 0.5934538, 0.5946159, 
    0.5971429, 0.6012216, 0.5996841, 0.60251, 0.6030792, 0.5987871, 
    0.6014184, 0.5930204, 0.5943686, 0.5935653, 0.5906426, 0.6000383, 
    0.5951958, 0.6041727, 0.601523, 0.6092943, 0.6054151, 0.613063, 
    0.6163687, 0.619499, 0.623184, 0.5928354, 0.5918184, 0.5936404, 
    0.5961721, 0.5985312, 0.6016843, 0.6020079, 0.6026012, 0.6041408, 
    0.6054389, 0.6027891, 0.6057648, 0.5946822, 0.6004606, 0.5914346, 
    0.5941368, 0.5960224, 0.5951942, 0.5995085, 0.6005306, 0.6047048, 
    0.6025427, 0.615551, 0.6097547, 0.6260078, 0.6214116, 0.5914636, 
    0.5928317, 0.5976212, 0.595337, 0.6018954, 0.6035225, 0.6048487, 
    0.6065495, 0.6067333, 0.607744, 0.6060889, 0.6076784, 0.6016911, 
    0.6043581, 0.5970713, 0.5988357, 0.5980232, 0.5971336, 0.5998841, 
    0.6028308, 0.6028935, 0.6038421, 0.6065252, 0.6019221, 0.6163048, 
    0.6073753, 0.5943276, 0.5969808, 0.5973604, 0.5963304, 0.6033591, 
    0.6008015, 0.6077192, 0.6058404, 0.6089224, 0.6073886, 0.6071634, 
    0.6052009, 0.603983, 0.6009186, 0.5984383, 0.5964796, 0.5969344, 
    0.5990883, 0.6030115, 0.6067501, 0.6059289, 0.6086875, 0.6014171, 
    0.6044534, 0.6032779, 0.6063486, 0.5996433, 0.6053489, 0.598195, 
    0.5988182, 0.6007509, 0.6046603, 0.6055287, 0.6064581, 0.6058843, 
    0.6031114, 0.6026583, 0.6007037, 0.6001655, 0.5986825, 0.5974579, 
    0.5985767, 0.5997543, 0.6031124, 0.6061576, 0.6094982, 0.6103189, 
    0.6142576, 0.6110495, 0.6163551, 0.6118417, 0.6196803, 0.6056809, 
    0.6117087, 0.6008388, 0.6019989, 0.604104, 0.6089641, 0.6063341, 
    0.609411, 0.6026406, 0.5991629, 0.5982664, 0.5965986, 0.5983046, 
    0.5981656, 0.5998029, 0.5992761, 0.6032243, 0.6010998, 0.6071578, 
    0.6093865, 0.6157336, 0.6196651, 0.623699, 0.6254908, 0.6260375, 0.6262662,
  0.6622251, 0.667787, 0.6666976, 0.6712429, 0.6687129, 0.6717016, 0.6633443, 
    0.6680101, 0.6650231, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987642, 0.6887959, 0.7008165, 0.6984711, 0.7055877, 
    0.7035307, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626507, 0.6661011, 0.6740712, 
    0.6713416, 0.6782681, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034775, 0.7026251, 0.7034886, 
    0.6991889, 0.7010233, 0.6972684, 0.683092, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616562, 0.6661214, 
    0.6703799, 0.6736662, 0.6758848, 0.6780871, 0.6848564, 0.688502, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978275, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.669309, 0.6669068, 0.6611419, 0.6651114, 0.6635405, 
    0.6672908, 0.6696985, 0.6685052, 0.6759457, 0.6730312, 0.6887196, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115249, 0.6985729, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.665608, 0.665367, 
    0.6617807, 0.6649695, 0.6663378, 0.6698384, 0.6719288, 0.6739292, 
    0.6783753, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972994, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108743, 
    0.710321, 0.7058374, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668458, 0.6613927, 0.6644333, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826057, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002691, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075859, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.6694789, 0.6755454, 0.6773884, 
    0.6861679, 0.6825325, 0.6883391, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870038, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.713842, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750265, 0.6776467, 0.6795995, 
    0.6838763, 0.6908692, 0.6882198, 0.6931019, 0.6940922, 0.6866817, 
    0.6912096, 0.6769205, 0.6791831, 0.6778337, 0.6729575, 0.6888287, 
    0.6805774, 0.6960008, 0.6913906, 0.7050577, 0.69818, 0.711851, 0.7179045, 
    0.7237219, 0.7306815, 0.6766108, 0.6749127, 0.6779597, 0.6822283, 
    0.6862438, 0.6916698, 0.6922304, 0.6932604, 0.6959449, 0.6982217, 
    0.6935872, 0.6987953, 0.6797112, 0.6895558, 0.6742736, 0.6787933, 
    0.6819748, 0.6805746, 0.6879184, 0.6896765, 0.6969327, 0.6931587, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846905, 0.6808156, 0.6920354, 0.6948648, 0.6971852, 0.7001796, 
    0.7005044, 0.7022954, 0.6993665, 0.702179, 0.6916814, 0.6963252, 
    0.6837546, 0.6867649, 0.685376, 0.6838604, 0.6885635, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016412, 
    0.6791143, 0.6836007, 0.6842464, 0.6824967, 0.6945799, 0.6901437, 
    0.7022516, 0.6989285, 0.7043934, 0.7016648, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.6860851, 0.6827497, 0.6835218, 0.6871974, 
    0.6939742, 0.7005342, 0.6990844, 0.7039744, 0.6912072, 0.6964923, 
    0.6944383, 0.6998248, 0.6881498, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863217, 
    0.6883404, 0.6941499, 0.6994876, 0.7054225, 0.7068936, 0.7140281, 
    0.7082077, 0.7178792, 0.7096372, 0.7240614, 0.6986477, 0.709397, 
    0.6902081, 0.6922148, 0.6958807, 0.7044679, 0.6997992, 0.7052665, 
    0.6933289, 0.6873254, 0.6857913, 0.6829515, 0.6858565, 0.6856191, 
    0.6884239, 0.6875196, 0.6943448, 0.6906587, 0.7012558, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.462176e-11, 3.477718e-11, 3.474688e-11, 3.487233e-11, 3.48027e-11, 
    3.488479e-11, 3.465309e-11, 3.478307e-11, 3.470003e-11, 3.463545e-11, 
    3.511576e-11, 3.487763e-11, 3.536388e-11, 3.521152e-11, 3.559451e-11, 
    3.534002e-11, 3.564586e-11, 3.558712e-11, 3.576395e-11, 3.571321e-11, 
    3.593947e-11, 3.578725e-11, 3.605698e-11, 3.590307e-11, 3.592706e-11, 
    3.578203e-11, 3.492585e-11, 3.508635e-11, 3.491625e-11, 3.493914e-11, 
    3.492884e-11, 3.480395e-11, 3.474104e-11, 3.460958e-11, 3.463339e-11, 
    3.472994e-11, 3.494915e-11, 3.487466e-11, 3.506242e-11, 3.505819e-11, 
    3.52675e-11, 3.517305e-11, 3.552555e-11, 3.54252e-11, 3.571528e-11, 
    3.564219e-11, 3.571176e-11, 3.56906e-11, 3.571192e-11, 3.560485e-11, 
    3.565063e-11, 3.555647e-11, 3.519117e-11, 3.529858e-11, 3.49783e-11, 
    3.4786e-11, 3.465861e-11, 3.45683e-11, 3.458098e-11, 3.460531e-11, 
    3.473043e-11, 3.484824e-11, 3.49381e-11, 3.49982e-11, 3.505746e-11, 
    3.523702e-11, 3.533225e-11, 3.554572e-11, 3.55072e-11, 3.557242e-11, 
    3.563488e-11, 3.573972e-11, 3.572244e-11, 3.57686e-11, 3.557054e-11, 
    3.570209e-11, 3.548492e-11, 3.554426e-11, 3.507375e-11, 3.489492e-11, 
    3.48188e-11, 3.475235e-11, 3.459076e-11, 3.470229e-11, 3.465826e-11, 
    3.47629e-11, 3.482944e-11, 3.479647e-11, 3.499981e-11, 3.492064e-11, 
    3.533784e-11, 3.515794e-11, 3.562765e-11, 3.551502e-11, 3.565454e-11, 
    3.558332e-11, 3.570529e-11, 3.559545e-11, 3.578575e-11, 3.582722e-11, 
    3.579879e-11, 3.590779e-11, 3.558911e-11, 3.571135e-11, 3.479576e-11, 
    3.480113e-11, 3.482611e-11, 3.471608e-11, 3.470935e-11, 3.460869e-11, 
    3.469817e-11, 3.473631e-11, 3.483322e-11, 3.48905e-11, 3.4945e-11, 
    3.506504e-11, 3.519917e-11, 3.538704e-11, 3.552227e-11, 3.561294e-11, 
    3.555729e-11, 3.560634e-11, 3.555142e-11, 3.552564e-11, 3.581156e-11, 
    3.565089e-11, 3.5892e-11, 3.587866e-11, 3.576939e-11, 3.588005e-11, 
    3.480483e-11, 3.477389e-11, 3.466665e-11, 3.47505e-11, 3.459767e-11, 
    3.468314e-11, 3.473224e-11, 3.492219e-11, 3.496398e-11, 3.500273e-11, 
    3.507928e-11, 3.517759e-11, 3.53503e-11, 3.550078e-11, 3.563837e-11, 
    3.562823e-11, 3.563176e-11, 3.566244e-11, 3.558627e-11, 3.567487e-11, 
    3.568969e-11, 3.56508e-11, 3.587676e-11, 3.581215e-11, 3.587822e-11, 
    3.583609e-11, 3.478389e-11, 3.483581e-11, 3.480767e-11, 3.48605e-11, 
    3.482318e-11, 3.498879e-11, 3.503843e-11, 3.527126e-11, 3.517563e-11, 
    3.532786e-11, 3.519103e-11, 3.521524e-11, 3.53326e-11, 3.519833e-11, 
    3.549231e-11, 3.529276e-11, 3.566359e-11, 3.546395e-11, 3.567603e-11, 
    3.563746e-11, 3.570119e-11, 3.575833e-11, 3.583019e-11, 3.596299e-11, 
    3.593215e-11, 3.604333e-11, 3.491333e-11, 3.498075e-11, 3.497483e-11, 
    3.504546e-11, 3.509771e-11, 3.521121e-11, 3.539335e-11, 3.532476e-11, 
    3.54506e-11, 3.547588e-11, 3.528457e-11, 3.540191e-11, 3.502557e-11, 
    3.508618e-11, 3.505007e-11, 3.491804e-11, 3.534017e-11, 3.512324e-11, 
    3.552404e-11, 3.540627e-11, 3.575006e-11, 3.557891e-11, 3.591519e-11, 
    3.605915e-11, 3.619492e-11, 3.635353e-11, 3.50176e-11, 3.497166e-11, 
    3.505381e-11, 3.516755e-11, 3.527322e-11, 3.54139e-11, 3.542828e-11, 
    3.545458e-11, 3.552289e-11, 3.558039e-11, 3.546278e-11, 3.55947e-11, 
    3.510013e-11, 3.535902e-11, 3.495378e-11, 3.50756e-11, 3.516033e-11, 
    3.512316e-11, 3.531644e-11, 3.536198e-11, 3.554737e-11, 3.545151e-11, 
    3.602345e-11, 3.577005e-11, 3.647454e-11, 3.627724e-11, 3.495559e-11, 
    3.50173e-11, 3.523244e-11, 3.513002e-11, 3.542321e-11, 3.54955e-11, 
    3.555424e-11, 3.562942e-11, 3.563749e-11, 3.568206e-11, 3.560895e-11, 
    3.567912e-11, 3.541379e-11, 3.553226e-11, 3.520745e-11, 3.528633e-11, 
    3.525001e-11, 3.521011e-11, 3.533306e-11, 3.546419e-11, 3.546701e-11, 
    3.550901e-11, 3.562748e-11, 3.542369e-11, 3.605592e-11, 3.56649e-11, 
    3.508465e-11, 3.520365e-11, 3.522069e-11, 3.517455e-11, 3.548814e-11, 
    3.537439e-11, 3.568099e-11, 3.559799e-11, 3.573388e-11, 3.566631e-11, 
    3.565628e-11, 3.556958e-11, 3.551552e-11, 3.537928e-11, 3.526848e-11, 
    3.51808e-11, 3.52011e-11, 3.529746e-11, 3.547212e-11, 3.563772e-11, 
    3.560137e-11, 3.572306e-11, 3.540113e-11, 3.553597e-11, 3.548373e-11, 
    3.561979e-11, 3.532277e-11, 3.557613e-11, 3.525802e-11, 3.528583e-11, 
    3.537202e-11, 3.554566e-11, 3.558412e-11, 3.562518e-11, 3.559978e-11, 
    3.547686e-11, 3.545671e-11, 3.536969e-11, 3.53456e-11, 3.527943e-11, 
    3.522454e-11, 3.52746e-11, 3.532709e-11, 3.547663e-11, 3.561147e-11, 
    3.575865e-11, 3.579473e-11, 3.59668e-11, 3.582655e-11, 3.605789e-11, 
    3.586096e-11, 3.620203e-11, 3.559082e-11, 3.585611e-11, 3.537598e-11, 
    3.542756e-11, 3.552094e-11, 3.573552e-11, 3.561962e-11, 3.575515e-11, 
    3.54559e-11, 3.530081e-11, 3.526077e-11, 3.518606e-11, 3.52624e-11, 
    3.52562e-11, 3.532932e-11, 3.530574e-11, 3.548149e-11, 3.538704e-11, 
    3.565551e-11, 3.575364e-11, 3.60312e-11, 3.620157e-11, 3.637539e-11, 
    3.64521e-11, 3.647546e-11, 3.648519e-11,
  1.775611e-11, 1.789055e-11, 1.786439e-11, 1.797303e-11, 1.791274e-11, 
    1.798391e-11, 1.778335e-11, 1.789588e-11, 1.782402e-11, 1.776822e-11, 
    1.818451e-11, 1.797788e-11, 1.840021e-11, 1.826772e-11, 1.860125e-11, 
    1.837955e-11, 1.864608e-11, 1.859487e-11, 1.874922e-11, 1.870495e-11, 
    1.890281e-11, 1.876966e-11, 1.900572e-11, 1.8871e-11, 1.889204e-11, 
    1.876527e-11, 1.801942e-11, 1.815873e-11, 1.801118e-11, 1.803101e-11, 
    1.802212e-11, 1.791398e-11, 1.785956e-11, 1.774587e-11, 1.77665e-11, 
    1.785001e-11, 1.803994e-11, 1.79754e-11, 1.813827e-11, 1.813459e-11, 
    1.831652e-11, 1.823441e-11, 1.854122e-11, 1.845384e-11, 1.87068e-11, 
    1.864306e-11, 1.87038e-11, 1.868538e-11, 1.870404e-11, 1.861059e-11, 
    1.865061e-11, 1.856846e-11, 1.824977e-11, 1.834321e-11, 1.806504e-11, 
    1.78985e-11, 1.778827e-11, 1.771019e-11, 1.772122e-11, 1.774225e-11, 
    1.78505e-11, 1.795253e-11, 1.803043e-11, 1.80826e-11, 1.813406e-11, 
    1.829009e-11, 1.837294e-11, 1.85589e-11, 1.852531e-11, 1.858224e-11, 
    1.863672e-11, 1.872829e-11, 1.871321e-11, 1.875359e-11, 1.858076e-11, 
    1.869555e-11, 1.850619e-11, 1.85579e-11, 1.814796e-11, 1.799281e-11, 
    1.792693e-11, 1.786941e-11, 1.77297e-11, 1.782614e-11, 1.77881e-11, 
    1.787867e-11, 1.793629e-11, 1.790779e-11, 1.808402e-11, 1.801543e-11, 
    1.837785e-11, 1.822141e-11, 1.863037e-11, 1.853221e-11, 1.865393e-11, 
    1.859178e-11, 1.86983e-11, 1.860243e-11, 1.876863e-11, 1.880488e-11, 
    1.878011e-11, 1.887539e-11, 1.859711e-11, 1.870379e-11, 1.790698e-11, 
    1.791163e-11, 1.79333e-11, 1.783812e-11, 1.783231e-11, 1.77453e-11, 
    1.782273e-11, 1.785573e-11, 1.793964e-11, 1.798933e-11, 1.803662e-11, 
    1.814075e-11, 1.82573e-11, 1.842077e-11, 1.853856e-11, 1.861767e-11, 
    1.856915e-11, 1.861198e-11, 1.85641e-11, 1.854168e-11, 1.879129e-11, 
    1.865097e-11, 1.886167e-11, 1.884999e-11, 1.875454e-11, 1.885131e-11, 
    1.79149e-11, 1.788815e-11, 1.77954e-11, 1.786797e-11, 1.773584e-11, 
    1.780974e-11, 1.785228e-11, 1.801684e-11, 1.805309e-11, 1.80867e-11, 
    1.815318e-11, 1.823861e-11, 1.838883e-11, 1.851991e-11, 1.86399e-11, 
    1.86311e-11, 1.86342e-11, 1.866103e-11, 1.859458e-11, 1.867194e-11, 
    1.868493e-11, 1.865097e-11, 1.884843e-11, 1.879194e-11, 1.884974e-11, 
    1.881296e-11, 1.789685e-11, 1.794187e-11, 1.791753e-11, 1.796329e-11, 
    1.793104e-11, 1.807459e-11, 1.811771e-11, 1.832002e-11, 1.823692e-11, 
    1.836927e-11, 1.825035e-11, 1.82714e-11, 1.837355e-11, 1.825678e-11, 
    1.851266e-11, 1.8339e-11, 1.866207e-11, 1.848809e-11, 1.867299e-11, 
    1.863938e-11, 1.869505e-11, 1.874494e-11, 1.880781e-11, 1.892396e-11, 
    1.889705e-11, 1.899436e-11, 1.800907e-11, 1.806759e-11, 1.806246e-11, 
    1.812379e-11, 1.816919e-11, 1.826777e-11, 1.842627e-11, 1.836661e-11, 
    1.847621e-11, 1.849823e-11, 1.833176e-11, 1.843389e-11, 1.810682e-11, 
    1.815949e-11, 1.812814e-11, 1.801367e-11, 1.838033e-11, 1.81918e-11, 
    1.854051e-11, 1.843796e-11, 1.873783e-11, 1.858846e-11, 1.888223e-11, 
    1.900828e-11, 1.912728e-11, 1.926657e-11, 1.809958e-11, 1.805978e-11, 
    1.813109e-11, 1.822989e-11, 1.832179e-11, 1.844421e-11, 1.845676e-11, 
    1.847973e-11, 1.853929e-11, 1.858941e-11, 1.848697e-11, 1.860199e-11, 
    1.817168e-11, 1.839673e-11, 1.804472e-11, 1.815043e-11, 1.822407e-11, 
    1.819177e-11, 1.83598e-11, 1.839948e-11, 1.856105e-11, 1.847747e-11, 
    1.897712e-11, 1.875546e-11, 1.937294e-11, 1.919964e-11, 1.804588e-11, 
    1.809946e-11, 1.828637e-11, 1.819735e-11, 1.84524e-11, 1.851537e-11, 
    1.856664e-11, 1.863222e-11, 1.863932e-11, 1.867823e-11, 1.861449e-11, 
    1.867571e-11, 1.844447e-11, 1.854768e-11, 1.826499e-11, 1.833363e-11, 
    1.830205e-11, 1.826741e-11, 1.837439e-11, 1.848858e-11, 1.849105e-11, 
    1.852772e-11, 1.863113e-11, 1.845344e-11, 1.900574e-11, 1.86639e-11, 
    1.815795e-11, 1.82614e-11, 1.827623e-11, 1.823611e-11, 1.850906e-11, 
    1.840998e-11, 1.867728e-11, 1.860491e-11, 1.872355e-11, 1.866456e-11, 
    1.865588e-11, 1.858023e-11, 1.853318e-11, 1.841451e-11, 1.831818e-11, 
    1.824193e-11, 1.825965e-11, 1.834344e-11, 1.849558e-11, 1.863995e-11, 
    1.860829e-11, 1.871453e-11, 1.843386e-11, 1.855134e-11, 1.850589e-11, 
    1.862449e-11, 1.836502e-11, 1.85858e-11, 1.830873e-11, 1.833297e-11, 
    1.840802e-11, 1.85593e-11, 1.859288e-11, 1.86287e-11, 1.86066e-11, 
    1.849945e-11, 1.848193e-11, 1.84062e-11, 1.838529e-11, 1.83277e-11, 
    1.828005e-11, 1.832357e-11, 1.836932e-11, 1.849951e-11, 1.861711e-11, 
    1.874565e-11, 1.877717e-11, 1.892777e-11, 1.88051e-11, 1.900764e-11, 
    1.883533e-11, 1.913401e-11, 1.859867e-11, 1.883033e-11, 1.841144e-11, 
    1.845641e-11, 1.853782e-11, 1.872509e-11, 1.862394e-11, 1.874227e-11, 
    1.848125e-11, 1.834632e-11, 1.831151e-11, 1.824656e-11, 1.831299e-11, 
    1.830759e-11, 1.837124e-11, 1.835077e-11, 1.850384e-11, 1.842156e-11, 
    1.865566e-11, 1.874134e-11, 1.898414e-11, 1.913352e-11, 1.928606e-11, 
    1.935352e-11, 1.937408e-11, 1.938267e-11,
  1.677678e-11, 1.692554e-11, 1.689658e-11, 1.701688e-11, 1.695011e-11, 
    1.702894e-11, 1.68069e-11, 1.693145e-11, 1.68519e-11, 1.679016e-11, 
    1.725135e-11, 1.702226e-11, 1.749078e-11, 1.734365e-11, 1.771427e-11, 
    1.746784e-11, 1.776415e-11, 1.770717e-11, 1.787894e-11, 1.782966e-11, 
    1.805009e-11, 1.790171e-11, 1.816483e-11, 1.801462e-11, 1.803808e-11, 
    1.789682e-11, 1.706827e-11, 1.722276e-11, 1.705914e-11, 1.708112e-11, 
    1.707126e-11, 1.695148e-11, 1.689125e-11, 1.676544e-11, 1.678826e-11, 
    1.688068e-11, 1.709102e-11, 1.70195e-11, 1.720002e-11, 1.719593e-11, 
    1.739782e-11, 1.730667e-11, 1.76475e-11, 1.755034e-11, 1.783172e-11, 
    1.776078e-11, 1.782838e-11, 1.780787e-11, 1.782865e-11, 1.772465e-11, 
    1.776918e-11, 1.767779e-11, 1.732372e-11, 1.742746e-11, 1.711883e-11, 
    1.693436e-11, 1.681235e-11, 1.672599e-11, 1.673819e-11, 1.676145e-11, 
    1.688122e-11, 1.699417e-11, 1.708046e-11, 1.713829e-11, 1.719534e-11, 
    1.73685e-11, 1.746048e-11, 1.766716e-11, 1.76298e-11, 1.769312e-11, 
    1.775373e-11, 1.785565e-11, 1.783886e-11, 1.788382e-11, 1.769146e-11, 
    1.78192e-11, 1.760853e-11, 1.766604e-11, 1.721081e-11, 1.703879e-11, 
    1.696584e-11, 1.690214e-11, 1.674757e-11, 1.685425e-11, 1.681216e-11, 
    1.691238e-11, 1.697618e-11, 1.694462e-11, 1.713987e-11, 1.706384e-11, 
    1.746594e-11, 1.729226e-11, 1.774665e-11, 1.763747e-11, 1.777287e-11, 
    1.770372e-11, 1.782226e-11, 1.771557e-11, 1.790057e-11, 1.794095e-11, 
    1.791335e-11, 1.80195e-11, 1.770966e-11, 1.782837e-11, 1.694373e-11, 
    1.694888e-11, 1.697287e-11, 1.686751e-11, 1.686108e-11, 1.676482e-11, 
    1.685047e-11, 1.688699e-11, 1.697989e-11, 1.703493e-11, 1.708733e-11, 
    1.720277e-11, 1.733209e-11, 1.751362e-11, 1.764454e-11, 1.773252e-11, 
    1.767855e-11, 1.77262e-11, 1.767294e-11, 1.7648e-11, 1.792581e-11, 
    1.776959e-11, 1.800421e-11, 1.79912e-11, 1.788488e-11, 1.799267e-11, 
    1.695249e-11, 1.692288e-11, 1.682023e-11, 1.690054e-11, 1.675435e-11, 
    1.683611e-11, 1.688319e-11, 1.706542e-11, 1.710558e-11, 1.714284e-11, 
    1.721655e-11, 1.731133e-11, 1.747812e-11, 1.762381e-11, 1.775726e-11, 
    1.774746e-11, 1.775091e-11, 1.778077e-11, 1.770684e-11, 1.779292e-11, 
    1.780738e-11, 1.776958e-11, 1.798946e-11, 1.792652e-11, 1.799092e-11, 
    1.794994e-11, 1.69325e-11, 1.698235e-11, 1.695541e-11, 1.700609e-11, 
    1.697037e-11, 1.712943e-11, 1.717724e-11, 1.740172e-11, 1.730946e-11, 
    1.745641e-11, 1.732436e-11, 1.734773e-11, 1.746119e-11, 1.733149e-11, 
    1.761575e-11, 1.74228e-11, 1.778193e-11, 1.758845e-11, 1.779408e-11, 
    1.775668e-11, 1.781863e-11, 1.787419e-11, 1.79442e-11, 1.807366e-11, 
    1.804365e-11, 1.815215e-11, 1.70568e-11, 1.712166e-11, 1.711596e-11, 
    1.718395e-11, 1.723431e-11, 1.734369e-11, 1.751972e-11, 1.745344e-11, 
    1.757521e-11, 1.759969e-11, 1.741473e-11, 1.752819e-11, 1.716514e-11, 
    1.722357e-11, 1.718878e-11, 1.70619e-11, 1.746869e-11, 1.725941e-11, 
    1.76467e-11, 1.753271e-11, 1.786626e-11, 1.770004e-11, 1.802714e-11, 
    1.81677e-11, 1.830046e-11, 1.845605e-11, 1.715712e-11, 1.7113e-11, 
    1.719205e-11, 1.730167e-11, 1.740367e-11, 1.753965e-11, 1.75536e-11, 
    1.757913e-11, 1.764534e-11, 1.770109e-11, 1.758719e-11, 1.771508e-11, 
    1.723711e-11, 1.748691e-11, 1.709631e-11, 1.721352e-11, 1.72952e-11, 
    1.725936e-11, 1.744587e-11, 1.748995e-11, 1.766955e-11, 1.757662e-11, 
    1.813295e-11, 1.788592e-11, 1.857492e-11, 1.838128e-11, 1.709759e-11, 
    1.715698e-11, 1.736434e-11, 1.726555e-11, 1.754875e-11, 1.761875e-11, 
    1.767576e-11, 1.774872e-11, 1.775661e-11, 1.779991e-11, 1.772898e-11, 
    1.779711e-11, 1.753994e-11, 1.765467e-11, 1.73406e-11, 1.741682e-11, 
    1.738174e-11, 1.734329e-11, 1.746207e-11, 1.758898e-11, 1.759171e-11, 
    1.763249e-11, 1.774756e-11, 1.75499e-11, 1.816491e-11, 1.778402e-11, 
    1.722184e-11, 1.733664e-11, 1.735309e-11, 1.730855e-11, 1.761173e-11, 
    1.750162e-11, 1.779886e-11, 1.771832e-11, 1.785037e-11, 1.77847e-11, 
    1.777505e-11, 1.769088e-11, 1.763855e-11, 1.750666e-11, 1.739965e-11, 
    1.731501e-11, 1.733468e-11, 1.742771e-11, 1.759676e-11, 1.775732e-11, 
    1.772209e-11, 1.784032e-11, 1.752815e-11, 1.765876e-11, 1.760822e-11, 
    1.774012e-11, 1.745168e-11, 1.769712e-11, 1.738916e-11, 1.741608e-11, 
    1.749944e-11, 1.766762e-11, 1.770495e-11, 1.77448e-11, 1.772021e-11, 
    1.760106e-11, 1.758158e-11, 1.749741e-11, 1.747419e-11, 1.741022e-11, 
    1.735732e-11, 1.740564e-11, 1.745645e-11, 1.760112e-11, 1.773191e-11, 
    1.787498e-11, 1.791007e-11, 1.807793e-11, 1.794121e-11, 1.816703e-11, 
    1.797493e-11, 1.830803e-11, 1.771142e-11, 1.796933e-11, 1.750324e-11, 
    1.755321e-11, 1.764373e-11, 1.78521e-11, 1.77395e-11, 1.787123e-11, 
    1.758082e-11, 1.743092e-11, 1.739224e-11, 1.732015e-11, 1.739389e-11, 
    1.738789e-11, 1.745857e-11, 1.743584e-11, 1.760593e-11, 1.751448e-11, 
    1.77748e-11, 1.787019e-11, 1.814076e-11, 1.830745e-11, 1.84778e-11, 
    1.855321e-11, 1.857619e-11, 1.85858e-11,
  1.722123e-11, 1.738505e-11, 1.735315e-11, 1.748571e-11, 1.741212e-11, 
    1.7499e-11, 1.725439e-11, 1.739157e-11, 1.730393e-11, 1.723595e-11, 
    1.774434e-11, 1.749163e-11, 1.800873e-11, 1.784619e-11, 1.825586e-11, 
    1.798339e-11, 1.831105e-11, 1.824798e-11, 1.843812e-11, 1.838356e-11, 
    1.862778e-11, 1.846334e-11, 1.8755e-11, 1.858845e-11, 1.861445e-11, 
    1.845792e-11, 1.754235e-11, 1.771278e-11, 1.753228e-11, 1.755653e-11, 
    1.754565e-11, 1.741363e-11, 1.734728e-11, 1.720874e-11, 1.723386e-11, 
    1.733563e-11, 1.756744e-11, 1.748859e-11, 1.768765e-11, 1.768314e-11, 
    1.790601e-11, 1.780536e-11, 1.818198e-11, 1.807455e-11, 1.838583e-11, 
    1.830731e-11, 1.838214e-11, 1.835943e-11, 1.838243e-11, 1.826733e-11, 
    1.83166e-11, 1.821548e-11, 1.782419e-11, 1.793876e-11, 1.75981e-11, 
    1.739479e-11, 1.726039e-11, 1.716532e-11, 1.717875e-11, 1.720435e-11, 
    1.733623e-11, 1.746067e-11, 1.755579e-11, 1.761955e-11, 1.76825e-11, 
    1.787366e-11, 1.797525e-11, 1.820373e-11, 1.81624e-11, 1.823245e-11, 
    1.82995e-11, 1.841233e-11, 1.839374e-11, 1.844353e-11, 1.823061e-11, 
    1.837198e-11, 1.813888e-11, 1.820249e-11, 1.76996e-11, 1.750984e-11, 
    1.742947e-11, 1.735928e-11, 1.718907e-11, 1.730652e-11, 1.726018e-11, 
    1.737054e-11, 1.744085e-11, 1.740606e-11, 1.76213e-11, 1.753747e-11, 
    1.798128e-11, 1.778946e-11, 1.829167e-11, 1.817088e-11, 1.832069e-11, 
    1.824417e-11, 1.837537e-11, 1.825727e-11, 1.846208e-11, 1.850682e-11, 
    1.847624e-11, 1.859385e-11, 1.825074e-11, 1.838213e-11, 1.740508e-11, 
    1.741075e-11, 1.743719e-11, 1.732114e-11, 1.731405e-11, 1.720806e-11, 
    1.730236e-11, 1.734259e-11, 1.744493e-11, 1.750559e-11, 1.756336e-11, 
    1.76907e-11, 1.783343e-11, 1.803396e-11, 1.81787e-11, 1.827604e-11, 
    1.821632e-11, 1.826904e-11, 1.821011e-11, 1.818253e-11, 1.849005e-11, 
    1.831706e-11, 1.857691e-11, 1.856248e-11, 1.844471e-11, 1.856411e-11, 
    1.741474e-11, 1.738211e-11, 1.726906e-11, 1.73575e-11, 1.719653e-11, 
    1.728654e-11, 1.73384e-11, 1.753921e-11, 1.758349e-11, 1.762458e-11, 
    1.770589e-11, 1.78105e-11, 1.799474e-11, 1.815578e-11, 1.830341e-11, 
    1.829257e-11, 1.829639e-11, 1.832944e-11, 1.824762e-11, 1.834288e-11, 
    1.835889e-11, 1.831705e-11, 1.856055e-11, 1.849083e-11, 1.856218e-11, 
    1.851676e-11, 1.739271e-11, 1.744765e-11, 1.741795e-11, 1.747381e-11, 
    1.743445e-11, 1.76098e-11, 1.766254e-11, 1.791033e-11, 1.780844e-11, 
    1.797074e-11, 1.78249e-11, 1.78507e-11, 1.797604e-11, 1.783276e-11, 
    1.814688e-11, 1.793362e-11, 1.833072e-11, 1.811671e-11, 1.834417e-11, 
    1.830277e-11, 1.837134e-11, 1.843287e-11, 1.851041e-11, 1.865389e-11, 
    1.862062e-11, 1.874092e-11, 1.752969e-11, 1.760123e-11, 1.759493e-11, 
    1.766993e-11, 1.77255e-11, 1.784623e-11, 1.80407e-11, 1.796745e-11, 
    1.810204e-11, 1.812911e-11, 1.792469e-11, 1.805007e-11, 1.764919e-11, 
    1.771366e-11, 1.767526e-11, 1.753533e-11, 1.798431e-11, 1.775321e-11, 
    1.81811e-11, 1.805506e-11, 1.842409e-11, 1.824011e-11, 1.860232e-11, 
    1.875819e-11, 1.890549e-11, 1.90783e-11, 1.764034e-11, 1.759166e-11, 
    1.767886e-11, 1.779985e-11, 1.791248e-11, 1.806273e-11, 1.807814e-11, 
    1.810637e-11, 1.817959e-11, 1.824126e-11, 1.81153e-11, 1.825673e-11, 
    1.772862e-11, 1.800444e-11, 1.757327e-11, 1.770257e-11, 1.779271e-11, 
    1.775314e-11, 1.795909e-11, 1.80078e-11, 1.820638e-11, 1.810359e-11, 
    1.871966e-11, 1.844587e-11, 1.921041e-11, 1.899524e-11, 1.757467e-11, 
    1.764017e-11, 1.786905e-11, 1.775997e-11, 1.807279e-11, 1.815019e-11, 
    1.821323e-11, 1.829397e-11, 1.83027e-11, 1.835063e-11, 1.827212e-11, 
    1.834752e-11, 1.806305e-11, 1.818991e-11, 1.784282e-11, 1.7927e-11, 
    1.788825e-11, 1.784579e-11, 1.797699e-11, 1.811727e-11, 1.812028e-11, 
    1.816538e-11, 1.829273e-11, 1.807406e-11, 1.875512e-11, 1.833307e-11, 
    1.771173e-11, 1.783847e-11, 1.785661e-11, 1.780744e-11, 1.814242e-11, 
    1.80207e-11, 1.834946e-11, 1.826033e-11, 1.840648e-11, 1.833378e-11, 
    1.83231e-11, 1.822996e-11, 1.817209e-11, 1.802627e-11, 1.790804e-11, 
    1.781457e-11, 1.783628e-11, 1.793904e-11, 1.812587e-11, 1.830349e-11, 
    1.826451e-11, 1.839535e-11, 1.805002e-11, 1.819444e-11, 1.813855e-11, 
    1.828445e-11, 1.796551e-11, 1.823691e-11, 1.789645e-11, 1.792618e-11, 
    1.801828e-11, 1.820425e-11, 1.824552e-11, 1.828963e-11, 1.826241e-11, 
    1.813063e-11, 1.810909e-11, 1.801604e-11, 1.799039e-11, 1.79197e-11, 
    1.786128e-11, 1.791465e-11, 1.797079e-11, 1.813069e-11, 1.827537e-11, 
    1.843374e-11, 1.84726e-11, 1.865865e-11, 1.850712e-11, 1.875749e-11, 
    1.854452e-11, 1.891393e-11, 1.825271e-11, 1.853828e-11, 1.802248e-11, 
    1.807771e-11, 1.817782e-11, 1.840842e-11, 1.828376e-11, 1.842959e-11, 
    1.810824e-11, 1.794259e-11, 1.789985e-11, 1.782024e-11, 1.790167e-11, 
    1.789504e-11, 1.797312e-11, 1.794801e-11, 1.813601e-11, 1.803491e-11, 
    1.832283e-11, 1.842844e-11, 1.872829e-11, 1.891326e-11, 1.910245e-11, 
    1.918626e-11, 1.921181e-11, 1.922249e-11,
  1.879543e-11, 1.897097e-11, 1.893677e-11, 1.907889e-11, 1.899998e-11, 
    1.909315e-11, 1.883094e-11, 1.897796e-11, 1.888403e-11, 1.88112e-11, 
    1.935646e-11, 1.908525e-11, 1.964051e-11, 1.946582e-11, 1.990637e-11, 
    1.961327e-11, 1.996578e-11, 1.989788e-11, 2.010264e-11, 2.004385e-11, 
    2.03071e-11, 2.012981e-11, 2.044435e-11, 2.026468e-11, 2.029272e-11, 
    2.012397e-11, 1.913965e-11, 1.932258e-11, 1.912884e-11, 1.915486e-11, 
    1.914318e-11, 1.900161e-11, 1.89305e-11, 1.878205e-11, 1.880895e-11, 
    1.8918e-11, 1.916656e-11, 1.908198e-11, 1.929556e-11, 1.929072e-11, 
    1.953009e-11, 1.942196e-11, 1.982684e-11, 1.971127e-11, 2.00463e-11, 
    1.996174e-11, 2.004233e-11, 2.001787e-11, 2.004265e-11, 1.991871e-11, 
    1.997175e-11, 1.986289e-11, 1.944218e-11, 1.956528e-11, 1.919946e-11, 
    1.898142e-11, 1.883738e-11, 1.873555e-11, 1.874993e-11, 1.877735e-11, 
    1.891864e-11, 1.905204e-11, 1.915406e-11, 1.922247e-11, 1.929003e-11, 
    1.949535e-11, 1.960452e-11, 1.985026e-11, 1.980578e-11, 1.988117e-11, 
    1.995334e-11, 2.007485e-11, 2.005482e-11, 2.010847e-11, 1.987917e-11, 
    2.003139e-11, 1.978046e-11, 1.984891e-11, 1.930843e-11, 1.910477e-11, 
    1.90186e-11, 1.894335e-11, 1.876099e-11, 1.888681e-11, 1.883715e-11, 
    1.895541e-11, 1.903078e-11, 1.899348e-11, 1.922435e-11, 1.91344e-11, 
    1.9611e-11, 1.940488e-11, 1.994491e-11, 1.98149e-11, 1.997614e-11, 
    1.989377e-11, 2.003504e-11, 1.990787e-11, 2.012845e-11, 2.017667e-11, 
    2.014371e-11, 2.027049e-11, 1.990084e-11, 2.004233e-11, 1.899244e-11, 
    1.899852e-11, 1.902686e-11, 1.890247e-11, 1.889487e-11, 1.878132e-11, 
    1.888234e-11, 1.892545e-11, 1.903516e-11, 1.910022e-11, 1.916218e-11, 
    1.929884e-11, 1.945212e-11, 1.966763e-11, 1.982331e-11, 1.992807e-11, 
    1.986379e-11, 1.992053e-11, 1.985711e-11, 1.982743e-11, 2.01586e-11, 
    1.997225e-11, 2.025223e-11, 2.023667e-11, 2.010975e-11, 2.023843e-11, 
    1.900279e-11, 1.896781e-11, 1.884667e-11, 1.894144e-11, 1.876897e-11, 
    1.88654e-11, 1.892098e-11, 1.913628e-11, 1.918377e-11, 1.922788e-11, 
    1.931514e-11, 1.942748e-11, 1.962546e-11, 1.979866e-11, 1.995754e-11, 
    1.994587e-11, 1.994998e-11, 1.998557e-11, 1.989748e-11, 2.000005e-11, 
    2.00173e-11, 1.997223e-11, 2.023459e-11, 2.015943e-11, 2.023634e-11, 
    2.018738e-11, 1.897918e-11, 1.903807e-11, 1.900624e-11, 1.906613e-11, 
    1.902392e-11, 1.921202e-11, 1.926862e-11, 1.953475e-11, 1.942527e-11, 
    1.959967e-11, 1.944294e-11, 1.947066e-11, 1.960538e-11, 1.945139e-11, 
    1.978909e-11, 1.955978e-11, 1.998695e-11, 1.975664e-11, 2.000144e-11, 
    1.995685e-11, 2.00307e-11, 2.009698e-11, 2.018054e-11, 2.033525e-11, 
    2.029937e-11, 2.042915e-11, 1.912607e-11, 1.920282e-11, 1.919605e-11, 
    1.927654e-11, 1.93362e-11, 1.946586e-11, 1.967487e-11, 1.959612e-11, 
    1.974083e-11, 1.976996e-11, 1.955016e-11, 1.968495e-11, 1.925428e-11, 
    1.932349e-11, 1.928227e-11, 1.913212e-11, 1.961426e-11, 1.936596e-11, 
    1.982589e-11, 1.969031e-11, 2.008752e-11, 1.988941e-11, 2.027963e-11, 
    2.04478e-11, 2.060681e-11, 2.079357e-11, 1.924478e-11, 1.919254e-11, 
    1.928613e-11, 1.941605e-11, 1.953704e-11, 1.969856e-11, 1.971513e-11, 
    1.97455e-11, 1.982426e-11, 1.989064e-11, 1.975511e-11, 1.990729e-11, 
    1.933957e-11, 1.963589e-11, 1.917282e-11, 1.931159e-11, 1.940838e-11, 
    1.936588e-11, 1.958713e-11, 1.963949e-11, 1.98531e-11, 1.974251e-11, 
    2.040622e-11, 2.0111e-11, 2.093642e-11, 2.070379e-11, 1.917431e-11, 
    1.92446e-11, 1.949038e-11, 1.937321e-11, 1.970937e-11, 1.979264e-11, 
    1.986047e-11, 1.994738e-11, 1.995678e-11, 2.000839e-11, 1.992385e-11, 
    2.000505e-11, 1.969891e-11, 1.983538e-11, 1.946219e-11, 1.955264e-11, 
    1.9511e-11, 1.946538e-11, 1.960637e-11, 1.975724e-11, 1.976046e-11, 
    1.980898e-11, 1.99461e-11, 1.971074e-11, 2.044452e-11, 1.998953e-11, 
    1.932141e-11, 1.945753e-11, 1.947701e-11, 1.942419e-11, 1.978428e-11, 
    1.965336e-11, 2.000713e-11, 1.991116e-11, 2.006855e-11, 1.999025e-11, 
    1.997874e-11, 1.987847e-11, 1.981619e-11, 1.965936e-11, 1.953228e-11, 
    1.943184e-11, 1.945517e-11, 1.956559e-11, 1.976649e-11, 1.995763e-11, 
    1.991567e-11, 2.005656e-11, 1.968489e-11, 1.984025e-11, 1.978012e-11, 
    1.993712e-11, 1.959403e-11, 1.9886e-11, 1.951981e-11, 1.955176e-11, 
    1.965077e-11, 1.985082e-11, 1.989522e-11, 1.994272e-11, 1.99134e-11, 
    1.97716e-11, 1.974842e-11, 1.964836e-11, 1.962078e-11, 1.95448e-11, 
    1.948202e-11, 1.953937e-11, 1.959971e-11, 1.977165e-11, 1.992736e-11, 
    2.009792e-11, 2.013979e-11, 2.034041e-11, 2.017702e-11, 2.044707e-11, 
    2.021736e-11, 2.061597e-11, 1.990298e-11, 2.021061e-11, 1.965528e-11, 
    1.971467e-11, 1.982237e-11, 2.007066e-11, 1.993639e-11, 2.009347e-11, 
    1.974751e-11, 1.956941e-11, 1.952347e-11, 1.943794e-11, 1.952542e-11, 
    1.95183e-11, 1.960221e-11, 1.957522e-11, 1.977738e-11, 1.966864e-11, 
    1.997846e-11, 2.009222e-11, 2.041553e-11, 2.061522e-11, 2.081966e-11, 
    2.09103e-11, 2.093793e-11, 2.094949e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
